magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1260 -1238 2498 2638
<< nwell >>
rect 0 581 1238 1378
rect 0 538 986 581
<< pwell >>
rect 64 36 1187 70
<< mvnmos >>
rect 122 144 322 344
rect 378 144 578 344
rect 764 144 864 344
rect 1056 200 1140 400
<< mvpmos >>
rect 122 604 322 1204
rect 378 604 578 1204
rect 764 604 864 1204
rect 1088 947 1172 1147
<< mvndiff >>
rect 1056 445 1140 456
rect 1056 411 1094 445
rect 1128 411 1140 445
rect 1056 400 1140 411
rect 66 326 122 344
rect 66 292 77 326
rect 111 292 122 326
rect 66 258 122 292
rect 66 224 77 258
rect 111 224 122 258
rect 66 190 122 224
rect 66 156 77 190
rect 111 156 122 190
rect 66 144 122 156
rect 322 326 378 344
rect 322 292 333 326
rect 367 292 378 326
rect 322 258 378 292
rect 322 224 333 258
rect 367 224 378 258
rect 322 190 378 224
rect 322 156 333 190
rect 367 156 378 190
rect 322 144 378 156
rect 578 326 634 344
rect 578 292 589 326
rect 623 292 634 326
rect 578 258 634 292
rect 578 224 589 258
rect 623 224 634 258
rect 578 190 634 224
rect 578 156 589 190
rect 623 156 634 190
rect 578 144 634 156
rect 708 326 764 344
rect 708 292 719 326
rect 753 292 764 326
rect 708 258 764 292
rect 708 224 719 258
rect 753 224 764 258
rect 708 190 764 224
rect 708 156 719 190
rect 753 156 764 190
rect 708 144 764 156
rect 864 326 920 344
rect 864 292 875 326
rect 909 292 920 326
rect 864 258 920 292
rect 864 224 875 258
rect 909 224 920 258
rect 864 190 920 224
rect 864 156 875 190
rect 909 156 920 190
rect 864 144 920 156
rect 1056 189 1140 200
rect 1056 155 1094 189
rect 1128 155 1140 189
rect 1056 144 1140 155
<< mvpdiff >>
rect 66 1192 122 1204
rect 66 1158 77 1192
rect 111 1158 122 1192
rect 66 1124 122 1158
rect 66 1090 77 1124
rect 111 1090 122 1124
rect 66 1056 122 1090
rect 66 1022 77 1056
rect 111 1022 122 1056
rect 66 988 122 1022
rect 66 954 77 988
rect 111 954 122 988
rect 66 920 122 954
rect 66 886 77 920
rect 111 886 122 920
rect 66 852 122 886
rect 66 818 77 852
rect 111 818 122 852
rect 66 784 122 818
rect 66 750 77 784
rect 111 750 122 784
rect 66 716 122 750
rect 66 682 77 716
rect 111 682 122 716
rect 66 604 122 682
rect 322 1192 378 1204
rect 322 1158 333 1192
rect 367 1158 378 1192
rect 322 1124 378 1158
rect 322 1090 333 1124
rect 367 1090 378 1124
rect 322 1056 378 1090
rect 322 1022 333 1056
rect 367 1022 378 1056
rect 322 988 378 1022
rect 322 954 333 988
rect 367 954 378 988
rect 322 920 378 954
rect 322 886 333 920
rect 367 886 378 920
rect 322 852 378 886
rect 322 818 333 852
rect 367 818 378 852
rect 322 784 378 818
rect 322 750 333 784
rect 367 750 378 784
rect 322 716 378 750
rect 322 682 333 716
rect 367 682 378 716
rect 322 604 378 682
rect 578 1192 634 1204
rect 578 1158 589 1192
rect 623 1158 634 1192
rect 578 1124 634 1158
rect 578 1090 589 1124
rect 623 1090 634 1124
rect 578 1056 634 1090
rect 578 1022 589 1056
rect 623 1022 634 1056
rect 578 988 634 1022
rect 578 954 589 988
rect 623 954 634 988
rect 578 920 634 954
rect 578 886 589 920
rect 623 886 634 920
rect 578 852 634 886
rect 578 818 589 852
rect 623 818 634 852
rect 578 784 634 818
rect 578 750 589 784
rect 623 750 634 784
rect 578 716 634 750
rect 578 682 589 716
rect 623 682 634 716
rect 578 604 634 682
rect 708 1192 764 1204
rect 708 1158 719 1192
rect 753 1158 764 1192
rect 708 1124 764 1158
rect 708 1090 719 1124
rect 753 1090 764 1124
rect 708 1056 764 1090
rect 708 1022 719 1056
rect 753 1022 764 1056
rect 708 988 764 1022
rect 708 954 719 988
rect 753 954 764 988
rect 708 920 764 954
rect 708 886 719 920
rect 753 886 764 920
rect 708 852 764 886
rect 708 818 719 852
rect 753 818 764 852
rect 708 784 764 818
rect 708 750 719 784
rect 753 750 764 784
rect 708 716 764 750
rect 708 682 719 716
rect 753 682 764 716
rect 708 604 764 682
rect 864 1192 920 1204
rect 864 1158 875 1192
rect 909 1158 920 1192
rect 864 1124 920 1158
rect 1088 1192 1172 1203
rect 1088 1158 1126 1192
rect 1160 1158 1172 1192
rect 1088 1147 1172 1158
rect 864 1090 875 1124
rect 909 1090 920 1124
rect 864 1056 920 1090
rect 864 1022 875 1056
rect 909 1022 920 1056
rect 864 988 920 1022
rect 864 954 875 988
rect 909 954 920 988
rect 864 920 920 954
rect 864 886 875 920
rect 909 886 920 920
rect 1088 936 1172 947
rect 1088 902 1126 936
rect 1160 902 1172 936
rect 1088 891 1172 902
rect 864 852 920 886
rect 864 818 875 852
rect 909 818 920 852
rect 864 784 920 818
rect 864 750 875 784
rect 909 750 920 784
rect 864 716 920 750
rect 864 682 875 716
rect 909 682 920 716
rect 864 604 920 682
<< mvndiffc >>
rect 1094 411 1128 445
rect 77 292 111 326
rect 77 224 111 258
rect 77 156 111 190
rect 333 292 367 326
rect 333 224 367 258
rect 333 156 367 190
rect 589 292 623 326
rect 589 224 623 258
rect 589 156 623 190
rect 719 292 753 326
rect 719 224 753 258
rect 719 156 753 190
rect 875 292 909 326
rect 875 224 909 258
rect 875 156 909 190
rect 1094 155 1128 189
<< mvpdiffc >>
rect 77 1158 111 1192
rect 77 1090 111 1124
rect 77 1022 111 1056
rect 77 954 111 988
rect 77 886 111 920
rect 77 818 111 852
rect 77 750 111 784
rect 77 682 111 716
rect 333 1158 367 1192
rect 333 1090 367 1124
rect 333 1022 367 1056
rect 333 954 367 988
rect 333 886 367 920
rect 333 818 367 852
rect 333 750 367 784
rect 333 682 367 716
rect 589 1158 623 1192
rect 589 1090 623 1124
rect 589 1022 623 1056
rect 589 954 623 988
rect 589 886 623 920
rect 589 818 623 852
rect 589 750 623 784
rect 589 682 623 716
rect 719 1158 753 1192
rect 719 1090 753 1124
rect 719 1022 753 1056
rect 719 954 753 988
rect 719 886 753 920
rect 719 818 753 852
rect 719 750 753 784
rect 719 682 753 716
rect 875 1158 909 1192
rect 1126 1158 1160 1192
rect 875 1090 909 1124
rect 875 1022 909 1056
rect 875 954 909 988
rect 875 886 909 920
rect 1126 902 1160 936
rect 875 818 909 852
rect 875 750 909 784
rect 875 682 909 716
<< mvpsubdiff >>
rect 64 36 88 70
rect 122 36 156 70
rect 190 36 224 70
rect 258 36 292 70
rect 326 36 360 70
rect 394 36 428 70
rect 462 36 496 70
rect 530 36 564 70
rect 598 36 632 70
rect 666 36 700 70
rect 734 36 768 70
rect 802 36 836 70
rect 870 36 904 70
rect 938 36 972 70
rect 1006 36 1040 70
rect 1074 36 1108 70
rect 1142 36 1187 70
<< mvnsubdiff >>
rect 68 1278 92 1312
rect 126 1278 160 1312
rect 194 1278 228 1312
rect 262 1278 296 1312
rect 330 1278 364 1312
rect 398 1278 432 1312
rect 466 1278 500 1312
rect 534 1278 568 1312
rect 602 1278 636 1312
rect 670 1278 704 1312
rect 738 1278 772 1312
rect 806 1278 840 1312
rect 874 1278 908 1312
rect 942 1278 976 1312
rect 1010 1278 1044 1312
rect 1078 1278 1112 1312
rect 1146 1278 1172 1312
<< mvpsubdiffcont >>
rect 88 36 122 70
rect 156 36 190 70
rect 224 36 258 70
rect 292 36 326 70
rect 360 36 394 70
rect 428 36 462 70
rect 496 36 530 70
rect 564 36 598 70
rect 632 36 666 70
rect 700 36 734 70
rect 768 36 802 70
rect 836 36 870 70
rect 904 36 938 70
rect 972 36 1006 70
rect 1040 36 1074 70
rect 1108 36 1142 70
<< mvnsubdiffcont >>
rect 92 1278 126 1312
rect 160 1278 194 1312
rect 228 1278 262 1312
rect 296 1278 330 1312
rect 364 1278 398 1312
rect 432 1278 466 1312
rect 500 1278 534 1312
rect 568 1278 602 1312
rect 636 1278 670 1312
rect 704 1278 738 1312
rect 772 1278 806 1312
rect 840 1278 874 1312
rect 908 1278 942 1312
rect 976 1278 1010 1312
rect 1044 1278 1078 1312
rect 1112 1278 1146 1312
<< poly >>
rect 122 1204 322 1236
rect 378 1204 578 1236
rect 764 1204 864 1236
rect 990 1131 1088 1147
rect 990 1097 1006 1131
rect 1040 1097 1088 1131
rect 990 997 1088 1097
rect 990 963 1006 997
rect 1040 963 1088 997
rect 990 947 1088 963
rect 1172 947 1204 1147
rect 122 572 322 604
rect 378 572 578 604
rect 764 572 864 604
rect 122 521 579 572
rect 122 487 138 521
rect 172 487 216 521
rect 250 487 294 521
rect 328 487 372 521
rect 406 487 450 521
rect 484 487 529 521
rect 563 487 579 521
rect 122 447 579 487
rect 122 413 138 447
rect 172 413 216 447
rect 250 413 294 447
rect 328 413 372 447
rect 406 413 450 447
rect 484 413 529 447
rect 563 413 579 447
rect 122 376 579 413
rect 697 521 864 572
rect 697 487 713 521
rect 747 487 802 521
rect 836 487 864 521
rect 697 447 864 487
rect 697 413 713 447
rect 747 413 802 447
rect 836 413 864 447
rect 697 376 864 413
rect 1024 399 1056 400
rect 122 344 322 376
rect 378 344 578 376
rect 764 344 864 376
rect 958 383 1056 399
rect 958 349 974 383
rect 1008 349 1056 383
rect 958 249 1056 349
rect 958 215 974 249
rect 1008 215 1056 249
rect 958 200 1056 215
rect 1140 200 1172 400
rect 958 199 1024 200
rect 122 112 322 144
rect 378 112 578 144
rect 764 112 864 144
<< polycont >>
rect 1006 1097 1040 1131
rect 1006 963 1040 997
rect 138 487 172 521
rect 216 487 250 521
rect 294 487 328 521
rect 372 487 406 521
rect 450 487 484 521
rect 529 487 563 521
rect 138 413 172 447
rect 216 413 250 447
rect 294 413 328 447
rect 372 413 406 447
rect 450 413 484 447
rect 529 413 563 447
rect 713 487 747 521
rect 802 487 836 521
rect 713 413 747 447
rect 802 413 836 447
rect 974 349 1008 383
rect 974 215 1008 249
<< locali >>
rect 68 1278 80 1312
rect 126 1278 152 1312
rect 194 1278 224 1312
rect 262 1278 296 1312
rect 330 1278 364 1312
rect 402 1278 432 1312
rect 474 1278 500 1312
rect 546 1278 568 1312
rect 618 1278 636 1312
rect 690 1278 704 1312
rect 762 1278 772 1312
rect 834 1278 840 1312
rect 906 1278 908 1312
rect 942 1278 944 1312
rect 1010 1278 1016 1312
rect 1078 1278 1088 1312
rect 1146 1278 1172 1312
rect 77 1136 111 1158
rect 77 1064 111 1090
rect 77 992 111 1022
rect 77 920 111 954
rect 77 852 111 886
rect 77 784 111 814
rect 77 716 111 742
rect 77 666 111 670
rect 333 1136 367 1158
rect 333 1064 367 1090
rect 333 992 367 1022
rect 333 920 367 954
rect 333 852 367 886
rect 333 784 367 814
rect 333 716 367 742
rect 333 666 367 670
rect 589 1136 623 1158
rect 589 1064 623 1090
rect 589 992 623 1022
rect 589 920 623 954
rect 589 852 623 886
rect 589 784 623 814
rect 589 716 623 742
rect 589 666 623 670
rect 719 1136 753 1158
rect 719 1064 753 1090
rect 719 992 753 1022
rect 719 920 753 954
rect 719 852 753 886
rect 719 784 753 814
rect 719 716 753 742
rect 719 666 753 670
rect 1110 1158 1126 1192
rect 875 1136 909 1158
rect 875 1064 909 1090
rect 875 992 909 1022
rect 875 920 909 954
rect 1006 1135 1040 1147
rect 1006 997 1040 1097
rect 1006 947 1040 959
rect 1110 902 1126 936
rect 875 852 909 886
rect 875 784 909 814
rect 875 716 909 742
rect 875 666 909 670
rect 122 521 579 523
rect 122 487 138 521
rect 172 492 216 521
rect 250 492 294 521
rect 180 487 216 492
rect 252 487 294 492
rect 328 487 372 521
rect 406 487 450 521
rect 484 487 529 521
rect 563 487 579 521
rect 122 458 146 487
rect 180 458 218 487
rect 252 458 579 487
rect 122 447 579 458
rect 122 413 138 447
rect 172 413 216 447
rect 250 413 294 447
rect 328 413 372 447
rect 406 413 450 447
rect 484 413 529 447
rect 563 413 579 447
rect 122 410 579 413
rect 697 521 864 523
rect 697 492 713 521
rect 747 492 802 521
rect 697 458 710 492
rect 747 487 782 492
rect 836 487 864 521
rect 744 458 782 487
rect 816 458 864 487
rect 697 447 864 458
rect 697 413 713 447
rect 747 413 802 447
rect 836 413 864 447
rect 697 410 864 413
rect 1078 411 1094 445
rect 974 383 1008 399
rect 77 326 111 342
rect 77 258 111 284
rect 77 190 111 212
rect 333 326 367 342
rect 333 258 367 284
rect 333 190 367 212
rect 589 326 623 342
rect 589 258 623 284
rect 589 190 623 212
rect 719 326 753 342
rect 719 258 753 284
rect 719 190 753 212
rect 875 326 909 342
rect 875 258 909 284
rect 875 190 909 212
rect 974 317 1008 349
rect 974 249 1008 283
rect 974 175 1008 215
rect 1078 155 1094 189
rect 64 36 76 70
rect 122 36 148 70
rect 190 36 220 70
rect 258 36 292 70
rect 326 36 360 70
rect 398 36 428 70
rect 470 36 496 70
rect 542 36 564 70
rect 614 36 632 70
rect 686 36 700 70
rect 758 36 768 70
rect 830 36 836 70
rect 902 36 904 70
rect 938 36 940 70
rect 1006 36 1012 70
rect 1074 36 1084 70
rect 1142 36 1187 70
<< viali >>
rect 80 1278 92 1312
rect 92 1278 114 1312
rect 152 1278 160 1312
rect 160 1278 186 1312
rect 224 1278 228 1312
rect 228 1278 258 1312
rect 296 1278 330 1312
rect 368 1278 398 1312
rect 398 1278 402 1312
rect 440 1278 466 1312
rect 466 1278 474 1312
rect 512 1278 534 1312
rect 534 1278 546 1312
rect 584 1278 602 1312
rect 602 1278 618 1312
rect 656 1278 670 1312
rect 670 1278 690 1312
rect 728 1278 738 1312
rect 738 1278 762 1312
rect 800 1278 806 1312
rect 806 1278 834 1312
rect 872 1278 874 1312
rect 874 1278 906 1312
rect 944 1278 976 1312
rect 976 1278 978 1312
rect 1016 1278 1044 1312
rect 1044 1278 1050 1312
rect 1088 1278 1112 1312
rect 1112 1278 1122 1312
rect 77 1192 111 1208
rect 77 1174 111 1192
rect 77 1124 111 1136
rect 77 1102 111 1124
rect 77 1056 111 1064
rect 77 1030 111 1056
rect 77 988 111 992
rect 77 958 111 988
rect 77 886 111 920
rect 77 818 111 848
rect 77 814 111 818
rect 77 750 111 776
rect 77 742 111 750
rect 77 682 111 704
rect 77 670 111 682
rect 333 1192 367 1208
rect 333 1174 367 1192
rect 333 1124 367 1136
rect 333 1102 367 1124
rect 333 1056 367 1064
rect 333 1030 367 1056
rect 333 988 367 992
rect 333 958 367 988
rect 333 886 367 920
rect 333 818 367 848
rect 333 814 367 818
rect 333 750 367 776
rect 333 742 367 750
rect 333 682 367 704
rect 333 670 367 682
rect 589 1192 623 1208
rect 589 1174 623 1192
rect 589 1124 623 1136
rect 589 1102 623 1124
rect 589 1056 623 1064
rect 589 1030 623 1056
rect 589 988 623 992
rect 589 958 623 988
rect 589 886 623 920
rect 589 818 623 848
rect 589 814 623 818
rect 589 750 623 776
rect 589 742 623 750
rect 589 682 623 704
rect 589 670 623 682
rect 719 1192 753 1208
rect 719 1174 753 1192
rect 719 1124 753 1136
rect 719 1102 753 1124
rect 719 1056 753 1064
rect 719 1030 753 1056
rect 719 988 753 992
rect 719 958 753 988
rect 719 886 753 920
rect 719 818 753 848
rect 719 814 753 818
rect 719 750 753 776
rect 719 742 753 750
rect 719 682 753 704
rect 719 670 753 682
rect 875 1192 909 1208
rect 875 1174 909 1192
rect 1142 1158 1160 1192
rect 1160 1158 1176 1192
rect 875 1124 909 1136
rect 875 1102 909 1124
rect 875 1056 909 1064
rect 875 1030 909 1056
rect 875 988 909 992
rect 875 958 909 988
rect 1006 1131 1040 1135
rect 1006 1101 1040 1131
rect 1006 963 1040 993
rect 1006 959 1040 963
rect 875 886 909 920
rect 1142 902 1160 936
rect 1160 902 1176 936
rect 875 818 909 848
rect 875 814 909 818
rect 875 750 909 776
rect 875 742 909 750
rect 875 682 909 704
rect 875 670 909 682
rect 146 487 172 492
rect 172 487 180 492
rect 218 487 250 492
rect 250 487 252 492
rect 146 458 180 487
rect 218 458 252 487
rect 710 487 713 492
rect 713 487 744 492
rect 782 487 802 492
rect 802 487 816 492
rect 710 458 744 487
rect 782 458 816 487
rect 1110 411 1128 445
rect 1128 411 1144 445
rect 77 292 111 318
rect 77 284 111 292
rect 77 224 111 246
rect 77 212 111 224
rect 77 156 111 174
rect 77 140 111 156
rect 333 292 367 318
rect 333 284 367 292
rect 333 224 367 246
rect 333 212 367 224
rect 333 156 367 174
rect 333 140 367 156
rect 589 292 623 318
rect 589 284 623 292
rect 589 224 623 246
rect 589 212 623 224
rect 589 156 623 174
rect 589 140 623 156
rect 719 292 753 318
rect 719 284 753 292
rect 719 224 753 246
rect 719 212 753 224
rect 719 156 753 174
rect 719 140 753 156
rect 875 292 909 318
rect 875 284 909 292
rect 875 224 909 246
rect 875 212 909 224
rect 875 156 909 174
rect 875 140 909 156
rect 974 283 1008 317
rect 974 141 1008 175
rect 1110 155 1128 189
rect 1128 155 1144 189
rect 76 36 88 70
rect 88 36 110 70
rect 148 36 156 70
rect 156 36 182 70
rect 220 36 224 70
rect 224 36 254 70
rect 292 36 326 70
rect 364 36 394 70
rect 394 36 398 70
rect 436 36 462 70
rect 462 36 470 70
rect 508 36 530 70
rect 530 36 542 70
rect 580 36 598 70
rect 598 36 614 70
rect 652 36 666 70
rect 666 36 686 70
rect 724 36 734 70
rect 734 36 758 70
rect 796 36 802 70
rect 802 36 830 70
rect 868 36 870 70
rect 870 36 902 70
rect 940 36 972 70
rect 972 36 974 70
rect 1012 36 1040 70
rect 1040 36 1046 70
rect 1084 36 1108 70
rect 1108 36 1118 70
<< metal1 >>
rect 68 1321 1172 1324
rect 68 1318 144 1321
rect 120 1269 144 1318
rect 196 1269 209 1321
rect 261 1269 274 1321
rect 326 1312 339 1321
rect 391 1312 404 1321
rect 456 1312 469 1321
rect 521 1312 534 1321
rect 586 1312 599 1321
rect 651 1312 664 1321
rect 716 1312 729 1321
rect 330 1278 339 1312
rect 402 1278 404 1312
rect 651 1278 656 1312
rect 716 1278 728 1312
rect 326 1269 339 1278
rect 391 1269 404 1278
rect 456 1269 469 1278
rect 521 1269 534 1278
rect 586 1269 599 1278
rect 651 1269 664 1278
rect 716 1269 729 1278
rect 781 1269 794 1321
rect 846 1269 858 1321
rect 910 1269 922 1321
rect 974 1312 986 1321
rect 1038 1312 1050 1321
rect 1102 1312 1114 1321
rect 978 1278 986 1312
rect 974 1269 986 1278
rect 1038 1269 1050 1278
rect 1102 1269 1114 1278
rect 1166 1269 1172 1321
rect 120 1266 1172 1269
rect 68 1234 131 1266
rect 120 1220 131 1234
tri 131 1220 177 1266 nw
tri 120 1209 131 1220 nw
rect 68 1174 77 1182
rect 111 1174 120 1182
rect 68 1149 120 1174
rect 68 1064 120 1097
rect 68 1006 120 1012
tri 68 1003 71 1006 ne
rect 71 992 117 1006
tri 117 1003 120 1006 nw
rect 327 1208 373 1220
rect 327 1174 333 1208
rect 367 1174 373 1208
rect 327 1136 373 1174
rect 327 1102 333 1136
rect 367 1102 373 1136
rect 327 1064 373 1102
rect 327 1030 333 1064
rect 367 1030 373 1064
rect 71 958 77 992
rect 111 958 117 992
rect 327 992 373 1030
rect 583 1208 629 1220
rect 583 1174 589 1208
rect 623 1174 629 1208
rect 583 1136 629 1174
rect 583 1102 589 1136
rect 623 1102 629 1136
rect 583 1064 629 1102
rect 583 1030 589 1064
rect 623 1030 629 1064
rect 583 992 629 1030
rect 710 1214 762 1220
rect 710 1139 762 1162
rect 710 1064 762 1087
rect 710 1006 762 1012
tri 710 1003 713 1006 ne
tri 303 958 327 982 se
rect 327 958 333 992
rect 367 958 373 992
tri 373 958 407 992 sw
rect 583 958 589 992
rect 623 958 629 992
rect 71 920 117 958
rect 71 886 77 920
rect 111 886 117 920
tri 291 946 303 958 se
rect 303 946 407 958
tri 407 946 419 958 sw
rect 291 894 297 946
rect 349 920 361 946
rect 413 894 419 946
tri 291 886 299 894 ne
rect 299 886 333 894
rect 367 886 411 894
tri 411 886 419 894 nw
rect 583 920 629 958
rect 583 886 589 920
rect 623 886 629 920
rect 71 848 117 886
tri 299 858 327 886 ne
rect 327 883 408 886
tri 408 883 411 886 nw
rect 71 814 77 848
rect 111 814 117 848
rect 71 776 117 814
rect 71 742 77 776
rect 111 742 117 776
rect 71 704 117 742
rect 71 670 77 704
rect 111 670 117 704
rect 71 658 117 670
rect 327 848 373 883
tri 373 848 408 883 nw
rect 583 848 629 886
rect 327 814 333 848
rect 367 814 373 848
rect 327 776 373 814
rect 327 742 333 776
rect 367 742 373 776
rect 327 704 373 742
rect 327 670 333 704
rect 367 670 373 704
rect 327 658 373 670
rect 583 814 589 848
rect 623 814 629 848
rect 583 776 629 814
rect 583 742 589 776
rect 623 742 629 776
rect 583 704 629 742
rect 583 670 589 704
rect 623 670 629 704
rect 583 498 629 670
rect 713 992 759 1006
tri 759 1003 762 1006 nw
rect 869 1208 915 1220
rect 869 1174 875 1208
rect 909 1192 915 1208
tri 915 1192 943 1220 sw
rect 909 1174 943 1192
rect 869 1158 943 1174
tri 943 1158 977 1192 sw
rect 869 1147 977 1158
tri 977 1147 988 1158 sw
rect 1097 1152 1103 1204
rect 1155 1192 1167 1204
rect 1155 1152 1167 1158
rect 1219 1152 1225 1204
rect 869 1136 1046 1147
rect 869 1102 875 1136
rect 909 1135 1046 1136
rect 909 1102 1006 1135
rect 869 1101 1006 1102
rect 1040 1101 1046 1135
rect 869 1064 1046 1101
rect 869 1030 875 1064
rect 909 1030 1046 1064
rect 713 958 719 992
rect 753 958 759 992
rect 713 920 759 958
rect 713 886 719 920
rect 753 886 759 920
rect 713 848 759 886
rect 713 814 719 848
rect 753 814 759 848
rect 713 776 759 814
rect 713 742 719 776
rect 753 742 759 776
rect 713 704 759 742
rect 713 670 719 704
rect 753 670 759 704
rect 713 658 759 670
rect 869 993 1046 1030
rect 869 992 1006 993
rect 869 958 875 992
rect 909 959 1006 992
rect 1040 959 1046 993
rect 909 958 1046 959
rect 869 947 1046 958
rect 869 936 968 947
tri 968 936 979 947 nw
rect 869 920 934 936
rect 869 886 875 920
rect 909 902 934 920
tri 934 902 968 936 nw
rect 909 886 915 902
rect 869 848 915 886
tri 915 883 934 902 nw
rect 1093 894 1099 946
rect 1151 936 1163 946
rect 1151 894 1163 902
rect 1215 894 1221 946
rect 869 814 875 848
rect 909 814 915 848
rect 869 776 915 814
rect 869 742 875 776
rect 909 742 915 776
rect 869 704 915 742
tri 915 708 963 756 sw
rect 869 670 875 704
rect 909 670 915 704
tri 629 498 668 537 sw
rect 134 492 264 498
rect 134 458 146 492
rect 180 458 218 492
rect 252 458 264 492
rect 134 452 264 458
rect 583 492 828 498
rect 583 458 710 492
rect 744 458 782 492
rect 816 458 828 492
rect 583 452 828 458
rect 583 445 661 452
tri 661 445 668 452 nw
rect 71 318 117 330
rect 71 284 77 318
rect 111 284 117 318
tri 68 248 71 251 se
rect 71 248 117 284
rect 291 294 297 346
rect 349 318 361 346
rect 413 294 419 346
rect 291 284 333 294
rect 367 284 409 294
tri 409 284 419 294 nw
rect 583 318 629 445
tri 629 413 661 445 nw
rect 869 330 915 670
tri 915 529 963 577 nw
rect 1028 401 1034 453
rect 1086 401 1098 453
rect 1150 401 1156 453
tri 915 330 975 390 sw
rect 583 284 589 318
rect 623 284 629 318
tri 291 283 292 284 ne
rect 292 283 408 284
tri 408 283 409 284 nw
tri 292 251 324 283 ne
rect 324 251 376 283
tri 376 251 408 283 nw
tri 117 248 120 251 sw
tri 324 248 327 251 ne
rect 68 246 120 248
rect 68 242 77 246
rect 111 242 120 246
rect 68 178 120 190
rect 327 246 373 251
tri 373 248 376 251 nw
rect 327 212 333 246
rect 367 212 373 246
rect 327 174 373 212
rect 327 140 333 174
rect 367 140 373 174
tri 120 129 125 134 sw
rect 120 126 125 129
rect 68 120 125 126
tri 125 120 134 129 sw
rect 327 128 373 140
rect 583 246 629 284
rect 713 318 759 330
rect 713 284 719 318
rect 753 284 759 318
rect 583 212 589 246
rect 623 212 629 246
rect 583 174 629 212
rect 583 140 589 174
rect 623 140 629 174
rect 583 128 629 140
tri 710 248 713 251 se
rect 713 248 759 284
rect 869 329 975 330
tri 975 329 976 330 sw
rect 869 318 1014 329
rect 869 284 875 318
rect 909 317 1014 318
rect 909 284 974 317
rect 869 283 974 284
rect 1008 283 1014 317
tri 759 248 762 251 sw
rect 710 246 762 248
rect 710 242 719 246
rect 753 242 762 246
rect 710 178 762 190
rect 869 246 1014 283
rect 869 212 875 246
rect 909 212 1014 246
rect 869 175 1014 212
rect 869 174 974 175
rect 869 140 875 174
rect 909 141 974 174
rect 1008 141 1014 175
rect 1073 146 1079 198
rect 1131 189 1143 198
rect 1131 146 1143 155
rect 1195 146 1201 198
rect 909 140 1014 141
rect 869 128 1014 140
rect 710 120 762 126
tri 64 82 68 86 se
rect 68 82 134 120
tri 134 82 172 120 sw
rect 64 79 1187 82
rect 64 27 70 79
rect 122 27 137 79
rect 189 27 204 79
rect 256 27 271 79
rect 323 70 337 79
rect 389 70 403 79
rect 455 70 469 79
rect 521 70 535 79
rect 587 70 601 79
rect 653 70 667 79
rect 719 70 733 79
rect 785 70 799 79
rect 326 36 337 70
rect 398 36 403 70
rect 719 36 724 70
rect 785 36 796 70
rect 323 27 337 36
rect 389 27 403 36
rect 455 27 469 36
rect 521 27 535 36
rect 587 27 601 36
rect 653 27 667 36
rect 719 27 733 36
rect 785 27 799 36
rect 851 27 865 79
rect 917 27 931 79
rect 983 27 997 79
rect 1049 27 1063 79
rect 1115 70 1129 79
rect 1118 36 1129 70
rect 1115 27 1129 36
rect 1181 27 1187 79
rect 64 24 1187 27
<< via1 >>
rect 68 1312 120 1318
rect 68 1278 80 1312
rect 80 1278 114 1312
rect 114 1278 120 1312
rect 68 1266 120 1278
rect 144 1312 196 1321
rect 144 1278 152 1312
rect 152 1278 186 1312
rect 186 1278 196 1312
rect 144 1269 196 1278
rect 209 1312 261 1321
rect 209 1278 224 1312
rect 224 1278 258 1312
rect 258 1278 261 1312
rect 209 1269 261 1278
rect 274 1312 326 1321
rect 339 1312 391 1321
rect 404 1312 456 1321
rect 469 1312 521 1321
rect 534 1312 586 1321
rect 599 1312 651 1321
rect 664 1312 716 1321
rect 729 1312 781 1321
rect 274 1278 296 1312
rect 296 1278 326 1312
rect 339 1278 368 1312
rect 368 1278 391 1312
rect 404 1278 440 1312
rect 440 1278 456 1312
rect 469 1278 474 1312
rect 474 1278 512 1312
rect 512 1278 521 1312
rect 534 1278 546 1312
rect 546 1278 584 1312
rect 584 1278 586 1312
rect 599 1278 618 1312
rect 618 1278 651 1312
rect 664 1278 690 1312
rect 690 1278 716 1312
rect 729 1278 762 1312
rect 762 1278 781 1312
rect 274 1269 326 1278
rect 339 1269 391 1278
rect 404 1269 456 1278
rect 469 1269 521 1278
rect 534 1269 586 1278
rect 599 1269 651 1278
rect 664 1269 716 1278
rect 729 1269 781 1278
rect 794 1312 846 1321
rect 794 1278 800 1312
rect 800 1278 834 1312
rect 834 1278 846 1312
rect 794 1269 846 1278
rect 858 1312 910 1321
rect 858 1278 872 1312
rect 872 1278 906 1312
rect 906 1278 910 1312
rect 858 1269 910 1278
rect 922 1312 974 1321
rect 986 1312 1038 1321
rect 1050 1312 1102 1321
rect 1114 1312 1166 1321
rect 922 1278 944 1312
rect 944 1278 974 1312
rect 986 1278 1016 1312
rect 1016 1278 1038 1312
rect 1050 1278 1088 1312
rect 1088 1278 1102 1312
rect 1114 1278 1122 1312
rect 1122 1278 1166 1312
rect 922 1269 974 1278
rect 986 1269 1038 1278
rect 1050 1269 1102 1278
rect 1114 1269 1166 1278
rect 68 1208 120 1234
rect 68 1182 77 1208
rect 77 1182 111 1208
rect 111 1182 120 1208
rect 68 1136 120 1149
rect 68 1102 77 1136
rect 77 1102 111 1136
rect 111 1102 120 1136
rect 68 1097 120 1102
rect 68 1030 77 1064
rect 77 1030 111 1064
rect 111 1030 120 1064
rect 68 1012 120 1030
rect 710 1208 762 1214
rect 710 1174 719 1208
rect 719 1174 753 1208
rect 753 1174 762 1208
rect 710 1162 762 1174
rect 710 1136 762 1139
rect 710 1102 719 1136
rect 719 1102 753 1136
rect 753 1102 762 1136
rect 710 1087 762 1102
rect 710 1030 719 1064
rect 719 1030 753 1064
rect 753 1030 762 1064
rect 710 1012 762 1030
rect 297 920 349 946
rect 361 920 413 946
rect 297 894 333 920
rect 333 894 349 920
rect 361 894 367 920
rect 367 894 413 920
rect 1103 1192 1155 1204
rect 1167 1192 1219 1204
rect 1103 1158 1142 1192
rect 1142 1158 1155 1192
rect 1167 1158 1176 1192
rect 1176 1158 1219 1192
rect 1103 1152 1155 1158
rect 1167 1152 1219 1158
rect 1099 936 1151 946
rect 1163 936 1215 946
rect 1099 902 1142 936
rect 1142 902 1151 936
rect 1163 902 1176 936
rect 1176 902 1215 936
rect 1099 894 1151 902
rect 1163 894 1215 902
rect 297 318 349 346
rect 361 318 413 346
rect 297 294 333 318
rect 333 294 349 318
rect 361 294 367 318
rect 367 294 413 318
rect 1034 401 1086 453
rect 1098 445 1150 453
rect 1098 411 1110 445
rect 1110 411 1144 445
rect 1144 411 1150 445
rect 1098 401 1150 411
rect 68 212 77 242
rect 77 212 111 242
rect 111 212 120 242
rect 68 190 120 212
rect 68 174 120 178
rect 68 140 77 174
rect 77 140 111 174
rect 111 140 120 174
rect 68 126 120 140
rect 710 212 719 242
rect 719 212 753 242
rect 753 212 762 242
rect 710 190 762 212
rect 710 174 762 178
rect 710 140 719 174
rect 719 140 753 174
rect 753 140 762 174
rect 710 126 762 140
rect 1079 189 1131 198
rect 1143 189 1195 198
rect 1079 155 1110 189
rect 1110 155 1131 189
rect 1143 155 1144 189
rect 1144 155 1195 189
rect 1079 146 1131 155
rect 1143 146 1195 155
rect 70 70 122 79
rect 70 36 76 70
rect 76 36 110 70
rect 110 36 122 70
rect 70 27 122 36
rect 137 70 189 79
rect 137 36 148 70
rect 148 36 182 70
rect 182 36 189 70
rect 137 27 189 36
rect 204 70 256 79
rect 204 36 220 70
rect 220 36 254 70
rect 254 36 256 70
rect 204 27 256 36
rect 271 70 323 79
rect 337 70 389 79
rect 403 70 455 79
rect 469 70 521 79
rect 535 70 587 79
rect 601 70 653 79
rect 667 70 719 79
rect 733 70 785 79
rect 799 70 851 79
rect 271 36 292 70
rect 292 36 323 70
rect 337 36 364 70
rect 364 36 389 70
rect 403 36 436 70
rect 436 36 455 70
rect 469 36 470 70
rect 470 36 508 70
rect 508 36 521 70
rect 535 36 542 70
rect 542 36 580 70
rect 580 36 587 70
rect 601 36 614 70
rect 614 36 652 70
rect 652 36 653 70
rect 667 36 686 70
rect 686 36 719 70
rect 733 36 758 70
rect 758 36 785 70
rect 799 36 830 70
rect 830 36 851 70
rect 271 27 323 36
rect 337 27 389 36
rect 403 27 455 36
rect 469 27 521 36
rect 535 27 587 36
rect 601 27 653 36
rect 667 27 719 36
rect 733 27 785 36
rect 799 27 851 36
rect 865 70 917 79
rect 865 36 868 70
rect 868 36 902 70
rect 902 36 917 70
rect 865 27 917 36
rect 931 70 983 79
rect 931 36 940 70
rect 940 36 974 70
rect 974 36 983 70
rect 931 27 983 36
rect 997 70 1049 79
rect 997 36 1012 70
rect 1012 36 1046 70
rect 1046 36 1049 70
rect 997 27 1049 36
rect 1063 70 1115 79
rect 1063 36 1084 70
rect 1084 36 1115 70
rect 1063 27 1115 36
rect 1129 27 1181 79
<< metal2 >>
rect 8 1321 1232 1360
rect 8 1318 144 1321
rect 8 1266 68 1318
rect 120 1269 144 1318
rect 196 1269 209 1321
rect 261 1269 274 1321
rect 326 1269 339 1321
rect 391 1269 404 1321
rect 456 1269 469 1321
rect 521 1269 534 1321
rect 586 1269 599 1321
rect 651 1269 664 1321
rect 716 1269 729 1321
rect 781 1269 794 1321
rect 846 1269 858 1321
rect 910 1269 922 1321
rect 974 1269 986 1321
rect 1038 1269 1050 1321
rect 1102 1269 1114 1321
rect 1166 1269 1232 1321
rect 120 1266 1232 1269
rect 8 1234 1232 1266
rect 8 1182 68 1234
rect 120 1214 1232 1234
rect 120 1182 710 1214
rect 8 1162 710 1182
rect 762 1204 1232 1214
rect 762 1162 1103 1204
rect 8 1152 1103 1162
rect 1155 1152 1167 1204
rect 1219 1152 1232 1204
rect 8 1149 1232 1152
rect 8 1097 68 1149
rect 120 1139 1232 1149
rect 120 1097 710 1139
rect 8 1087 710 1097
rect 762 1087 1232 1139
rect 8 1064 1232 1087
rect 8 1012 68 1064
rect 120 1012 710 1064
rect 762 1012 1232 1064
rect 8 1006 1232 1012
rect 291 894 297 946
rect 349 894 361 946
rect 413 894 1099 946
rect 1151 894 1163 946
rect 1215 894 1221 946
rect 1028 401 1034 453
rect 1086 401 1098 453
rect 1150 401 1156 453
tri 1013 356 1028 371 se
rect 1028 356 1156 401
tri 1003 346 1013 356 se
rect 1013 346 1094 356
rect 291 294 297 346
rect 349 294 361 346
rect 413 294 1094 346
tri 1094 294 1156 356 nw
rect 53 242 1212 248
rect 53 190 68 242
rect 120 190 710 242
rect 762 198 1212 242
rect 762 190 1079 198
rect 53 178 1079 190
rect 53 126 68 178
rect 120 126 710 178
rect 762 146 1079 178
rect 1131 146 1143 198
rect 1195 146 1212 198
rect 762 126 1212 146
rect 53 79 1212 126
rect 53 27 70 79
rect 122 27 137 79
rect 189 27 204 79
rect 256 27 271 79
rect 323 27 337 79
rect 389 27 403 79
rect 455 27 469 79
rect 521 27 535 79
rect 587 27 601 79
rect 653 27 667 79
rect 719 27 733 79
rect 785 27 799 79
rect 851 27 865 79
rect 917 27 931 79
rect 983 27 997 79
rect 1049 27 1063 79
rect 1115 27 1129 79
rect 1181 27 1212 79
rect 53 22 1212 27
use sky130_fd_pr__nfet_01v8__example_55959141808723  sky130_fd_pr__nfet_01v8__example_55959141808723_0
timestamp 1619729480
transform 1 0 122 0 1 144
box -28 0 228 85
use sky130_fd_pr__nfet_01v8__example_55959141808723  sky130_fd_pr__nfet_01v8__example_55959141808723_1
timestamp 1619729480
transform 1 0 378 0 1 144
box -28 0 228 85
use sky130_fd_pr__nfet_01v8__example_55959141808722  sky130_fd_pr__nfet_01v8__example_55959141808722_0
timestamp 1619729480
transform 1 0 764 0 1 144
box -28 0 128 85
use sky130_fd_pr__nfet_01v8__example_55959141808721  sky130_fd_pr__nfet_01v8__example_55959141808721_0
timestamp 1619729480
transform 0 -1 1140 1 0 200
box -28 0 228 13
use sky130_fd_pr__pfet_01v8__example_55959141808720  sky130_fd_pr__pfet_01v8__example_55959141808720_0
timestamp 1619729480
transform 1 0 378 0 -1 1204
box -28 0 228 265
use sky130_fd_pr__pfet_01v8__example_55959141808720  sky130_fd_pr__pfet_01v8__example_55959141808720_1
timestamp 1619729480
transform 1 0 122 0 -1 1204
box -28 0 228 265
use sky130_fd_pr__pfet_01v8__example_55959141808718  sky130_fd_pr__pfet_01v8__example_55959141808718_0
timestamp 1619729480
transform 1 0 764 0 -1 1204
box -28 0 128 265
use sky130_fd_pr__pfet_01v8__example_55959141808716  sky130_fd_pr__pfet_01v8__example_55959141808716_0
timestamp 1619729480
transform 0 -1 1172 -1 0 1147
box -28 0 228 13
<< labels >>
flabel metal2 s 14 1006 329 1360 3 FreeSans 520 0 0 0 VCC_IO
flabel metal2 s 208 69 322 190 3 FreeSans 520 0 0 0 VSSD
flabel metal1 s 870 409 909 550 3 FreeSans 520 0 0 0 OUT_H
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 5015808
string GDS_START 4999354
<< end >>
