magic
tech sky130A
magscale 1 2
timestamp 1640697675
<< dnwell >>
rect 80 80 1644 1844
<< nwell >>
rect 0 1564 1724 1924
rect 0 360 360 1564
rect 1364 360 1724 1564
rect 0 0 1724 360
<< pbase >>
rect 360 360 1364 1564
<< npn2p00 >>
rect 360 360 1364 1564
<< ndiff >>
rect 762 1149 962 1162
rect 762 775 777 1149
rect 947 775 962 1149
rect 762 762 962 775
<< ndiffc >>
rect 777 775 947 1149
<< psubdiff >>
rect 520 1380 1204 1404
rect 520 1346 544 1380
rect 578 1346 641 1380
rect 675 1346 709 1380
rect 743 1346 777 1380
rect 811 1346 845 1380
rect 879 1346 913 1380
rect 947 1346 981 1380
rect 1015 1346 1049 1380
rect 1083 1346 1146 1380
rect 1180 1346 1204 1380
rect 520 1322 1204 1346
rect 520 1285 602 1322
rect 520 1251 544 1285
rect 578 1251 602 1285
rect 520 1217 602 1251
rect 520 1183 544 1217
rect 578 1183 602 1217
rect 520 1149 602 1183
rect 1122 1285 1204 1322
rect 1122 1251 1146 1285
rect 1180 1251 1204 1285
rect 1122 1217 1204 1251
rect 1122 1183 1146 1217
rect 1180 1183 1204 1217
rect 520 1115 544 1149
rect 578 1115 602 1149
rect 520 1081 602 1115
rect 520 1047 544 1081
rect 578 1047 602 1081
rect 520 1013 602 1047
rect 520 979 544 1013
rect 578 979 602 1013
rect 520 945 602 979
rect 520 911 544 945
rect 578 911 602 945
rect 520 877 602 911
rect 520 843 544 877
rect 578 843 602 877
rect 520 809 602 843
rect 520 775 544 809
rect 578 775 602 809
rect 520 741 602 775
rect 1122 1149 1204 1183
rect 1122 1115 1146 1149
rect 1180 1115 1204 1149
rect 1122 1081 1204 1115
rect 1122 1047 1146 1081
rect 1180 1047 1204 1081
rect 1122 1013 1204 1047
rect 1122 979 1146 1013
rect 1180 979 1204 1013
rect 1122 945 1204 979
rect 1122 911 1146 945
rect 1180 911 1204 945
rect 1122 877 1204 911
rect 1122 843 1146 877
rect 1180 843 1204 877
rect 1122 809 1204 843
rect 1122 775 1146 809
rect 1180 775 1204 809
rect 520 707 544 741
rect 578 707 602 741
rect 520 673 602 707
rect 520 639 544 673
rect 578 639 602 673
rect 520 602 602 639
rect 1122 741 1204 775
rect 1122 707 1146 741
rect 1180 707 1204 741
rect 1122 673 1204 707
rect 1122 639 1146 673
rect 1180 639 1204 673
rect 1122 602 1204 639
rect 520 578 1204 602
rect 520 544 544 578
rect 578 544 641 578
rect 675 544 709 578
rect 743 544 777 578
rect 811 544 845 578
rect 879 544 913 578
rect 947 544 981 578
rect 1015 544 1049 578
rect 1083 544 1146 578
rect 1180 544 1204 578
rect 520 520 1204 544
<< nsubdiff >>
rect 118 1782 1606 1806
rect 118 1748 142 1782
rect 176 1748 233 1782
rect 267 1748 301 1782
rect 335 1748 369 1782
rect 403 1748 437 1782
rect 471 1748 505 1782
rect 539 1748 573 1782
rect 607 1748 641 1782
rect 675 1748 709 1782
rect 743 1748 777 1782
rect 811 1748 845 1782
rect 879 1748 913 1782
rect 947 1748 981 1782
rect 1015 1748 1049 1782
rect 1083 1748 1117 1782
rect 1151 1748 1185 1782
rect 1219 1748 1253 1782
rect 1287 1748 1321 1782
rect 1355 1748 1389 1782
rect 1423 1748 1457 1782
rect 1491 1748 1548 1782
rect 1582 1748 1606 1782
rect 118 1724 1606 1748
rect 118 1693 200 1724
rect 118 1659 142 1693
rect 176 1659 200 1693
rect 118 1625 200 1659
rect 118 1591 142 1625
rect 176 1591 200 1625
rect 118 1557 200 1591
rect 118 1523 142 1557
rect 176 1523 200 1557
rect 118 1489 200 1523
rect 118 1455 142 1489
rect 176 1455 200 1489
rect 118 1421 200 1455
rect 118 1387 142 1421
rect 176 1387 200 1421
rect 1524 1693 1606 1724
rect 1524 1659 1548 1693
rect 1582 1659 1606 1693
rect 1524 1625 1606 1659
rect 1524 1591 1548 1625
rect 1582 1591 1606 1625
rect 1524 1557 1606 1591
rect 1524 1523 1548 1557
rect 1582 1523 1606 1557
rect 1524 1489 1606 1523
rect 1524 1455 1548 1489
rect 1582 1455 1606 1489
rect 1524 1421 1606 1455
rect 118 1353 200 1387
rect 118 1319 142 1353
rect 176 1319 200 1353
rect 118 1285 200 1319
rect 118 1251 142 1285
rect 176 1251 200 1285
rect 118 1217 200 1251
rect 118 1183 142 1217
rect 176 1183 200 1217
rect 118 1149 200 1183
rect 118 1115 142 1149
rect 176 1115 200 1149
rect 118 1081 200 1115
rect 118 1047 142 1081
rect 176 1047 200 1081
rect 118 1013 200 1047
rect 118 979 142 1013
rect 176 979 200 1013
rect 118 945 200 979
rect 118 911 142 945
rect 176 911 200 945
rect 118 877 200 911
rect 118 843 142 877
rect 176 843 200 877
rect 118 809 200 843
rect 118 775 142 809
rect 176 775 200 809
rect 118 741 200 775
rect 118 707 142 741
rect 176 707 200 741
rect 118 673 200 707
rect 118 639 142 673
rect 176 639 200 673
rect 118 605 200 639
rect 118 571 142 605
rect 176 571 200 605
rect 118 537 200 571
rect 118 503 142 537
rect 176 503 200 537
rect 1524 1387 1548 1421
rect 1582 1387 1606 1421
rect 1524 1353 1606 1387
rect 1524 1319 1548 1353
rect 1582 1319 1606 1353
rect 1524 1285 1606 1319
rect 1524 1251 1548 1285
rect 1582 1251 1606 1285
rect 1524 1217 1606 1251
rect 1524 1183 1548 1217
rect 1582 1183 1606 1217
rect 1524 1149 1606 1183
rect 1524 1115 1548 1149
rect 1582 1115 1606 1149
rect 1524 1081 1606 1115
rect 1524 1047 1548 1081
rect 1582 1047 1606 1081
rect 1524 1013 1606 1047
rect 1524 979 1548 1013
rect 1582 979 1606 1013
rect 1524 945 1606 979
rect 1524 911 1548 945
rect 1582 911 1606 945
rect 1524 877 1606 911
rect 1524 843 1548 877
rect 1582 843 1606 877
rect 1524 809 1606 843
rect 1524 775 1548 809
rect 1582 775 1606 809
rect 1524 741 1606 775
rect 1524 707 1548 741
rect 1582 707 1606 741
rect 1524 673 1606 707
rect 1524 639 1548 673
rect 1582 639 1606 673
rect 1524 605 1606 639
rect 1524 571 1548 605
rect 1582 571 1606 605
rect 1524 537 1606 571
rect 118 469 200 503
rect 118 435 142 469
rect 176 435 200 469
rect 118 401 200 435
rect 118 367 142 401
rect 176 367 200 401
rect 118 333 200 367
rect 118 299 142 333
rect 176 299 200 333
rect 118 265 200 299
rect 118 231 142 265
rect 176 231 200 265
rect 118 200 200 231
rect 1524 503 1548 537
rect 1582 503 1606 537
rect 1524 469 1606 503
rect 1524 435 1548 469
rect 1582 435 1606 469
rect 1524 401 1606 435
rect 1524 367 1548 401
rect 1582 367 1606 401
rect 1524 333 1606 367
rect 1524 299 1548 333
rect 1582 299 1606 333
rect 1524 265 1606 299
rect 1524 231 1548 265
rect 1582 231 1606 265
rect 1524 200 1606 231
rect 118 176 1606 200
rect 118 142 142 176
rect 176 142 233 176
rect 267 142 301 176
rect 335 142 369 176
rect 403 142 437 176
rect 471 142 505 176
rect 539 142 573 176
rect 607 142 641 176
rect 675 142 709 176
rect 743 142 777 176
rect 811 142 845 176
rect 879 142 913 176
rect 947 142 981 176
rect 1015 142 1049 176
rect 1083 142 1117 176
rect 1151 142 1185 176
rect 1219 142 1253 176
rect 1287 142 1321 176
rect 1355 142 1389 176
rect 1423 142 1457 176
rect 1491 142 1548 176
rect 1582 142 1606 176
rect 118 118 1606 142
<< psubdiffcont >>
rect 544 1346 578 1380
rect 641 1346 675 1380
rect 709 1346 743 1380
rect 777 1346 811 1380
rect 845 1346 879 1380
rect 913 1346 947 1380
rect 981 1346 1015 1380
rect 1049 1346 1083 1380
rect 1146 1346 1180 1380
rect 544 1251 578 1285
rect 544 1183 578 1217
rect 1146 1251 1180 1285
rect 1146 1183 1180 1217
rect 544 1115 578 1149
rect 544 1047 578 1081
rect 544 979 578 1013
rect 544 911 578 945
rect 544 843 578 877
rect 544 775 578 809
rect 1146 1115 1180 1149
rect 1146 1047 1180 1081
rect 1146 979 1180 1013
rect 1146 911 1180 945
rect 1146 843 1180 877
rect 1146 775 1180 809
rect 544 707 578 741
rect 544 639 578 673
rect 1146 707 1180 741
rect 1146 639 1180 673
rect 544 544 578 578
rect 641 544 675 578
rect 709 544 743 578
rect 777 544 811 578
rect 845 544 879 578
rect 913 544 947 578
rect 981 544 1015 578
rect 1049 544 1083 578
rect 1146 544 1180 578
<< nsubdiffcont >>
rect 142 1748 176 1782
rect 233 1748 267 1782
rect 301 1748 335 1782
rect 369 1748 403 1782
rect 437 1748 471 1782
rect 505 1748 539 1782
rect 573 1748 607 1782
rect 641 1748 675 1782
rect 709 1748 743 1782
rect 777 1748 811 1782
rect 845 1748 879 1782
rect 913 1748 947 1782
rect 981 1748 1015 1782
rect 1049 1748 1083 1782
rect 1117 1748 1151 1782
rect 1185 1748 1219 1782
rect 1253 1748 1287 1782
rect 1321 1748 1355 1782
rect 1389 1748 1423 1782
rect 1457 1748 1491 1782
rect 1548 1748 1582 1782
rect 142 1659 176 1693
rect 142 1591 176 1625
rect 142 1523 176 1557
rect 142 1455 176 1489
rect 142 1387 176 1421
rect 1548 1659 1582 1693
rect 1548 1591 1582 1625
rect 1548 1523 1582 1557
rect 1548 1455 1582 1489
rect 142 1319 176 1353
rect 142 1251 176 1285
rect 142 1183 176 1217
rect 142 1115 176 1149
rect 142 1047 176 1081
rect 142 979 176 1013
rect 142 911 176 945
rect 142 843 176 877
rect 142 775 176 809
rect 142 707 176 741
rect 142 639 176 673
rect 142 571 176 605
rect 142 503 176 537
rect 1548 1387 1582 1421
rect 1548 1319 1582 1353
rect 1548 1251 1582 1285
rect 1548 1183 1582 1217
rect 1548 1115 1582 1149
rect 1548 1047 1582 1081
rect 1548 979 1582 1013
rect 1548 911 1582 945
rect 1548 843 1582 877
rect 1548 775 1582 809
rect 1548 707 1582 741
rect 1548 639 1582 673
rect 1548 571 1582 605
rect 142 435 176 469
rect 142 367 176 401
rect 142 299 176 333
rect 142 231 176 265
rect 1548 503 1582 537
rect 1548 435 1582 469
rect 1548 367 1582 401
rect 1548 299 1582 333
rect 1548 231 1582 265
rect 142 142 176 176
rect 233 142 267 176
rect 301 142 335 176
rect 369 142 403 176
rect 437 142 471 176
rect 505 142 539 176
rect 573 142 607 176
rect 641 142 675 176
rect 709 142 743 176
rect 777 142 811 176
rect 845 142 879 176
rect 913 142 947 176
rect 981 142 1015 176
rect 1049 142 1083 176
rect 1117 142 1151 176
rect 1185 142 1219 176
rect 1253 142 1287 176
rect 1321 142 1355 176
rect 1389 142 1423 176
rect 1457 142 1491 176
rect 1548 142 1582 176
<< locali >>
rect 126 1782 1598 1798
rect 126 1748 142 1782
rect 176 1748 233 1782
rect 267 1748 301 1782
rect 339 1748 369 1782
rect 411 1748 437 1782
rect 483 1748 505 1782
rect 555 1748 573 1782
rect 627 1748 641 1782
rect 699 1748 709 1782
rect 771 1748 777 1782
rect 843 1748 845 1782
rect 879 1748 881 1782
rect 947 1748 953 1782
rect 1015 1748 1025 1782
rect 1083 1748 1097 1782
rect 1151 1748 1169 1782
rect 1219 1748 1241 1782
rect 1287 1748 1313 1782
rect 1355 1748 1385 1782
rect 1423 1748 1457 1782
rect 1491 1748 1548 1782
rect 1582 1748 1598 1782
rect 126 1732 1598 1748
rect 126 1699 192 1732
rect 126 1659 142 1699
rect 176 1659 192 1699
rect 126 1627 192 1659
rect 126 1591 142 1627
rect 176 1591 192 1627
rect 126 1557 192 1591
rect 126 1521 142 1557
rect 176 1521 192 1557
rect 126 1489 192 1521
rect 126 1449 142 1489
rect 176 1449 192 1489
rect 126 1421 192 1449
rect 126 1377 142 1421
rect 176 1377 192 1421
rect 1532 1699 1598 1732
rect 1532 1659 1548 1699
rect 1582 1659 1598 1699
rect 1532 1627 1598 1659
rect 1532 1591 1548 1627
rect 1582 1591 1598 1627
rect 1532 1557 1598 1591
rect 1532 1521 1548 1557
rect 1582 1521 1598 1557
rect 1532 1489 1598 1521
rect 1532 1449 1548 1489
rect 1582 1449 1598 1489
rect 1532 1421 1598 1449
rect 126 1353 192 1377
rect 126 1305 142 1353
rect 176 1305 192 1353
rect 126 1285 192 1305
rect 126 1233 142 1285
rect 176 1233 192 1285
rect 126 1217 192 1233
rect 126 1161 142 1217
rect 176 1161 192 1217
rect 126 1149 192 1161
rect 126 1089 142 1149
rect 176 1089 192 1149
rect 126 1081 192 1089
rect 126 1017 142 1081
rect 176 1017 192 1081
rect 126 1013 192 1017
rect 126 911 142 1013
rect 176 911 192 1013
rect 126 907 192 911
rect 126 843 142 907
rect 176 843 192 907
rect 126 835 192 843
rect 126 775 142 835
rect 176 775 192 835
rect 126 763 192 775
rect 126 707 142 763
rect 176 707 192 763
rect 126 691 192 707
rect 126 639 142 691
rect 176 639 192 691
rect 126 619 192 639
rect 126 571 142 619
rect 176 571 192 619
rect 126 547 192 571
rect 126 503 142 547
rect 176 503 192 547
rect 528 1380 1196 1396
rect 528 1346 544 1380
rect 578 1346 629 1380
rect 675 1346 701 1380
rect 743 1346 773 1380
rect 811 1346 845 1380
rect 879 1346 913 1380
rect 951 1346 981 1380
rect 1023 1346 1049 1380
rect 1095 1346 1146 1380
rect 1180 1346 1196 1380
rect 528 1330 1196 1346
rect 528 1303 594 1330
rect 528 1251 544 1303
rect 578 1251 594 1303
rect 528 1231 594 1251
rect 528 1183 544 1231
rect 578 1183 594 1231
rect 528 1159 594 1183
rect 1130 1303 1196 1330
rect 1130 1251 1146 1303
rect 1180 1251 1196 1303
rect 1130 1231 1196 1251
rect 1130 1183 1146 1231
rect 1180 1183 1196 1231
rect 528 1115 544 1159
rect 578 1115 594 1159
rect 528 1087 594 1115
rect 528 1047 544 1087
rect 578 1047 594 1087
rect 528 1015 594 1047
rect 528 979 544 1015
rect 578 979 594 1015
rect 528 945 594 979
rect 528 909 544 945
rect 578 909 594 945
rect 528 877 594 909
rect 528 837 544 877
rect 578 837 594 877
rect 528 809 594 837
rect 528 765 544 809
rect 578 765 594 809
rect 528 741 594 765
rect 761 1149 963 1165
rect 761 1123 777 1149
rect 947 1123 963 1149
rect 761 801 773 1123
rect 951 801 963 1123
rect 761 775 777 801
rect 947 775 963 801
rect 761 759 963 775
rect 1130 1159 1196 1183
rect 1130 1115 1146 1159
rect 1180 1115 1196 1159
rect 1130 1087 1196 1115
rect 1130 1047 1146 1087
rect 1180 1047 1196 1087
rect 1130 1015 1196 1047
rect 1130 979 1146 1015
rect 1180 979 1196 1015
rect 1130 945 1196 979
rect 1130 909 1146 945
rect 1180 909 1196 945
rect 1130 877 1196 909
rect 1130 837 1146 877
rect 1180 837 1196 877
rect 1130 809 1196 837
rect 1130 765 1146 809
rect 1180 765 1196 809
rect 528 693 544 741
rect 578 693 594 741
rect 528 673 594 693
rect 528 621 544 673
rect 578 621 594 673
rect 528 594 594 621
rect 1130 741 1196 765
rect 1130 693 1146 741
rect 1180 693 1196 741
rect 1130 673 1196 693
rect 1130 621 1146 673
rect 1180 621 1196 673
rect 1130 594 1196 621
rect 528 578 1196 594
rect 528 544 544 578
rect 578 544 629 578
rect 675 544 701 578
rect 743 544 773 578
rect 811 544 845 578
rect 879 544 913 578
rect 951 544 981 578
rect 1023 544 1049 578
rect 1095 544 1146 578
rect 1180 544 1196 578
rect 528 528 1196 544
rect 1532 1377 1548 1421
rect 1582 1377 1598 1421
rect 1532 1353 1598 1377
rect 1532 1305 1548 1353
rect 1582 1305 1598 1353
rect 1532 1285 1598 1305
rect 1532 1233 1548 1285
rect 1582 1233 1598 1285
rect 1532 1217 1598 1233
rect 1532 1161 1548 1217
rect 1582 1161 1598 1217
rect 1532 1149 1598 1161
rect 1532 1089 1548 1149
rect 1582 1089 1598 1149
rect 1532 1081 1598 1089
rect 1532 1017 1548 1081
rect 1582 1017 1598 1081
rect 1532 1013 1598 1017
rect 1532 911 1548 1013
rect 1582 911 1598 1013
rect 1532 907 1598 911
rect 1532 843 1548 907
rect 1582 843 1598 907
rect 1532 835 1598 843
rect 1532 775 1548 835
rect 1582 775 1598 835
rect 1532 763 1598 775
rect 1532 707 1548 763
rect 1582 707 1598 763
rect 1532 691 1598 707
rect 1532 639 1548 691
rect 1582 639 1598 691
rect 1532 619 1598 639
rect 1532 571 1548 619
rect 1582 571 1598 619
rect 1532 547 1598 571
rect 126 475 192 503
rect 126 435 142 475
rect 176 435 192 475
rect 126 403 192 435
rect 126 367 142 403
rect 176 367 192 403
rect 126 333 192 367
rect 126 297 142 333
rect 176 297 192 333
rect 126 265 192 297
rect 126 225 142 265
rect 176 225 192 265
rect 126 192 192 225
rect 1532 503 1548 547
rect 1582 503 1598 547
rect 1532 475 1598 503
rect 1532 435 1548 475
rect 1582 435 1598 475
rect 1532 403 1598 435
rect 1532 367 1548 403
rect 1582 367 1598 403
rect 1532 333 1598 367
rect 1532 297 1548 333
rect 1582 297 1598 333
rect 1532 265 1598 297
rect 1532 225 1548 265
rect 1582 225 1598 265
rect 1532 192 1598 225
rect 126 176 1598 192
rect 126 142 142 176
rect 176 142 233 176
rect 267 142 301 176
rect 339 142 369 176
rect 411 142 437 176
rect 483 142 505 176
rect 555 142 573 176
rect 627 142 641 176
rect 699 142 709 176
rect 771 142 777 176
rect 843 142 845 176
rect 879 142 881 176
rect 947 142 953 176
rect 1015 142 1025 176
rect 1083 142 1097 176
rect 1151 142 1169 176
rect 1219 142 1241 176
rect 1287 142 1313 176
rect 1355 142 1385 176
rect 1423 142 1457 176
rect 1491 142 1548 176
rect 1582 142 1598 176
rect 126 126 1598 142
<< viali >>
rect 142 1748 176 1782
rect 233 1748 267 1782
rect 305 1748 335 1782
rect 335 1748 339 1782
rect 377 1748 403 1782
rect 403 1748 411 1782
rect 449 1748 471 1782
rect 471 1748 483 1782
rect 521 1748 539 1782
rect 539 1748 555 1782
rect 593 1748 607 1782
rect 607 1748 627 1782
rect 665 1748 675 1782
rect 675 1748 699 1782
rect 737 1748 743 1782
rect 743 1748 771 1782
rect 809 1748 811 1782
rect 811 1748 843 1782
rect 881 1748 913 1782
rect 913 1748 915 1782
rect 953 1748 981 1782
rect 981 1748 987 1782
rect 1025 1748 1049 1782
rect 1049 1748 1059 1782
rect 1097 1748 1117 1782
rect 1117 1748 1131 1782
rect 1169 1748 1185 1782
rect 1185 1748 1203 1782
rect 1241 1748 1253 1782
rect 1253 1748 1275 1782
rect 1313 1748 1321 1782
rect 1321 1748 1347 1782
rect 1385 1748 1389 1782
rect 1389 1748 1419 1782
rect 1457 1748 1491 1782
rect 1548 1748 1582 1782
rect 142 1693 176 1699
rect 142 1665 176 1693
rect 142 1625 176 1627
rect 142 1593 176 1625
rect 142 1523 176 1555
rect 142 1521 176 1523
rect 142 1455 176 1483
rect 142 1449 176 1455
rect 142 1387 176 1411
rect 142 1377 176 1387
rect 1548 1693 1582 1699
rect 1548 1665 1582 1693
rect 1548 1625 1582 1627
rect 1548 1593 1582 1625
rect 1548 1523 1582 1555
rect 1548 1521 1582 1523
rect 1548 1455 1582 1483
rect 1548 1449 1582 1455
rect 142 1319 176 1339
rect 142 1305 176 1319
rect 142 1251 176 1267
rect 142 1233 176 1251
rect 142 1183 176 1195
rect 142 1161 176 1183
rect 142 1115 176 1123
rect 142 1089 176 1115
rect 142 1047 176 1051
rect 142 1017 176 1047
rect 142 945 176 979
rect 142 877 176 907
rect 142 873 176 877
rect 142 809 176 835
rect 142 801 176 809
rect 142 741 176 763
rect 142 729 176 741
rect 142 673 176 691
rect 142 657 176 673
rect 142 605 176 619
rect 142 585 176 605
rect 142 537 176 547
rect 142 513 176 537
rect 544 1346 578 1380
rect 629 1346 641 1380
rect 641 1346 663 1380
rect 701 1346 709 1380
rect 709 1346 735 1380
rect 773 1346 777 1380
rect 777 1346 807 1380
rect 845 1346 879 1380
rect 917 1346 947 1380
rect 947 1346 951 1380
rect 989 1346 1015 1380
rect 1015 1346 1023 1380
rect 1061 1346 1083 1380
rect 1083 1346 1095 1380
rect 1146 1346 1180 1380
rect 544 1285 578 1303
rect 544 1269 578 1285
rect 544 1217 578 1231
rect 544 1197 578 1217
rect 1146 1285 1180 1303
rect 1146 1269 1180 1285
rect 1146 1217 1180 1231
rect 1146 1197 1180 1217
rect 544 1149 578 1159
rect 544 1125 578 1149
rect 544 1081 578 1087
rect 544 1053 578 1081
rect 544 1013 578 1015
rect 544 981 578 1013
rect 544 911 578 943
rect 544 909 578 911
rect 544 843 578 871
rect 544 837 578 843
rect 544 775 578 799
rect 544 765 578 775
rect 773 801 777 1123
rect 777 801 947 1123
rect 947 801 951 1123
rect 1146 1149 1180 1159
rect 1146 1125 1180 1149
rect 1146 1081 1180 1087
rect 1146 1053 1180 1081
rect 1146 1013 1180 1015
rect 1146 981 1180 1013
rect 1146 911 1180 943
rect 1146 909 1180 911
rect 1146 843 1180 871
rect 1146 837 1180 843
rect 1146 775 1180 799
rect 1146 765 1180 775
rect 544 707 578 727
rect 544 693 578 707
rect 544 639 578 655
rect 544 621 578 639
rect 1146 707 1180 727
rect 1146 693 1180 707
rect 1146 639 1180 655
rect 1146 621 1180 639
rect 544 544 578 578
rect 629 544 641 578
rect 641 544 663 578
rect 701 544 709 578
rect 709 544 735 578
rect 773 544 777 578
rect 777 544 807 578
rect 845 544 879 578
rect 917 544 947 578
rect 947 544 951 578
rect 989 544 1015 578
rect 1015 544 1023 578
rect 1061 544 1083 578
rect 1083 544 1095 578
rect 1146 544 1180 578
rect 1548 1387 1582 1411
rect 1548 1377 1582 1387
rect 1548 1319 1582 1339
rect 1548 1305 1582 1319
rect 1548 1251 1582 1267
rect 1548 1233 1582 1251
rect 1548 1183 1582 1195
rect 1548 1161 1582 1183
rect 1548 1115 1582 1123
rect 1548 1089 1582 1115
rect 1548 1047 1582 1051
rect 1548 1017 1582 1047
rect 1548 945 1582 979
rect 1548 877 1582 907
rect 1548 873 1582 877
rect 1548 809 1582 835
rect 1548 801 1582 809
rect 1548 741 1582 763
rect 1548 729 1582 741
rect 1548 673 1582 691
rect 1548 657 1582 673
rect 1548 605 1582 619
rect 1548 585 1582 605
rect 142 469 176 475
rect 142 441 176 469
rect 142 401 176 403
rect 142 369 176 401
rect 142 299 176 331
rect 142 297 176 299
rect 142 231 176 259
rect 142 225 176 231
rect 1548 537 1582 547
rect 1548 513 1582 537
rect 1548 469 1582 475
rect 1548 441 1582 469
rect 1548 401 1582 403
rect 1548 369 1582 401
rect 1548 299 1582 331
rect 1548 297 1582 299
rect 1548 231 1582 259
rect 1548 225 1582 231
rect 142 142 176 176
rect 233 142 267 176
rect 305 142 335 176
rect 335 142 339 176
rect 377 142 403 176
rect 403 142 411 176
rect 449 142 471 176
rect 471 142 483 176
rect 521 142 539 176
rect 539 142 555 176
rect 593 142 607 176
rect 607 142 627 176
rect 665 142 675 176
rect 675 142 699 176
rect 737 142 743 176
rect 743 142 771 176
rect 809 142 811 176
rect 811 142 843 176
rect 881 142 913 176
rect 913 142 915 176
rect 953 142 981 176
rect 981 142 987 176
rect 1025 142 1049 176
rect 1049 142 1059 176
rect 1097 142 1117 176
rect 1117 142 1131 176
rect 1169 142 1185 176
rect 1185 142 1203 176
rect 1241 142 1253 176
rect 1253 142 1275 176
rect 1313 142 1321 176
rect 1321 142 1347 176
rect 1385 142 1389 176
rect 1389 142 1419 176
rect 1457 142 1491 176
rect 1548 142 1582 176
<< metal1 >>
rect 130 1782 1594 1794
rect 130 1748 142 1782
rect 176 1748 233 1782
rect 267 1748 305 1782
rect 339 1748 377 1782
rect 411 1748 449 1782
rect 483 1748 521 1782
rect 555 1748 593 1782
rect 627 1748 665 1782
rect 699 1748 737 1782
rect 771 1748 809 1782
rect 843 1748 881 1782
rect 915 1748 953 1782
rect 987 1748 1025 1782
rect 1059 1748 1097 1782
rect 1131 1748 1169 1782
rect 1203 1748 1241 1782
rect 1275 1748 1313 1782
rect 1347 1748 1385 1782
rect 1419 1748 1457 1782
rect 1491 1748 1548 1782
rect 1582 1748 1594 1782
rect 130 1736 1594 1748
rect 130 1699 188 1736
rect 130 1665 142 1699
rect 176 1665 188 1699
rect 130 1627 188 1665
rect 130 1593 142 1627
rect 176 1593 188 1627
rect 130 1555 188 1593
rect 130 1521 142 1555
rect 176 1521 188 1555
rect 130 1483 188 1521
rect 130 1449 142 1483
rect 176 1449 188 1483
rect 130 1411 188 1449
rect 130 1377 142 1411
rect 176 1377 188 1411
rect 1536 1699 1594 1736
rect 1536 1665 1548 1699
rect 1582 1665 1594 1699
rect 1536 1627 1594 1665
rect 1536 1593 1548 1627
rect 1582 1593 1594 1627
rect 1536 1555 1594 1593
rect 1536 1521 1548 1555
rect 1582 1521 1594 1555
rect 1536 1483 1594 1521
rect 1536 1449 1548 1483
rect 1582 1449 1594 1483
rect 1536 1411 1594 1449
rect 130 1339 188 1377
rect 130 1305 142 1339
rect 176 1305 188 1339
rect 130 1267 188 1305
rect 130 1233 142 1267
rect 176 1233 188 1267
rect 130 1195 188 1233
rect 130 1161 142 1195
rect 176 1161 188 1195
rect 130 1123 188 1161
rect 130 1089 142 1123
rect 176 1089 188 1123
rect 130 1051 188 1089
rect 130 1017 142 1051
rect 176 1017 188 1051
rect 130 979 188 1017
rect 130 945 142 979
rect 176 945 188 979
rect 130 907 188 945
rect 130 873 142 907
rect 176 873 188 907
rect 130 835 188 873
rect 130 801 142 835
rect 176 801 188 835
rect 130 763 188 801
rect 130 729 142 763
rect 176 729 188 763
rect 130 691 188 729
rect 130 657 142 691
rect 176 657 188 691
rect 130 619 188 657
rect 130 585 142 619
rect 176 585 188 619
rect 130 547 188 585
rect 130 513 142 547
rect 176 513 188 547
rect 532 1380 1192 1392
rect 532 1346 544 1380
rect 578 1346 629 1380
rect 663 1346 701 1380
rect 735 1346 773 1380
rect 807 1346 845 1380
rect 879 1346 917 1380
rect 951 1346 989 1380
rect 1023 1346 1061 1380
rect 1095 1346 1146 1380
rect 1180 1346 1192 1380
rect 532 1334 1192 1346
rect 532 1303 590 1334
rect 532 1269 544 1303
rect 578 1269 590 1303
rect 532 1231 590 1269
rect 532 1197 544 1231
rect 578 1197 590 1231
rect 532 1159 590 1197
rect 532 1125 544 1159
rect 578 1125 590 1159
rect 1134 1303 1192 1334
rect 1134 1269 1146 1303
rect 1180 1269 1192 1303
rect 1134 1231 1192 1269
rect 1134 1197 1146 1231
rect 1180 1197 1192 1231
rect 1134 1159 1192 1197
rect 532 1087 590 1125
rect 532 1053 544 1087
rect 578 1053 590 1087
rect 532 1015 590 1053
rect 532 981 544 1015
rect 578 981 590 1015
rect 532 943 590 981
rect 532 909 544 943
rect 578 909 590 943
rect 532 871 590 909
rect 532 837 544 871
rect 578 837 590 871
rect 532 799 590 837
rect 532 765 544 799
rect 578 765 590 799
rect 761 1123 963 1135
rect 761 801 773 1123
rect 951 801 963 1123
rect 761 789 963 801
rect 1134 1125 1146 1159
rect 1180 1125 1192 1159
rect 1134 1087 1192 1125
rect 1134 1053 1146 1087
rect 1180 1053 1192 1087
rect 1134 1015 1192 1053
rect 1134 981 1146 1015
rect 1180 981 1192 1015
rect 1134 943 1192 981
rect 1134 909 1146 943
rect 1180 909 1192 943
rect 1134 871 1192 909
rect 1134 837 1146 871
rect 1180 837 1192 871
rect 1134 799 1192 837
rect 532 727 590 765
rect 532 693 544 727
rect 578 693 590 727
rect 532 655 590 693
rect 532 621 544 655
rect 578 621 590 655
rect 532 590 590 621
rect 1134 765 1146 799
rect 1180 765 1192 799
rect 1134 727 1192 765
rect 1134 693 1146 727
rect 1180 693 1192 727
rect 1134 655 1192 693
rect 1134 621 1146 655
rect 1180 621 1192 655
rect 1134 590 1192 621
rect 532 578 1192 590
rect 532 544 544 578
rect 578 544 629 578
rect 663 544 701 578
rect 735 544 773 578
rect 807 544 845 578
rect 879 544 917 578
rect 951 544 989 578
rect 1023 544 1061 578
rect 1095 544 1146 578
rect 1180 544 1192 578
rect 532 532 1192 544
rect 1536 1377 1548 1411
rect 1582 1377 1594 1411
rect 1536 1339 1594 1377
rect 1536 1305 1548 1339
rect 1582 1305 1594 1339
rect 1536 1267 1594 1305
rect 1536 1233 1548 1267
rect 1582 1233 1594 1267
rect 1536 1195 1594 1233
rect 1536 1161 1548 1195
rect 1582 1161 1594 1195
rect 1536 1123 1594 1161
rect 1536 1089 1548 1123
rect 1582 1089 1594 1123
rect 1536 1051 1594 1089
rect 1536 1017 1548 1051
rect 1582 1017 1594 1051
rect 1536 979 1594 1017
rect 1536 945 1548 979
rect 1582 945 1594 979
rect 1536 907 1594 945
rect 1536 873 1548 907
rect 1582 873 1594 907
rect 1536 835 1594 873
rect 1536 801 1548 835
rect 1582 801 1594 835
rect 1536 763 1594 801
rect 1536 729 1548 763
rect 1582 729 1594 763
rect 1536 691 1594 729
rect 1536 657 1548 691
rect 1582 657 1594 691
rect 1536 619 1594 657
rect 1536 585 1548 619
rect 1582 585 1594 619
rect 1536 547 1594 585
rect 130 475 188 513
rect 130 441 142 475
rect 176 441 188 475
rect 130 403 188 441
rect 130 369 142 403
rect 176 369 188 403
rect 130 331 188 369
rect 130 297 142 331
rect 176 297 188 331
rect 130 259 188 297
rect 130 225 142 259
rect 176 225 188 259
rect 130 188 188 225
rect 1536 513 1548 547
rect 1582 513 1594 547
rect 1536 475 1594 513
rect 1536 441 1548 475
rect 1582 441 1594 475
rect 1536 403 1594 441
rect 1536 369 1548 403
rect 1582 369 1594 403
rect 1536 331 1594 369
rect 1536 297 1548 331
rect 1582 297 1594 331
rect 1536 259 1594 297
rect 1536 225 1548 259
rect 1582 225 1594 259
rect 1536 188 1594 225
rect 130 176 1594 188
rect 130 142 142 176
rect 176 142 233 176
rect 267 142 305 176
rect 339 142 377 176
rect 411 142 449 176
rect 483 142 521 176
rect 555 142 593 176
rect 627 142 665 176
rect 699 142 737 176
rect 771 142 809 176
rect 843 142 881 176
rect 915 142 953 176
rect 987 142 1025 176
rect 1059 142 1097 176
rect 1131 142 1169 176
rect 1203 142 1241 176
rect 1275 142 1313 176
rect 1347 142 1385 176
rect 1419 142 1457 176
rect 1491 142 1548 176
rect 1582 142 1594 176
rect 130 130 1594 142
<< properties >>
string gencell sky130_fd_pr__rf_npn_05v5_W1p00L2p00
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 9104402
string GDS_START 9080134
string parameter m=1
string library sky130
string path 4.500 9.000 4.500 43.600 38.600 43.600 38.600 4.500 0.000 4.500 
<< end >>
