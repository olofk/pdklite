magic
tech sky130A
magscale 1 2
timestamp 1619729571
<< checkpaint >>
rect -1298 -1308 2494 1852
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 97 47 127 177
rect 181 47 211 177
rect 369 47 399 177
rect 453 47 483 177
rect 537 47 567 177
rect 621 47 651 177
rect 809 47 839 177
rect 893 47 923 177
rect 977 47 1007 177
rect 1061 47 1091 177
<< scpmoshvt >>
rect 201 297 231 497
rect 285 297 315 497
rect 369 297 399 497
rect 453 297 483 497
rect 537 297 567 497
rect 621 297 651 497
rect 709 297 739 497
rect 893 297 923 497
rect 977 297 1007 497
rect 1061 297 1091 497
<< ndiff >>
rect 45 93 97 177
rect 45 59 53 93
rect 87 59 97 93
rect 45 47 97 59
rect 127 101 181 177
rect 127 67 137 101
rect 171 67 181 101
rect 127 47 181 67
rect 211 93 263 177
rect 211 59 221 93
rect 255 59 263 93
rect 211 47 263 59
rect 317 93 369 177
rect 317 59 325 93
rect 359 59 369 93
rect 317 47 369 59
rect 399 163 453 177
rect 399 129 409 163
rect 443 129 453 163
rect 399 47 453 129
rect 483 147 537 177
rect 483 113 493 147
rect 527 113 537 147
rect 483 47 537 113
rect 567 93 621 177
rect 567 59 577 93
rect 611 59 621 93
rect 567 47 621 59
rect 651 163 703 177
rect 651 129 661 163
rect 695 129 703 163
rect 651 47 703 129
rect 757 163 809 177
rect 757 129 765 163
rect 799 129 809 163
rect 757 47 809 129
rect 839 93 893 177
rect 839 59 849 93
rect 883 59 893 93
rect 839 47 893 59
rect 923 163 977 177
rect 923 129 933 163
rect 967 129 977 163
rect 923 47 977 129
rect 1007 93 1061 177
rect 1007 59 1017 93
rect 1051 59 1061 93
rect 1007 47 1061 59
rect 1091 101 1143 177
rect 1091 67 1101 101
rect 1135 67 1143 101
rect 1091 47 1143 67
<< pdiff >>
rect 149 477 201 497
rect 149 443 157 477
rect 191 443 201 477
rect 149 409 201 443
rect 149 375 157 409
rect 191 375 201 409
rect 149 297 201 375
rect 231 425 285 497
rect 231 391 241 425
rect 275 391 285 425
rect 231 357 285 391
rect 231 323 241 357
rect 275 323 285 357
rect 231 297 285 323
rect 315 477 369 497
rect 315 443 325 477
rect 359 443 369 477
rect 315 409 369 443
rect 315 375 325 409
rect 359 375 369 409
rect 315 297 369 375
rect 399 485 453 497
rect 399 451 409 485
rect 443 451 453 485
rect 399 417 453 451
rect 399 383 409 417
rect 443 383 453 417
rect 399 297 453 383
rect 483 477 537 497
rect 483 443 493 477
rect 527 443 537 477
rect 483 409 537 443
rect 483 375 493 409
rect 527 375 537 409
rect 483 297 537 375
rect 567 485 621 497
rect 567 451 577 485
rect 611 451 621 485
rect 567 417 621 451
rect 567 383 577 417
rect 611 383 621 417
rect 567 297 621 383
rect 651 477 709 497
rect 651 443 665 477
rect 699 443 709 477
rect 651 409 709 443
rect 651 375 665 409
rect 699 375 709 409
rect 651 297 709 375
rect 739 485 893 497
rect 739 383 767 485
rect 869 383 893 485
rect 739 297 893 383
rect 923 477 977 497
rect 923 443 933 477
rect 967 443 977 477
rect 923 409 977 443
rect 923 375 933 409
rect 967 375 977 409
rect 923 297 977 375
rect 1007 485 1061 497
rect 1007 451 1017 485
rect 1051 451 1061 485
rect 1007 417 1061 451
rect 1007 383 1017 417
rect 1051 383 1061 417
rect 1007 297 1061 383
rect 1091 477 1143 497
rect 1091 443 1101 477
rect 1135 443 1143 477
rect 1091 409 1143 443
rect 1091 375 1101 409
rect 1135 375 1143 409
rect 1091 297 1143 375
<< ndiffc >>
rect 53 59 87 93
rect 137 67 171 101
rect 221 59 255 93
rect 325 59 359 93
rect 409 129 443 163
rect 493 113 527 147
rect 577 59 611 93
rect 661 129 695 163
rect 765 129 799 163
rect 849 59 883 93
rect 933 129 967 163
rect 1017 59 1051 93
rect 1101 67 1135 101
<< pdiffc >>
rect 157 443 191 477
rect 157 375 191 409
rect 241 391 275 425
rect 241 323 275 357
rect 325 443 359 477
rect 325 375 359 409
rect 409 451 443 485
rect 409 383 443 417
rect 493 443 527 477
rect 493 375 527 409
rect 577 451 611 485
rect 577 383 611 417
rect 665 443 699 477
rect 665 375 699 409
rect 767 383 869 485
rect 933 443 967 477
rect 933 375 967 409
rect 1017 451 1051 485
rect 1017 383 1051 417
rect 1101 443 1135 477
rect 1101 375 1135 409
<< poly >>
rect 201 497 231 523
rect 285 497 315 523
rect 369 497 399 523
rect 453 497 483 523
rect 537 497 567 523
rect 621 497 651 523
rect 709 497 739 523
rect 893 497 923 523
rect 977 497 1007 523
rect 1061 497 1091 523
rect 201 265 231 297
rect 285 265 315 297
rect 97 249 315 265
rect 369 265 399 297
rect 453 265 483 297
rect 369 259 483 265
rect 537 259 567 297
rect 621 259 651 297
rect 709 259 739 297
rect 893 259 923 297
rect 977 259 1007 297
rect 1061 261 1091 297
rect 1061 259 1175 261
rect 97 215 125 249
rect 159 215 193 249
rect 227 215 261 249
rect 295 215 315 249
rect 97 199 315 215
rect 357 249 491 259
rect 357 215 373 249
rect 407 215 441 249
rect 475 215 491 249
rect 357 205 491 215
rect 533 249 667 259
rect 533 215 549 249
rect 583 215 617 249
rect 651 215 667 249
rect 533 205 667 215
rect 709 249 923 259
rect 709 215 725 249
rect 759 215 797 249
rect 831 215 865 249
rect 899 215 923 249
rect 709 205 923 215
rect 965 249 1175 259
rect 965 215 989 249
rect 1023 215 1057 249
rect 1091 215 1125 249
rect 1159 215 1175 249
rect 965 205 1175 215
rect 369 199 483 205
rect 97 177 127 199
rect 181 177 211 199
rect 369 177 399 199
rect 453 177 483 199
rect 537 177 567 205
rect 621 177 651 205
rect 809 177 839 205
rect 893 177 923 205
rect 977 177 1007 205
rect 1061 203 1175 205
rect 1061 177 1091 203
rect 97 21 127 47
rect 181 21 211 47
rect 369 21 399 47
rect 453 21 483 47
rect 537 21 567 47
rect 621 21 651 47
rect 809 21 839 47
rect 893 21 923 47
rect 977 21 1007 47
rect 1061 21 1091 47
<< polycont >>
rect 125 215 159 249
rect 193 215 227 249
rect 261 215 295 249
rect 373 215 407 249
rect 441 215 475 249
rect 549 215 583 249
rect 617 215 651 249
rect 725 215 759 249
rect 797 215 831 249
rect 865 215 899 249
rect 989 215 1023 249
rect 1057 215 1091 249
rect 1125 215 1159 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 157 477 359 493
rect 191 459 325 477
rect 157 409 191 443
rect 157 359 191 375
rect 225 391 241 425
rect 275 391 291 425
rect 225 357 291 391
rect 225 325 241 357
rect 29 323 241 325
rect 275 323 291 357
rect 29 291 291 323
rect 325 409 359 443
rect 393 485 459 527
rect 393 451 409 485
rect 443 451 459 485
rect 393 417 459 451
rect 393 383 409 417
rect 443 383 459 417
rect 493 477 527 493
rect 493 409 527 443
rect 325 341 359 375
rect 561 485 627 527
rect 561 451 577 485
rect 611 451 627 485
rect 561 417 627 451
rect 561 383 577 417
rect 611 383 627 417
rect 665 477 699 493
rect 665 409 699 443
rect 493 341 527 375
rect 751 485 885 527
rect 751 383 767 485
rect 869 383 885 485
rect 933 477 967 493
rect 933 409 967 443
rect 665 341 699 375
rect 1001 485 1067 527
rect 1001 451 1017 485
rect 1051 451 1067 485
rect 1001 417 1067 451
rect 1001 383 1017 417
rect 1051 383 1067 417
rect 1101 477 1135 493
rect 1101 409 1135 443
rect 933 341 967 375
rect 1101 341 1135 375
rect 325 307 1152 341
rect 29 163 63 291
rect 109 249 311 256
rect 109 215 125 249
rect 159 215 193 249
rect 227 215 261 249
rect 295 215 311 249
rect 357 249 491 259
rect 357 215 373 249
rect 407 215 441 249
rect 475 215 491 249
rect 533 249 673 257
rect 533 215 549 249
rect 583 215 617 249
rect 651 215 673 249
rect 709 249 915 259
rect 709 215 725 249
rect 759 215 797 249
rect 831 215 865 249
rect 899 215 915 249
rect 951 249 1179 259
rect 951 215 989 249
rect 1023 215 1057 249
rect 1091 215 1125 249
rect 1159 215 1179 249
rect 29 129 409 163
rect 443 129 459 163
rect 493 147 661 163
rect 137 101 171 129
rect 37 59 53 93
rect 87 59 103 93
rect 37 17 103 59
rect 527 129 661 147
rect 695 129 711 163
rect 749 129 765 163
rect 799 129 933 163
rect 967 129 1135 163
rect 493 93 527 113
rect 1101 101 1135 129
rect 137 51 171 67
rect 205 59 221 93
rect 255 59 275 93
rect 309 59 325 93
rect 359 59 527 93
rect 561 59 577 93
rect 611 59 849 93
rect 883 59 899 93
rect 1001 59 1017 93
rect 1051 59 1067 93
rect 205 17 275 59
rect 1001 17 1067 59
rect 1101 51 1135 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 1133 221 1167 255 0 FreeSans 200 0 0 0 A4
port 4 nsew signal input
flabel locali s 953 221 987 255 0 FreeSans 200 0 0 0 A4
port 4 nsew signal input
flabel locali s 769 221 803 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1041 221 1075 255 0 FreeSans 200 0 0 0 A4
port 4 nsew signal input
flabel locali s 861 221 895 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 B1
port 5 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 B1
port 5 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 29 153 63 187 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 a41oi_2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 651636
string GDS_START 641566
string path 0.000 13.600 29.900 13.600 
<< end >>
