magic
tech sky130A
magscale 1 2
timestamp 1640697850
<< dnwell >>
rect -1000 1958 0 7825
<< poly >>
rect 149 9434 336 9467
rect 149 9400 166 9434
rect 200 9400 234 9434
rect 268 9400 302 9434
rect 149 9367 336 9400
rect 2376 9434 2563 9467
rect 2410 9400 2444 9434
rect 2478 9400 2512 9434
rect 2546 9400 2563 9434
rect 2376 9367 2563 9400
<< polycont >>
rect 166 9400 200 9434
rect 234 9400 268 9434
rect 302 9400 336 9434
rect 2376 9400 2410 9434
rect 2444 9400 2478 9434
rect 2512 9400 2546 9434
<< npolyres >>
rect 336 9367 2376 9467
<< locali >>
rect 150 9440 352 9450
rect 150 9434 353 9440
rect 150 9400 163 9434
rect 200 9400 234 9434
rect 269 9400 302 9434
rect 341 9400 353 9434
rect 150 9394 353 9400
rect 2359 9434 2562 9508
rect 2359 9400 2371 9434
rect 2410 9400 2443 9434
rect 2478 9400 2512 9434
rect 2549 9400 2562 9434
rect 2359 9394 2562 9400
rect 150 9384 352 9394
rect 2360 9384 2562 9394
rect 688 3618 702 7256
rect 14252 3618 14266 7256
rect 301 2962 12495 2978
<< viali >>
rect 163 9400 166 9434
rect 166 9400 197 9434
rect 235 9400 268 9434
rect 268 9400 269 9434
rect 307 9400 336 9434
rect 336 9400 341 9434
rect 2371 9400 2376 9434
rect 2376 9400 2405 9434
rect 2443 9400 2444 9434
rect 2444 9400 2477 9434
rect 2515 9400 2546 9434
rect 2546 9400 2549 9434
<< metal1 >>
rect 321 9512 373 9520
tri 287 9440 321 9474 se
rect 321 9448 373 9460
rect 150 9434 321 9440
rect 150 9400 163 9434
rect 197 9400 235 9434
rect 269 9400 307 9434
rect 150 9396 321 9400
rect 150 9394 373 9396
tri 317 9390 321 9394 ne
rect 321 9390 373 9394
rect 2359 9434 2562 9487
rect 2359 9400 2371 9434
rect 2405 9400 2443 9434
rect 2477 9400 2515 9434
rect 2549 9400 2562 9434
rect 2359 9357 2562 9400
rect 785 4021 1705 4028
rect 785 3969 791 4021
rect 843 3969 857 4021
rect 909 3969 1705 4021
rect 785 3957 1705 3969
rect 785 3905 791 3957
rect 843 3905 857 3957
rect 909 3905 1705 3957
rect 785 3898 1705 3905
rect 2135 3976 2141 4028
rect 2193 3976 2207 4028
rect 2259 3976 2265 4028
rect 2135 3950 2265 3976
rect 2135 3898 2141 3950
rect 2193 3898 2207 3950
rect 2259 3898 2265 3950
rect 2697 4021 2827 4028
rect 2697 3969 2703 4021
rect 2755 3969 2769 4021
rect 2821 3969 2827 4021
rect 2697 3957 2827 3969
rect 2697 3905 2703 3957
rect 2755 3905 2769 3957
rect 2821 3905 2827 3957
rect 2697 3898 2827 3905
rect 3257 3898 3757 4028
rect 3810 4021 4189 4028
rect 3810 3969 3816 4021
rect 3868 3969 3895 4021
rect 3947 3969 3974 4021
rect 4026 3969 4053 4021
rect 4105 3969 4131 4021
rect 4183 3969 4189 4021
rect 3810 3957 4189 3969
rect 3810 3905 3816 3957
rect 3868 3905 3895 3957
rect 3947 3905 3974 3957
rect 4026 3905 4053 3957
rect 4105 3905 4131 3957
rect 4183 3905 4189 3957
rect 3810 3898 4189 3905
rect 4249 3898 4681 4028
rect 4686 3898 5678 4028
rect 6103 3976 6109 4028
rect 6161 3976 6174 4028
rect 6226 3976 6239 4028
rect 6291 3976 6304 4028
rect 6356 3976 6368 4028
rect 6420 3976 6432 4028
rect 6484 3976 6496 4028
rect 6548 3976 6560 4028
rect 6612 3976 6624 4028
rect 6676 3976 6688 4028
rect 6740 3976 6752 4028
rect 6804 3976 7095 4028
rect 6103 3956 7095 3976
rect 6103 3904 6109 3956
rect 6161 3904 6174 3956
rect 6226 3904 6239 3956
rect 6291 3904 6304 3956
rect 6356 3904 6368 3956
rect 6420 3904 6432 3956
rect 6484 3904 6496 3956
rect 6548 3904 6560 3956
rect 6612 3904 6624 3956
rect 6676 3904 6688 3956
rect 6740 3904 6752 3956
rect 6804 3904 7095 3956
rect 6103 3898 7095 3904
rect 7657 3976 7663 4028
rect 7715 3976 7729 4028
rect 7781 3976 7787 4028
rect 7657 3950 7787 3976
rect 7657 3898 7663 3950
rect 7715 3898 7729 3950
rect 7781 3898 7787 3950
rect 8232 3976 8595 4028
rect 8647 3976 8660 4028
rect 8712 3976 8724 4028
rect 8776 3976 8788 4028
rect 8840 3976 9202 4028
rect 8232 3954 9202 3976
rect 8232 3902 8595 3954
rect 8647 3902 8660 3954
rect 8712 3902 8724 3954
rect 8776 3902 8788 3954
rect 8840 3902 9202 3954
rect 8232 3898 9202 3902
rect 9769 3986 10750 4028
rect 9769 3934 10220 3986
rect 10272 3934 10286 3986
rect 10338 3934 10352 3986
rect 10404 3934 10418 3986
rect 10470 3934 10483 3986
rect 10535 3934 10548 3986
rect 10600 3934 10613 3986
rect 10665 3934 10678 3986
rect 10730 3934 10750 3986
rect 9769 3898 10750 3934
rect 11193 3987 12185 4028
rect 11193 3935 11631 3987
rect 11683 3935 11696 3987
rect 11748 3935 11761 3987
rect 11813 3935 11826 3987
rect 11878 3935 11891 3987
rect 11943 3935 11956 3987
rect 12008 3935 12021 3987
rect 12073 3935 12185 3987
rect 11193 3898 12185 3935
rect 12747 3976 13053 4028
rect 13105 3976 13120 4028
rect 13172 3976 13187 4028
rect 13239 3976 13254 4028
rect 13306 3976 13321 4028
rect 13373 3976 13388 4028
rect 13440 3976 13455 4028
rect 13507 3976 14039 4028
rect 12747 3950 14039 3976
rect 12747 3898 13053 3950
rect 13105 3898 13120 3950
rect 13172 3898 13187 3950
rect 13239 3898 13254 3950
rect 13306 3898 13321 3950
rect 13373 3898 13388 3950
rect 13440 3898 13455 3950
rect 13507 3898 14039 3950
rect 441 2973 641 3074
rect 4511 2658 4997 2659
rect 4511 2606 4517 2658
rect 4569 2606 4602 2658
rect 4654 2606 4687 2658
rect 4739 2606 4771 2658
rect 4823 2606 4855 2658
rect 4907 2606 4939 2658
rect 4991 2606 4997 2658
tri 2390 2540 2396 2546 ne
rect 2396 2540 2402 2592
rect 2454 2540 2466 2592
rect 2518 2540 2524 2592
tri 2524 2540 2530 2546 nw
rect 4511 2542 4997 2606
tri 1845 2490 1851 2496 se
rect 1851 2444 1857 2496
rect 1909 2444 1921 2496
rect 1973 2444 1979 2496
tri 1979 2490 1985 2496 sw
tri 3519 2490 3525 2496 se
rect 3525 2444 3531 2496
rect 3583 2444 3595 2496
rect 3647 2444 3653 2496
tri 3653 2490 3659 2496 sw
rect 4511 2490 4517 2542
rect 4569 2490 4602 2542
rect 4654 2490 4687 2542
rect 4739 2490 4771 2542
rect 4823 2490 4855 2542
rect 4907 2490 4939 2542
rect 4991 2490 4997 2542
tri 9569 2540 9575 2546 ne
rect 9575 2540 9581 2592
rect 9633 2540 9645 2592
rect 9697 2540 9703 2592
tri 9703 2540 9709 2546 nw
tri 8092 2490 8098 2496 se
rect 4511 2426 4997 2490
rect 8098 2444 8104 2496
rect 8156 2444 8170 2496
rect 8222 2444 8228 2496
tri 8228 2490 8234 2496 sw
tri 9764 2490 9770 2496 se
rect 9770 2444 9776 2496
rect 9828 2444 9842 2496
rect 9894 2444 9900 2496
tri 9900 2490 9906 2496 sw
rect 4511 2374 4517 2426
rect 4569 2374 4602 2426
rect 4654 2374 4687 2426
rect 4739 2374 4771 2426
rect 4823 2374 4855 2426
rect 4907 2374 4939 2426
rect 4991 2374 4997 2426
rect 4511 2373 4997 2374
rect 2077 1882 2129 1888
tri 245 1812 291 1858 sw
tri 2043 1812 2077 1846 se
rect 2077 1818 2129 1830
rect 225 1766 2077 1812
tri 2129 1812 2163 1846 sw
rect 2129 1766 3531 1812
rect 225 1760 3531 1766
rect 3583 1760 3595 1812
rect 3647 1760 3653 1812
rect 320 1680 8106 1732
rect 8158 1680 8170 1732
rect 8222 1680 9776 1732
rect 9828 1680 9840 1732
rect 9892 1680 9898 1732
rect 10167 1680 10173 1732
rect 10225 1680 10237 1732
rect 10289 1680 14541 1732
rect 14593 1680 14605 1732
rect 14657 1680 14663 1732
rect 320 1652 326 1680
tri 326 1652 354 1680 nw
tri 320 1646 326 1652 nw
rect 2447 1600 2453 1652
rect 2505 1600 2517 1652
rect 2569 1600 14621 1652
rect 14673 1600 14685 1652
rect 14737 1600 14743 1652
rect 896 1491 904 1543
rect 956 1491 968 1543
rect 1020 1491 1266 1543
rect 1318 1491 1330 1543
rect 1382 1491 5653 1543
rect 5705 1491 5742 1543
rect 5794 1491 5831 1543
rect 5883 1491 5920 1543
rect 5972 1491 6809 1543
rect 6861 1491 6873 1543
rect 6925 1491 8511 1543
rect 8563 1491 8575 1543
rect 8627 1491 9991 1543
rect 10043 1491 10055 1543
rect 10107 1491 11334 1543
rect 11386 1491 11398 1543
rect 11450 1491 12768 1543
rect 12820 1491 12832 1543
rect 12884 1491 14701 1543
rect 14753 1491 14765 1543
rect 14817 1491 14823 1543
rect 300 1453 352 1459
tri 352 1411 358 1417 sw
rect 655 1411 663 1463
rect 715 1411 727 1463
rect 779 1411 1570 1463
rect 1622 1411 1634 1463
rect 1686 1411 3100 1463
rect 3152 1411 3164 1463
rect 3216 1411 3875 1463
rect 3927 1411 3939 1463
rect 3991 1411 4003 1463
rect 4055 1411 4067 1463
rect 4119 1411 4131 1463
rect 4183 1411 7239 1463
rect 7291 1411 7303 1463
rect 7355 1411 8941 1463
rect 8993 1411 9005 1463
rect 9057 1411 10421 1463
rect 10473 1411 10485 1463
rect 10537 1411 11764 1463
rect 11816 1411 11828 1463
rect 11880 1411 13198 1463
rect 13250 1411 13262 1463
rect 13314 1411 14781 1463
rect 14833 1411 14845 1463
rect 14897 1411 14903 1463
rect 352 1401 358 1411
rect 300 1389 358 1401
rect 352 1383 358 1389
tri 358 1383 386 1411 sw
rect 352 1337 421 1383
rect 300 1331 421 1337
rect 473 1331 485 1383
rect 537 1331 1853 1383
rect 1905 1331 1917 1383
rect 1969 1331 3383 1383
rect 3435 1331 3447 1383
rect 3499 1331 7669 1383
rect 7721 1331 7733 1383
rect 7785 1331 9371 1383
rect 9423 1331 9435 1383
rect 9487 1331 10851 1383
rect 10903 1331 10915 1383
rect 10967 1331 12194 1383
rect 12246 1331 12258 1383
rect 12310 1331 13628 1383
rect 13680 1331 13692 1383
rect 13744 1331 14861 1383
rect 14913 1331 14925 1383
rect 14977 1331 14983 1383
rect 487 1263 573 1286
rect 647 1263 692 1286
rect 773 1263 825 1286
<< via1 >>
rect 321 9460 373 9512
rect 321 9434 373 9448
rect 321 9400 341 9434
rect 341 9400 373 9434
rect 321 9396 373 9400
rect 791 3969 843 4021
rect 857 3969 909 4021
rect 791 3905 843 3957
rect 857 3905 909 3957
rect 2141 3976 2193 4028
rect 2207 3976 2259 4028
rect 2141 3898 2193 3950
rect 2207 3898 2259 3950
rect 2703 3969 2755 4021
rect 2769 3969 2821 4021
rect 2703 3905 2755 3957
rect 2769 3905 2821 3957
rect 3816 3969 3868 4021
rect 3895 3969 3947 4021
rect 3974 3969 4026 4021
rect 4053 3969 4105 4021
rect 4131 3969 4183 4021
rect 3816 3905 3868 3957
rect 3895 3905 3947 3957
rect 3974 3905 4026 3957
rect 4053 3905 4105 3957
rect 4131 3905 4183 3957
rect 6109 3976 6161 4028
rect 6174 3976 6226 4028
rect 6239 3976 6291 4028
rect 6304 3976 6356 4028
rect 6368 3976 6420 4028
rect 6432 3976 6484 4028
rect 6496 3976 6548 4028
rect 6560 3976 6612 4028
rect 6624 3976 6676 4028
rect 6688 3976 6740 4028
rect 6752 3976 6804 4028
rect 6109 3904 6161 3956
rect 6174 3904 6226 3956
rect 6239 3904 6291 3956
rect 6304 3904 6356 3956
rect 6368 3904 6420 3956
rect 6432 3904 6484 3956
rect 6496 3904 6548 3956
rect 6560 3904 6612 3956
rect 6624 3904 6676 3956
rect 6688 3904 6740 3956
rect 6752 3904 6804 3956
rect 7663 3976 7715 4028
rect 7729 3976 7781 4028
rect 7663 3898 7715 3950
rect 7729 3898 7781 3950
rect 8595 3976 8647 4028
rect 8660 3976 8712 4028
rect 8724 3976 8776 4028
rect 8788 3976 8840 4028
rect 8595 3902 8647 3954
rect 8660 3902 8712 3954
rect 8724 3902 8776 3954
rect 8788 3902 8840 3954
rect 10220 3934 10272 3986
rect 10286 3934 10338 3986
rect 10352 3934 10404 3986
rect 10418 3934 10470 3986
rect 10483 3934 10535 3986
rect 10548 3934 10600 3986
rect 10613 3934 10665 3986
rect 10678 3934 10730 3986
rect 11631 3935 11683 3987
rect 11696 3935 11748 3987
rect 11761 3935 11813 3987
rect 11826 3935 11878 3987
rect 11891 3935 11943 3987
rect 11956 3935 12008 3987
rect 12021 3935 12073 3987
rect 13053 3976 13105 4028
rect 13120 3976 13172 4028
rect 13187 3976 13239 4028
rect 13254 3976 13306 4028
rect 13321 3976 13373 4028
rect 13388 3976 13440 4028
rect 13455 3976 13507 4028
rect 13053 3898 13105 3950
rect 13120 3898 13172 3950
rect 13187 3898 13239 3950
rect 13254 3898 13306 3950
rect 13321 3898 13373 3950
rect 13388 3898 13440 3950
rect 13455 3898 13507 3950
rect 4517 2606 4569 2658
rect 4602 2606 4654 2658
rect 4687 2606 4739 2658
rect 4771 2606 4823 2658
rect 4855 2606 4907 2658
rect 4939 2606 4991 2658
rect 2402 2540 2454 2592
rect 2466 2540 2518 2592
rect 1857 2444 1909 2496
rect 1921 2444 1973 2496
rect 3531 2444 3583 2496
rect 3595 2444 3647 2496
rect 4517 2490 4569 2542
rect 4602 2490 4654 2542
rect 4687 2490 4739 2542
rect 4771 2490 4823 2542
rect 4855 2490 4907 2542
rect 4939 2490 4991 2542
rect 9581 2540 9633 2592
rect 9645 2540 9697 2592
rect 8104 2444 8156 2496
rect 8170 2444 8222 2496
rect 9776 2444 9828 2496
rect 9842 2444 9894 2496
rect 4517 2374 4569 2426
rect 4602 2374 4654 2426
rect 4687 2374 4739 2426
rect 4771 2374 4823 2426
rect 4855 2374 4907 2426
rect 4939 2374 4991 2426
rect 2077 1830 2129 1882
rect 2077 1766 2129 1818
rect 3531 1760 3583 1812
rect 3595 1760 3647 1812
rect 8106 1680 8158 1732
rect 8170 1680 8222 1732
rect 9776 1680 9828 1732
rect 9840 1680 9892 1732
rect 10173 1680 10225 1732
rect 10237 1680 10289 1732
rect 14541 1680 14593 1732
rect 14605 1680 14657 1732
rect 2453 1600 2505 1652
rect 2517 1600 2569 1652
rect 14621 1600 14673 1652
rect 14685 1600 14737 1652
rect 904 1491 956 1543
rect 968 1491 1020 1543
rect 1266 1491 1318 1543
rect 1330 1491 1382 1543
rect 5653 1491 5705 1543
rect 5742 1491 5794 1543
rect 5831 1491 5883 1543
rect 5920 1491 5972 1543
rect 6809 1491 6861 1543
rect 6873 1491 6925 1543
rect 8511 1491 8563 1543
rect 8575 1491 8627 1543
rect 9991 1491 10043 1543
rect 10055 1491 10107 1543
rect 11334 1491 11386 1543
rect 11398 1491 11450 1543
rect 12768 1491 12820 1543
rect 12832 1491 12884 1543
rect 14701 1491 14753 1543
rect 14765 1491 14817 1543
rect 300 1401 352 1453
rect 663 1411 715 1463
rect 727 1411 779 1463
rect 1570 1411 1622 1463
rect 1634 1411 1686 1463
rect 3100 1411 3152 1463
rect 3164 1411 3216 1463
rect 3875 1411 3927 1463
rect 3939 1411 3991 1463
rect 4003 1411 4055 1463
rect 4067 1411 4119 1463
rect 4131 1411 4183 1463
rect 7239 1411 7291 1463
rect 7303 1411 7355 1463
rect 8941 1411 8993 1463
rect 9005 1411 9057 1463
rect 10421 1411 10473 1463
rect 10485 1411 10537 1463
rect 11764 1411 11816 1463
rect 11828 1411 11880 1463
rect 13198 1411 13250 1463
rect 13262 1411 13314 1463
rect 14781 1411 14833 1463
rect 14845 1411 14897 1463
rect 300 1337 352 1389
rect 421 1331 473 1383
rect 485 1331 537 1383
rect 1853 1331 1905 1383
rect 1917 1331 1969 1383
rect 3383 1331 3435 1383
rect 3447 1331 3499 1383
rect 7669 1331 7721 1383
rect 7733 1331 7785 1383
rect 9371 1331 9423 1383
rect 9435 1331 9487 1383
rect 10851 1331 10903 1383
rect 10915 1331 10967 1383
rect 12194 1331 12246 1383
rect 12258 1331 12310 1383
rect 13628 1331 13680 1383
rect 13692 1331 13744 1383
rect 14861 1331 14913 1383
rect 14925 1331 14977 1383
<< metal2 >>
rect 12150 28507 12206 31368
tri 12206 28507 12226 28527 sw
rect 12150 28505 12226 28507
tri 12150 28429 12226 28505 ne
tri 12226 28429 12304 28507 sw
tri 12226 28351 12304 28429 ne
tri 12304 28351 12382 28429 sw
tri 12304 28273 12382 28351 ne
tri 12382 28273 12460 28351 sw
tri 12382 28239 12416 28273 ne
rect 12416 28239 12998 28273
tri 12998 28239 13032 28273 sw
tri 12416 28217 12438 28239 ne
rect 12438 28217 13032 28239
tri 12976 28161 13032 28217 ne
tri 13032 28161 13110 28239 sw
tri 13032 28083 13110 28161 ne
tri 13110 28083 13188 28161 sw
tri 13110 28061 13132 28083 ne
rect 13132 27555 13188 28083
tri 13188 27555 13193 27560 sw
rect 13132 27538 13193 27555
tri 13132 27490 13180 27538 ne
rect 13180 27499 13193 27538
tri 13193 27499 13249 27555 sw
tri 14274 27499 14330 27555 se
rect 14330 27499 14400 27555
rect 14456 27499 14480 27555
rect 14536 27499 14545 27555
rect 13180 27490 13249 27499
tri 13249 27490 13258 27499 sw
tri 14265 27490 14274 27499 se
rect 14274 27490 14330 27499
tri 13180 27482 13188 27490 ne
rect 13188 27482 13258 27490
tri 13188 27412 13258 27482 ne
tri 13258 27477 13271 27490 sw
tri 14252 27477 14265 27490 se
rect 14265 27477 14330 27490
tri 14330 27477 14352 27499 nw
rect 13258 27412 13271 27477
tri 13271 27412 13336 27477 sw
tri 14187 27412 14252 27477 se
tri 13258 27334 13336 27412 ne
tri 13336 27399 13349 27412 sw
tri 14174 27399 14187 27412 se
rect 14187 27399 14252 27412
tri 14252 27399 14330 27477 nw
rect 13336 27334 13349 27399
tri 13349 27334 13414 27399 sw
tri 14109 27334 14174 27399 se
rect 14174 27334 14187 27399
tri 14187 27334 14252 27399 nw
tri 13336 27278 13392 27334 ne
rect 13392 27278 14131 27334
tri 14131 27278 14187 27334 nw
rect 321 9512 373 9520
rect 321 9448 373 9460
rect 321 9375 373 9396
rect 321 1992 352 9375
tri 352 9354 373 9375 nw
rect 10509 5802 12816 6927
rect 5016 4408 6787 5353
rect 785 4021 915 4028
rect 785 3969 791 4021
rect 843 3969 857 4021
rect 909 3969 915 4021
tri 1750 3976 1802 4028 se
rect 1802 3976 2141 4028
rect 2193 3976 2207 4028
rect 2259 3976 2265 4028
tri 1743 3969 1750 3976 se
rect 1750 3969 2265 3976
rect 785 3957 915 3969
tri 1731 3957 1743 3969 se
rect 1743 3957 2265 3969
rect 785 3905 791 3957
rect 843 3905 857 3957
rect 909 3905 915 3957
tri 1724 3950 1731 3957 se
rect 1731 3950 2265 3957
tri 715 3387 785 3457 se
rect 785 3387 915 3905
tri 1676 3902 1724 3950 se
rect 1724 3902 2141 3950
tri 1672 3898 1676 3902 se
rect 1676 3898 2141 3902
rect 2193 3898 2207 3950
rect 2259 3898 2265 3950
rect 2697 4021 2827 4028
rect 2697 3969 2703 4021
rect 2755 3969 2769 4021
rect 2821 3969 2827 4021
rect 2697 3957 2827 3969
rect 2697 3905 2703 3957
rect 2755 3905 2769 3957
rect 2821 3905 2827 3957
tri 1618 3844 1672 3898 se
rect 1672 3844 1802 3898
tri 1802 3844 1856 3898 nw
rect 584 3257 915 3387
tri 1497 3723 1618 3844 se
rect 1618 3723 1681 3844
tri 1681 3723 1802 3844 nw
tri 524 2106 584 2166 se
rect 584 2106 714 3257
tri 714 3187 784 3257 nw
tri 1464 2160 1497 2193 se
rect 1497 2160 1627 3723
tri 1627 3669 1681 3723 nw
rect 2697 3319 2827 3905
rect 3810 4021 4189 4028
rect 3810 3969 3816 4021
rect 3868 3969 3895 4021
rect 3947 3969 3974 4021
rect 4026 3969 4053 4021
rect 4105 3969 4131 4021
rect 4183 3969 4189 4021
rect 3810 3957 4189 3969
rect 3810 3905 3816 3957
rect 3868 3905 3895 3957
rect 3947 3905 3974 3957
rect 4026 3905 4053 3957
rect 4105 3905 4131 3957
rect 4183 3905 4189 3957
tri 2827 3319 2852 3344 sw
rect 2697 3290 2852 3319
tri 2697 3135 2852 3290 ne
tri 2852 3135 3036 3319 sw
tri 2852 2951 3036 3135 ne
tri 3036 2951 3220 3135 sw
tri 3036 2897 3090 2951 ne
rect 2396 2540 2402 2592
rect 2454 2540 2466 2592
rect 2518 2540 2524 2592
tri 2396 2515 2421 2540 ne
rect 2421 2515 2499 2540
tri 2499 2515 2524 2540 nw
tri 2421 2496 2440 2515 ne
rect 2440 2496 2499 2515
rect 1851 2444 1857 2496
rect 1909 2444 1921 2496
rect 1973 2444 1979 2496
tri 2440 2489 2447 2496 ne
rect 1851 2401 1979 2444
tri 1851 2374 1878 2401 ne
rect 1878 2374 1979 2401
tri 1878 2347 1905 2374 ne
rect 1905 2347 1979 2374
tri 1905 2345 1907 2347 ne
rect 1907 2345 1979 2347
tri 1979 2345 1981 2347 sw
tri 1907 2273 1979 2345 ne
rect 1979 2273 1981 2345
tri 1979 2271 1981 2273 ne
tri 1981 2271 2055 2345 sw
tri 1981 2197 2055 2271 ne
tri 2055 2197 2129 2271 sw
tri 2055 2193 2059 2197 ne
rect 2059 2193 2129 2197
tri 714 2106 768 2160 sw
tri 1410 2106 1464 2160 se
rect 1464 2106 1627 2160
tri 1627 2106 1714 2193 sw
tri 2059 2175 2077 2193 ne
tri 352 1992 357 1997 sw
rect 413 1992 1026 2106
rect 321 1986 357 1992
tri 321 1965 342 1986 ne
rect 342 1965 357 1986
tri 357 1965 384 1992 sw
tri 342 1958 349 1965 ne
rect 349 1958 384 1965
tri 349 1956 351 1958 ne
rect 351 1956 384 1958
tri 351 1955 352 1956 ne
rect 352 1955 384 1956
tri 352 1953 354 1955 ne
tri 321 1551 354 1584 se
rect 354 1572 384 1955
rect 413 1940 543 1992
tri 543 1958 577 1992 nw
tri 621 1958 655 1992 ne
rect 414 1938 542 1939
rect 655 1940 785 1992
tri 785 1958 819 1992 nw
tri 862 1958 896 1992 ne
rect 656 1938 784 1939
rect 896 1940 1026 1992
rect 897 1938 1025 1939
rect 1260 1992 1977 2106
rect 1260 1958 1392 1992
tri 1392 1958 1426 1992 nw
tri 1528 1958 1562 1992 ne
rect 1562 1958 1696 1992
tri 1696 1958 1730 1992 nw
tri 1811 1958 1845 1992 ne
rect 1845 1958 1977 1992
rect 1260 1940 1390 1958
tri 1390 1956 1392 1958 nw
tri 1562 1956 1564 1958 ne
rect 1261 1938 1389 1939
rect 1564 1940 1694 1958
tri 1694 1956 1696 1958 nw
tri 1845 1956 1847 1958 ne
rect 1565 1938 1693 1939
rect 1847 1940 1977 1958
rect 1848 1938 1976 1939
rect 655 1638 785 1938
rect 1260 1638 1390 1938
rect 2077 1882 2129 2193
rect 2077 1818 2129 1830
rect 2077 1760 2129 1766
rect 2447 1680 2499 2496
tri 3003 2106 3090 2193 se
rect 3090 2106 3220 2951
rect 2790 1992 3220 2106
rect 3525 2444 3531 2496
rect 3583 2444 3595 2496
rect 3647 2444 3653 2496
rect 2790 1958 2922 1992
tri 2922 1958 2956 1992 nw
tri 2499 1680 2547 1728 sw
rect 2447 1652 2547 1680
tri 2547 1652 2575 1680 sw
rect 354 1551 363 1572
tri 363 1551 384 1572 nw
rect 414 1637 542 1638
rect 321 1543 355 1551
tri 355 1543 363 1551 nw
rect 321 1459 352 1543
tri 352 1540 355 1543 nw
rect 300 1453 352 1459
rect 300 1389 352 1401
rect 300 1331 352 1337
rect 413 1383 543 1636
rect 656 1637 784 1638
rect 655 1463 785 1636
rect 897 1637 1025 1638
rect 896 1543 1026 1636
rect 896 1491 904 1543
rect 956 1491 968 1543
rect 1020 1491 1026 1543
rect 1261 1637 1389 1638
rect 1260 1543 1390 1636
rect 1260 1491 1266 1543
rect 1318 1491 1330 1543
rect 1382 1491 1390 1543
rect 1565 1637 1693 1638
rect 655 1411 663 1463
rect 715 1411 727 1463
rect 779 1411 785 1463
rect 1564 1463 1694 1636
rect 1564 1411 1570 1463
rect 1622 1411 1634 1463
rect 1686 1411 1694 1463
rect 1848 1637 1976 1638
rect 413 1331 421 1383
rect 473 1331 485 1383
rect 537 1331 543 1383
rect 1847 1383 1977 1636
rect 2447 1600 2453 1652
rect 2505 1600 2517 1652
rect 2569 1600 2575 1652
rect 2790 1478 2920 1958
tri 2920 1956 2922 1958 nw
rect 3525 1812 3653 2444
rect 3525 1760 3531 1812
rect 3583 1760 3595 1812
rect 3647 1760 3653 1812
tri 2790 1463 2805 1478 ne
rect 2805 1463 2920 1478
tri 2805 1422 2846 1463 ne
rect 2846 1422 2920 1463
rect 3094 1463 3224 1584
tri 2846 1411 2857 1422 ne
rect 2857 1411 2920 1422
tri 2920 1411 2931 1422 sw
rect 3094 1411 3100 1463
rect 3152 1411 3164 1463
rect 3216 1411 3224 1463
tri 2857 1383 2885 1411 ne
rect 2885 1383 2931 1411
tri 2931 1383 2959 1411 sw
rect 3377 1383 3507 1584
rect 3810 1463 4189 3905
rect 5647 3976 6109 4028
rect 6161 3976 6174 4028
rect 6226 3976 6239 4028
rect 6291 3976 6304 4028
rect 6356 3976 6368 4028
rect 6420 3976 6432 4028
rect 6484 3976 6496 4028
rect 6548 3976 6560 4028
rect 6612 3976 6624 4028
rect 6676 3976 6688 4028
rect 6740 3976 6752 4028
rect 6804 3976 6810 4028
rect 5647 3956 6810 3976
rect 5647 3904 6109 3956
rect 6161 3904 6174 3956
rect 6226 3904 6239 3956
rect 6291 3904 6304 3956
rect 6356 3904 6368 3956
rect 6420 3904 6432 3956
rect 6484 3904 6496 3956
rect 6548 3904 6560 3956
rect 6612 3904 6624 3956
rect 6676 3904 6688 3956
rect 6740 3904 6752 3956
rect 6804 3904 6810 3956
rect 7657 3976 7663 4028
rect 7715 3976 7729 4028
rect 7781 3976 7787 4028
rect 7657 3950 7787 3976
rect 5647 3898 6107 3904
tri 6107 3898 6113 3904 nw
rect 7657 3898 7663 3950
rect 7715 3898 7729 3950
rect 7781 3898 7787 3950
rect 4511 2658 4520 2663
rect 4576 2658 4625 2663
rect 4681 2658 4730 2663
rect 4786 2658 4834 2663
rect 4890 2658 4938 2663
rect 4511 2606 4517 2658
rect 4576 2607 4602 2658
rect 4681 2607 4687 2658
rect 4823 2607 4834 2658
rect 4907 2607 4938 2658
rect 4994 2607 5003 2663
rect 4569 2606 4602 2607
rect 4654 2606 4687 2607
rect 4739 2606 4771 2607
rect 4823 2606 4855 2607
rect 4907 2606 4939 2607
rect 4991 2606 5003 2607
rect 4511 2543 5003 2606
rect 4511 2542 4520 2543
rect 4576 2542 4625 2543
rect 4681 2542 4730 2543
rect 4786 2542 4834 2543
rect 4890 2542 4938 2543
rect 4511 2490 4517 2542
rect 4576 2490 4602 2542
rect 4681 2490 4687 2542
rect 4823 2490 4834 2542
rect 4907 2490 4938 2542
rect 4511 2487 4520 2490
rect 4576 2487 4625 2490
rect 4681 2487 4730 2490
rect 4786 2487 4834 2490
rect 4890 2487 4938 2490
rect 4994 2487 5003 2543
rect 4511 2426 5003 2487
rect 4511 2374 4517 2426
rect 4569 2423 4602 2426
rect 4654 2423 4687 2426
rect 4739 2423 4771 2426
rect 4823 2423 4855 2426
rect 4907 2423 4939 2426
rect 4991 2423 5003 2426
rect 4576 2374 4602 2423
rect 4681 2374 4687 2423
rect 4823 2374 4834 2423
rect 4907 2374 4938 2423
rect 4511 2367 4520 2374
rect 4576 2367 4625 2374
rect 4681 2367 4730 2374
rect 4786 2367 4834 2374
rect 4890 2367 4938 2374
rect 4994 2367 5003 2423
rect 5647 1543 5978 3898
tri 5978 3769 6107 3898 nw
tri 7463 2224 7657 2418 se
rect 7657 2224 7787 3898
rect 8589 3976 8595 4028
rect 8647 3976 8660 4028
rect 8712 3976 8724 4028
rect 8776 3976 8788 4028
rect 8840 3976 8846 4028
rect 8589 3954 8846 3976
rect 8589 3902 8595 3954
rect 8647 3902 8660 3954
rect 8712 3902 8724 3954
rect 8776 3902 8788 3954
rect 8840 3902 8846 3954
rect 8098 2444 8104 2496
rect 8156 2444 8170 2496
rect 8222 2444 8228 2496
tri 7457 2218 7463 2224 se
rect 7463 2218 7787 2224
tri 7787 2218 7793 2224 sw
tri 7389 2150 7457 2218 se
rect 7457 2150 7793 2218
tri 7345 2106 7389 2150 se
rect 7389 2106 7793 2150
rect 6803 1992 7793 2106
rect 6803 1958 6935 1992
tri 6935 1958 6969 1992 nw
tri 7197 1958 7231 1992 ne
rect 7231 1958 7363 1992
rect 6803 1940 6933 1958
tri 6933 1956 6935 1958 nw
tri 7231 1956 7233 1958 ne
rect 6804 1938 6932 1939
rect 7233 1940 7363 1958
tri 7363 1956 7399 1992 nw
tri 7627 1956 7663 1992 ne
rect 7234 1938 7362 1939
rect 7663 1940 7793 1992
rect 7664 1938 7792 1939
rect 7233 1638 7363 1938
rect 8098 1732 8228 2444
tri 8545 2106 8589 2150 se
rect 8589 2106 8846 3902
rect 10214 3986 10736 4017
rect 10214 3934 10220 3986
rect 10272 3934 10286 3986
rect 10338 3934 10352 3986
rect 10404 3934 10418 3986
rect 10470 3934 10483 3986
rect 10535 3934 10548 3986
rect 10600 3934 10613 3986
rect 10665 3934 10678 3986
rect 10730 3934 10736 3986
rect 8958 2607 8967 2663
rect 9023 2607 9084 2663
rect 9140 2607 9201 2663
rect 9257 2607 9266 2663
rect 8958 2543 9266 2607
rect 8958 2487 8967 2543
rect 9023 2487 9084 2543
rect 9140 2487 9201 2543
rect 9257 2487 9266 2543
rect 9575 2540 9581 2592
rect 9633 2540 9645 2592
rect 9697 2540 9703 2592
tri 9575 2511 9604 2540 ne
rect 9604 2511 9674 2540
tri 9674 2511 9703 2540 nw
tri 9604 2496 9619 2511 ne
rect 9619 2496 9674 2511
tri 9619 2493 9622 2496 ne
rect 8958 2423 9266 2487
rect 8958 2367 8967 2423
rect 9023 2367 9084 2423
rect 9140 2367 9201 2423
rect 9257 2367 9266 2423
tri 8846 2106 8896 2156 sw
tri 8505 2066 8545 2106 se
rect 8545 2066 8896 2106
tri 8896 2066 8936 2106 sw
rect 8505 1992 9495 2066
rect 8505 1940 8635 1992
tri 8635 1956 8671 1992 nw
tri 8899 1956 8935 1992 ne
rect 8506 1938 8634 1939
rect 8935 1940 9065 1992
tri 9065 1956 9101 1992 nw
tri 9329 1956 9365 1992 ne
rect 8936 1938 9064 1939
rect 9365 1940 9495 1992
rect 9366 1938 9494 1939
rect 8098 1680 8106 1732
rect 8158 1680 8170 1732
rect 8222 1680 8228 1732
rect 8935 1638 9065 1938
rect 5647 1491 5653 1543
rect 5705 1491 5742 1543
rect 5794 1491 5831 1543
rect 5883 1491 5920 1543
rect 5972 1491 5978 1543
rect 6804 1637 6932 1638
rect 6803 1543 6933 1636
rect 6803 1491 6809 1543
rect 6861 1491 6873 1543
rect 6925 1491 6933 1543
rect 7234 1637 7362 1638
rect 3810 1411 3875 1463
rect 3927 1411 3939 1463
rect 3991 1411 4003 1463
rect 4055 1411 4067 1463
rect 4119 1411 4131 1463
rect 4183 1411 4189 1463
rect 7233 1463 7363 1636
rect 7233 1411 7239 1463
rect 7291 1411 7303 1463
rect 7355 1411 7363 1463
rect 7664 1637 7792 1638
rect 1847 1331 1853 1383
rect 1905 1331 1917 1383
rect 1969 1331 1977 1383
tri 2885 1354 2914 1383 ne
rect 2914 1354 2959 1383
tri 2959 1354 2988 1383 sw
tri 2914 1348 2920 1354 ne
rect 2920 1348 2988 1354
tri 2920 1331 2937 1348 ne
rect 2937 1331 2988 1348
tri 2988 1331 3011 1354 sw
rect 3377 1331 3383 1383
rect 3435 1331 3447 1383
rect 3499 1331 3507 1383
rect 7663 1383 7793 1636
rect 8506 1637 8634 1638
rect 8505 1543 8635 1636
rect 8505 1491 8511 1543
rect 8563 1491 8575 1543
rect 8627 1491 8635 1543
rect 8936 1637 9064 1638
rect 8935 1463 9065 1636
rect 8935 1411 8941 1463
rect 8993 1411 9005 1463
rect 9057 1411 9065 1463
rect 9366 1637 9494 1638
rect 7663 1331 7669 1383
rect 7721 1331 7733 1383
rect 7785 1331 7793 1383
rect 9365 1383 9495 1636
rect 9622 1463 9674 2496
rect 9770 2444 9776 2496
rect 9828 2444 9842 2496
rect 9894 2444 9900 2496
rect 9770 1732 9900 2444
tri 10082 2106 10214 2238 se
rect 10214 2106 10736 3934
rect 11625 3987 12079 4018
rect 11625 3935 11631 3987
rect 11683 3935 11696 3987
rect 11748 3935 11761 3987
rect 11813 3935 11826 3987
rect 11878 3935 11891 3987
rect 11943 3935 11956 3987
rect 12008 3935 12021 3987
rect 12073 3935 12079 3987
tri 11557 2238 11625 2306 se
rect 11625 2238 12079 3935
rect 13047 3976 13053 4028
rect 13105 3976 13120 4028
rect 13172 3976 13187 4028
rect 13239 3976 13254 4028
rect 13306 3976 13321 4028
rect 13373 3976 13388 4028
rect 13440 3976 13455 4028
rect 13507 3976 13513 4028
rect 13047 3950 13513 3976
rect 13047 3898 13053 3950
rect 13105 3898 13120 3950
rect 13172 3898 13187 3950
rect 13239 3898 13254 3950
rect 13306 3898 13321 3950
rect 13373 3898 13388 3950
rect 13440 3898 13455 3950
rect 13507 3898 13513 3950
tri 13017 2238 13047 2268 se
rect 13047 2238 13513 3898
tri 10736 2106 10868 2238 sw
tri 11425 2106 11557 2238 se
rect 11557 2106 12079 2238
tri 12079 2106 12211 2238 sw
tri 12991 2212 13017 2238 se
rect 13017 2212 13513 2238
tri 12885 2106 12991 2212 se
rect 12991 2106 13513 2212
tri 13513 2106 13619 2212 sw
rect 9985 1992 10975 2106
rect 9985 1940 10115 1992
tri 10115 1956 10151 1992 nw
tri 10379 1956 10415 1992 ne
rect 9986 1938 10114 1939
rect 10415 1940 10545 1992
tri 10545 1956 10581 1992 nw
tri 10809 1956 10845 1992 ne
rect 10416 1938 10544 1939
rect 10845 1940 10975 1992
rect 10846 1938 10974 1939
rect 11328 1992 12318 2106
rect 11328 1940 11458 1992
tri 11458 1956 11494 1992 nw
tri 11722 1956 11758 1992 ne
rect 11329 1938 11457 1939
rect 11758 1940 11888 1992
tri 11888 1956 11924 1992 nw
tri 12152 1956 12188 1992 ne
rect 11759 1938 11887 1939
rect 12188 1940 12318 1992
rect 12189 1938 12317 1939
rect 12762 1992 13752 2106
rect 12762 1940 12892 1992
tri 12892 1956 12928 1992 nw
tri 13156 1956 13192 1992 ne
rect 12763 1938 12891 1939
rect 13192 1940 13322 1992
tri 13322 1956 13358 1992 nw
tri 13586 1956 13622 1992 ne
rect 13193 1938 13321 1939
rect 13622 1940 13752 1992
rect 13623 1938 13751 1939
rect 9770 1680 9776 1732
rect 9828 1680 9840 1732
rect 9892 1680 9900 1732
rect 10167 1680 10173 1732
rect 10225 1680 10237 1732
rect 10289 1680 10295 1732
tri 10180 1652 10208 1680 ne
rect 10208 1652 10267 1680
tri 10267 1652 10295 1680 nw
tri 10208 1646 10214 1652 ne
rect 9986 1637 10114 1638
rect 9985 1543 10115 1636
rect 9985 1491 9991 1543
rect 10043 1491 10055 1543
rect 10107 1491 10115 1543
tri 9674 1463 9686 1475 sw
rect 9622 1453 9686 1463
tri 9622 1441 9634 1453 ne
rect 9634 1441 9686 1453
tri 9686 1441 9708 1463 sw
tri 9634 1411 9664 1441 ne
rect 9664 1426 9708 1441
tri 9708 1426 9723 1441 sw
rect 9664 1411 9723 1426
tri 9723 1411 9738 1426 sw
tri 10199 1411 10214 1426 se
rect 10214 1411 10266 1652
tri 10266 1651 10267 1652 nw
rect 10415 1638 10545 1938
rect 11758 1638 11888 1938
rect 13622 1638 13752 1938
tri 14589 1732 14623 1766 se
rect 14535 1680 14541 1732
rect 14593 1680 14605 1732
rect 14657 1680 14663 1732
tri 14675 1652 14703 1680 se
rect 10416 1637 10544 1638
rect 10415 1463 10545 1636
rect 10415 1411 10421 1463
rect 10473 1411 10485 1463
rect 10537 1411 10545 1463
rect 10846 1637 10974 1638
tri 9664 1401 9674 1411 ne
rect 9674 1401 9738 1411
tri 9674 1383 9692 1401 ne
rect 9692 1383 9738 1401
tri 9738 1383 9766 1411 sw
tri 10171 1383 10199 1411 se
rect 10199 1404 10266 1411
rect 10199 1383 10245 1404
tri 10245 1383 10266 1404 nw
rect 10845 1383 10975 1636
rect 11329 1637 11457 1638
rect 11328 1543 11458 1636
rect 11328 1491 11334 1543
rect 11386 1491 11398 1543
rect 11450 1491 11458 1543
rect 11759 1637 11887 1638
rect 11758 1463 11888 1636
rect 11758 1411 11764 1463
rect 11816 1411 11828 1463
rect 11880 1411 11888 1463
rect 12189 1637 12317 1638
rect 9365 1331 9371 1383
rect 9423 1331 9435 1383
rect 9487 1331 9495 1383
tri 9692 1367 9708 1383 ne
rect 9708 1367 9766 1383
tri 9766 1367 9782 1383 sw
tri 10155 1367 10171 1383 se
rect 10171 1367 10229 1383
tri 10229 1367 10245 1383 nw
tri 9708 1331 9744 1367 ne
rect 9744 1331 10193 1367
tri 10193 1331 10229 1367 nw
rect 10845 1331 10851 1383
rect 10903 1331 10915 1383
rect 10967 1331 10975 1383
rect 12188 1383 12318 1636
rect 12763 1637 12891 1638
rect 12762 1543 12892 1636
rect 12762 1491 12768 1543
rect 12820 1491 12832 1543
rect 12884 1491 12892 1543
rect 13193 1637 13321 1638
rect 13192 1463 13322 1636
rect 13192 1411 13198 1463
rect 13250 1411 13262 1463
rect 13314 1411 13322 1463
rect 13623 1637 13751 1638
rect 12188 1331 12194 1383
rect 12246 1331 12258 1383
rect 12310 1331 12318 1383
rect 13622 1383 13752 1636
rect 14615 1600 14621 1652
rect 14673 1600 14685 1652
rect 14737 1600 14743 1652
tri 14755 1543 14783 1571 se
rect 14695 1491 14701 1543
rect 14753 1491 14765 1543
rect 14817 1491 14823 1543
tri 14835 1463 14863 1491 se
rect 14775 1411 14781 1463
rect 14833 1411 14845 1463
rect 14897 1411 14903 1463
tri 14915 1383 14943 1411 se
rect 13622 1331 13628 1383
rect 13680 1331 13692 1383
rect 13744 1331 13752 1383
rect 14855 1331 14861 1383
rect 14913 1331 14925 1383
rect 14977 1331 14983 1383
tri 2937 1280 2988 1331 ne
rect 2988 1315 3011 1331
tri 3011 1315 3027 1331 sw
tri 9744 1315 9760 1331 ne
rect 9760 1315 10177 1331
tri 10177 1315 10193 1331 nw
rect 2988 1290 3027 1315
tri 3027 1290 3052 1315 sw
rect 2988 1280 3052 1290
tri 3052 1280 3062 1290 sw
rect 14506 1281 14562 1290
tri 2988 1206 3062 1280 ne
tri 3062 1242 3100 1280 sw
rect 3062 1206 3100 1242
tri 3100 1206 3136 1242 sw
tri 14470 1206 14506 1242 se
rect 14506 1206 14562 1225
tri 3062 1154 3114 1206 ne
rect 3114 1201 14562 1206
rect 3114 1154 14506 1201
tri 14488 1136 14506 1154 ne
rect 14506 1136 14562 1145
<< rmetal2 >>
rect 413 1939 543 1940
rect 413 1938 414 1939
rect 542 1938 543 1939
rect 655 1939 785 1940
rect 655 1938 656 1939
rect 784 1938 785 1939
rect 896 1939 1026 1940
rect 896 1938 897 1939
rect 1025 1938 1026 1939
rect 1260 1939 1390 1940
rect 1260 1938 1261 1939
rect 1389 1938 1390 1939
rect 1564 1939 1694 1940
rect 1564 1938 1565 1939
rect 1693 1938 1694 1939
rect 1847 1939 1977 1940
rect 1847 1938 1848 1939
rect 1976 1938 1977 1939
rect 413 1637 414 1638
rect 542 1637 543 1638
rect 413 1636 543 1637
rect 655 1637 656 1638
rect 784 1637 785 1638
rect 655 1636 785 1637
rect 896 1637 897 1638
rect 1025 1637 1026 1638
rect 896 1636 1026 1637
rect 1260 1637 1261 1638
rect 1389 1637 1390 1638
rect 1260 1636 1390 1637
rect 1564 1637 1565 1638
rect 1693 1637 1694 1638
rect 1564 1636 1694 1637
rect 1847 1637 1848 1638
rect 1976 1637 1977 1638
rect 1847 1636 1977 1637
rect 6803 1939 6933 1940
rect 6803 1938 6804 1939
rect 6932 1938 6933 1939
rect 7233 1939 7363 1940
rect 7233 1938 7234 1939
rect 7362 1938 7363 1939
rect 7663 1939 7793 1940
rect 7663 1938 7664 1939
rect 7792 1938 7793 1939
rect 8505 1939 8635 1940
rect 8505 1938 8506 1939
rect 8634 1938 8635 1939
rect 8935 1939 9065 1940
rect 8935 1938 8936 1939
rect 9064 1938 9065 1939
rect 9365 1939 9495 1940
rect 9365 1938 9366 1939
rect 9494 1938 9495 1939
rect 6803 1637 6804 1638
rect 6932 1637 6933 1638
rect 6803 1636 6933 1637
rect 7233 1637 7234 1638
rect 7362 1637 7363 1638
rect 7233 1636 7363 1637
rect 7663 1637 7664 1638
rect 7792 1637 7793 1638
rect 7663 1636 7793 1637
rect 8505 1637 8506 1638
rect 8634 1637 8635 1638
rect 8505 1636 8635 1637
rect 8935 1637 8936 1638
rect 9064 1637 9065 1638
rect 8935 1636 9065 1637
rect 9365 1637 9366 1638
rect 9494 1637 9495 1638
rect 9365 1636 9495 1637
rect 9985 1939 10115 1940
rect 9985 1938 9986 1939
rect 10114 1938 10115 1939
rect 10415 1939 10545 1940
rect 10415 1938 10416 1939
rect 10544 1938 10545 1939
rect 10845 1939 10975 1940
rect 10845 1938 10846 1939
rect 10974 1938 10975 1939
rect 11328 1939 11458 1940
rect 11328 1938 11329 1939
rect 11457 1938 11458 1939
rect 11758 1939 11888 1940
rect 11758 1938 11759 1939
rect 11887 1938 11888 1939
rect 12188 1939 12318 1940
rect 12188 1938 12189 1939
rect 12317 1938 12318 1939
rect 12762 1939 12892 1940
rect 12762 1938 12763 1939
rect 12891 1938 12892 1939
rect 13192 1939 13322 1940
rect 13192 1938 13193 1939
rect 13321 1938 13322 1939
rect 13622 1939 13752 1940
rect 13622 1938 13623 1939
rect 13751 1938 13752 1939
rect 9985 1637 9986 1638
rect 10114 1637 10115 1638
rect 9985 1636 10115 1637
rect 10415 1637 10416 1638
rect 10544 1637 10545 1638
rect 10415 1636 10545 1637
rect 10845 1637 10846 1638
rect 10974 1637 10975 1638
rect 10845 1636 10975 1637
rect 11328 1637 11329 1638
rect 11457 1637 11458 1638
rect 11328 1636 11458 1637
rect 11758 1637 11759 1638
rect 11887 1637 11888 1638
rect 11758 1636 11888 1637
rect 12188 1637 12189 1638
rect 12317 1637 12318 1638
rect 12188 1636 12318 1637
rect 12762 1637 12763 1638
rect 12891 1637 12892 1638
rect 12762 1636 12892 1637
rect 13192 1637 13193 1638
rect 13321 1637 13322 1638
rect 13192 1636 13322 1637
rect 13622 1637 13623 1638
rect 13751 1637 13752 1638
rect 13622 1636 13752 1637
<< via2 >>
rect 14400 27499 14456 27555
rect 14480 27499 14536 27555
rect 4520 2658 4576 2663
rect 4625 2658 4681 2663
rect 4730 2658 4786 2663
rect 4834 2658 4890 2663
rect 4938 2658 4994 2663
rect 4520 2607 4569 2658
rect 4569 2607 4576 2658
rect 4625 2607 4654 2658
rect 4654 2607 4681 2658
rect 4730 2607 4739 2658
rect 4739 2607 4771 2658
rect 4771 2607 4786 2658
rect 4834 2607 4855 2658
rect 4855 2607 4890 2658
rect 4938 2607 4939 2658
rect 4939 2607 4991 2658
rect 4991 2607 4994 2658
rect 4520 2542 4576 2543
rect 4625 2542 4681 2543
rect 4730 2542 4786 2543
rect 4834 2542 4890 2543
rect 4938 2542 4994 2543
rect 4520 2490 4569 2542
rect 4569 2490 4576 2542
rect 4625 2490 4654 2542
rect 4654 2490 4681 2542
rect 4730 2490 4739 2542
rect 4739 2490 4771 2542
rect 4771 2490 4786 2542
rect 4834 2490 4855 2542
rect 4855 2490 4890 2542
rect 4938 2490 4939 2542
rect 4939 2490 4991 2542
rect 4991 2490 4994 2542
rect 4520 2487 4576 2490
rect 4625 2487 4681 2490
rect 4730 2487 4786 2490
rect 4834 2487 4890 2490
rect 4938 2487 4994 2490
rect 4520 2374 4569 2423
rect 4569 2374 4576 2423
rect 4625 2374 4654 2423
rect 4654 2374 4681 2423
rect 4730 2374 4739 2423
rect 4739 2374 4771 2423
rect 4771 2374 4786 2423
rect 4834 2374 4855 2423
rect 4855 2374 4890 2423
rect 4938 2374 4939 2423
rect 4939 2374 4991 2423
rect 4991 2374 4994 2423
rect 4520 2367 4576 2374
rect 4625 2367 4681 2374
rect 4730 2367 4786 2374
rect 4834 2367 4890 2374
rect 4938 2367 4994 2374
rect 8967 2607 9023 2663
rect 9084 2607 9140 2663
rect 9201 2607 9257 2663
rect 8967 2487 9023 2543
rect 9084 2487 9140 2543
rect 9201 2487 9257 2543
rect 8967 2367 9023 2423
rect 9084 2367 9140 2423
rect 9201 2367 9257 2423
rect 14506 1225 14562 1281
rect 14506 1145 14562 1201
<< metal3 >>
rect 14395 27555 14567 27560
rect 14395 27499 14400 27555
rect 14456 27499 14480 27555
rect 14536 27499 14567 27555
rect 14395 27494 14567 27499
tri 14395 27388 14501 27494 ne
rect 4515 2663 4999 2668
rect 4515 2607 4520 2663
rect 4576 2607 4625 2663
rect 4681 2607 4730 2663
rect 4786 2607 4834 2663
rect 4890 2607 4938 2663
rect 4994 2607 4999 2663
rect 4515 2543 4999 2607
rect 4515 2487 4520 2543
rect 4576 2487 4625 2543
rect 4681 2487 4730 2543
rect 4786 2487 4834 2543
rect 4890 2487 4938 2543
rect 4994 2487 4999 2543
rect 4515 2423 4999 2487
rect 4515 2367 4520 2423
rect 4576 2367 4625 2423
rect 4681 2367 4730 2423
rect 4786 2367 4834 2423
rect 4890 2367 4938 2423
rect 4994 2367 4999 2423
rect 4515 2362 4999 2367
rect 8962 2663 9262 2668
rect 8962 2607 8967 2663
rect 9023 2607 9084 2663
rect 9140 2607 9201 2663
rect 9257 2607 9262 2663
rect 8962 2543 9262 2607
rect 8962 2487 8967 2543
rect 9023 2487 9084 2543
rect 9140 2487 9201 2543
rect 9257 2487 9262 2543
rect 8962 2423 9262 2487
rect 8962 2367 8967 2423
rect 9023 2367 9084 2423
rect 9140 2367 9201 2423
rect 9257 2367 9262 2423
rect 8962 2362 9262 2367
rect 14501 1281 14567 27494
rect 14501 1225 14506 1281
rect 14562 1225 14567 1281
rect 14501 1201 14567 1225
rect 14501 1145 14506 1201
rect 14562 1145 14567 1201
rect 14501 1140 14567 1145
use sky130_fd_pr__via_pol1_centered__example_559591418081  sky130_fd_pr__via_pol1_centered__example_559591418081_0
timestamp 1640697850
transform -1 0 2461 0 -1 9417
box 0 0 1 1
use sky130_fd_pr__via_pol1_centered__example_559591418081  sky130_fd_pr__via_pol1_centered__example_559591418081_1
timestamp 1640697850
transform 1 0 251 0 -1 9417
box 0 0 1 1
use sky130_fd_pr__res_generic_po__example_5595914180838  sky130_fd_pr__res_generic_po__example_5595914180838_0
timestamp 1640697850
transform 1 0 336 0 1 9367
box 15 17 2025 18
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_0
timestamp 1640697850
transform 0 -1 12892 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_1
timestamp 1640697850
transform 0 -1 11458 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_2
timestamp 1640697850
transform 0 -1 10115 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_3
timestamp 1640697850
transform 0 -1 8635 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_4
timestamp 1640697850
transform 0 -1 6933 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_5
timestamp 1640697850
transform 0 -1 13322 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_6
timestamp 1640697850
transform 0 -1 10975 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_7
timestamp 1640697850
transform 0 -1 9495 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_8
timestamp 1640697850
transform 0 -1 12318 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_9
timestamp 1640697850
transform 0 -1 7793 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_10
timestamp 1640697850
transform 0 -1 1977 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_11
timestamp 1640697850
transform 0 -1 1694 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_12
timestamp 1640697850
transform 0 1 413 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_13
timestamp 1640697850
transform 0 1 896 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_0
timestamp 1640697850
transform 0 -1 11888 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_1
timestamp 1640697850
transform 0 -1 7363 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_2
timestamp 1640697850
transform 0 -1 10545 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_3
timestamp 1640697850
transform 0 -1 9065 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_4
timestamp 1640697850
transform 0 -1 13752 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_5
timestamp 1640697850
transform 0 -1 1390 1 0 1584
box 0 24 408 28
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_6
timestamp 1640697850
transform 0 1 655 1 0 1584
box 0 24 408 28
use sky130_fd_io__nfet_con_diff_wo_abt_270v2  sky130_fd_io__nfet_con_diff_wo_abt_270v2_0
timestamp 1640697850
transform -1 0 15088 0 -1 8404
box 0 423 15173 5493
<< labels >>
flabel metal1 s 441 2973 641 3074 0 FreeSans 400 0 0 0 VCC_IO
port 1 nsew
flabel metal1 s 14692 1491 14777 1543 0 FreeSans 400 0 0 0 PD_H[2]
port 2 nsew
flabel metal1 s 14701 1411 14857 1463 0 FreeSans 400 0 0 0 PD_H[3]
port 3 nsew
flabel metal1 s 14833 1331 14937 1383 0 FreeSans 400 0 0 0 TIE_LO_ESD
port 4 nsew
flabel metal1 s 201 9395 292 9439 0 FreeSans 400 0 0 0 TIE_LO_ESD
port 4 nsew
flabel metal1 s 2427 9424 2499 9476 0 FreeSans 400 180 0 0 VGND_IO
port 5 nsew
flabel metal1 s 779 1270 819 1282 3 FreeSans 520 90 0 0 VSSIO_AMX
port 6 nsew
flabel metal1 s 653 1265 687 1275 3 FreeSans 520 90 0 0 FORCE_LOVOL_H
port 7 nsew
flabel metal1 s 490 1271 570 1286 3 FreeSans 520 90 0 0 FORCE_LO_H
port 8 nsew
flabel metal2 s 10509 5802 12816 6927 0 FreeSans 400 0 0 0 PAD
port 9 nsew
flabel metal2 s 5016 4408 6787 5353 0 FreeSans 400 0 0 0 VGND_IO
port 5 nsew
flabel metal2 s 2816 1991 2896 2063 3 FreeSans 520 0 0 0 PD_H_I2C
port 10 nsew
flabel comment s 1276 7506 1276 7506 0 FreeSans 440 180 0 0 CONDIODE
flabel comment s 1461 9429 1461 9429 0 FreeSans 440 0 0 0 LEAKER
flabel comment s 2310 1270 2310 1270 0 FreeSans 440 0 0 0 RES
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 4473848
string GDS_START 4438700
<< end >>
