magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1368 -1260 1405 1935
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_0
timestamp 1619729480
transform -1 0 -80 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808679  sky130_fd_pr__dfl1sd2__example_55959141808679_1
timestamp 1619729480
transform 1 0 117 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 145 675 145 675 0 FreeSans 300 0 0 0 D
flabel comment s -108 675 -108 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 9194500
string GDS_START 9193510
<< end >>
