magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1158 -3367 18499 39974
<< metal1 >>
rect 15049 7623 17239 7665
rect 15049 6931 15095 7623
rect 17195 6931 17239 7623
rect 15049 6891 17239 6931
rect 5107 -7 5683 57
rect 4099 -163 11313 -7
rect 15240 -163 17187 6891
rect 4099 -203 17187 -163
tri 3331 -603 3731 -203 se
rect 3731 -603 17187 -203
rect 3331 -1307 17187 -603
rect 3331 -1707 16387 -1307
tri 3331 -2107 3731 -1707 ne
rect 3731 -2107 16387 -1707
tri 16387 -2107 17187 -1307 nw
<< via1 >>
rect 15095 6931 17195 7623
<< metal2 >>
rect 132 38641 2749 38676
rect 132 34825 172 38641
rect 2708 34825 2749 38641
rect 132 34791 2749 34825
rect 14940 8802 17228 8840
rect 14940 7946 15165 8802
rect 16181 7946 17228 8802
rect 14940 7910 17228 7946
rect 15049 7623 17239 7665
rect 15049 6931 15095 7623
rect 17195 6931 17239 7623
rect 15049 6891 17239 6931
<< via2 >>
rect 172 34825 2708 38641
rect 15165 7946 16181 8802
rect 15136 6977 17192 7593
<< metal3 >>
rect 102 38645 2772 38714
rect 102 34821 168 38645
rect 2712 34821 2772 38645
rect 102 34753 2772 34821
rect 15121 8806 17228 8840
rect 15121 8802 15181 8806
rect 15121 7946 15165 8802
rect 15121 7942 15181 7946
rect 17165 7942 17228 8806
rect 15121 7910 17228 7942
rect 15088 7597 17228 7632
rect 15088 6973 15132 7597
rect 17196 6973 17228 7597
rect 15088 6939 17228 6973
rect 5228 2223 7341 2269
rect 5228 1439 5252 2223
rect 7316 1439 7341 2223
rect 5228 1394 7341 1439
rect 7705 2221 9818 2267
rect 7705 1437 7729 2221
rect 9793 1437 9818 2221
rect 7705 1392 9818 1437
<< via3 >>
rect 168 38641 2712 38645
rect 168 34825 172 38641
rect 172 34825 2708 38641
rect 2708 34825 2712 38641
rect 168 34821 2712 34825
rect 15181 8802 17165 8806
rect 15181 7946 16181 8802
rect 16181 7946 17165 8802
rect 15181 7942 17165 7946
rect 15132 7593 17196 7597
rect 15132 6977 15136 7593
rect 15136 6977 17192 7593
rect 17192 6977 17196 7593
rect 15132 6973 17196 6977
rect 5252 1439 7316 2223
rect 7729 1437 9793 2221
<< metal4 >>
rect 132 38645 2749 38676
rect 132 34821 168 38645
rect 2712 34821 2749 38645
rect 132 34791 2749 34821
rect 14940 8806 17228 8840
rect 14940 7942 15181 8806
rect 17165 7942 17228 8806
rect 14940 7910 17228 7942
rect 14985 7597 17233 7630
rect 14985 6973 15132 7597
rect 17196 6973 17233 7597
rect 14985 6940 17233 6973
rect 5228 2223 7341 2269
rect 5228 1439 5252 2223
rect 7316 1439 7341 2223
rect 5228 1394 7341 1439
rect 7705 2221 9818 2267
rect 7705 1437 7729 2221
rect 9793 1437 9818 2221
rect 7705 1392 9818 1437
<< properties >>
string FIXED_BBOX 0 -7 15000 39593
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_END 1552440
string GDS_START 1244300
<< end >>
