magic
tech sky130A
magscale 1 2
timestamp 1640697850
use sky130_fd_pr__hvdfm1sd2__example_55959141808210  sky130_fd_pr__hvdfm1sd2__example_55959141808210_0
timestamp 1640697850
transform 1 0 456 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808210  sky130_fd_pr__hvdfm1sd2__example_55959141808210_1
timestamp 1640697850
transform 1 0 968 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfm1sd2__example_55959141808219  sky130_fd_pr__dfm1sd2__example_55959141808219_0
timestamp 1640697850
transform 1 0 200 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfm1sd2__example_55959141808219  sky130_fd_pr__dfm1sd2__example_55959141808219_1
timestamp 1640697850
transform 1 0 712 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808207  sky130_fd_pr__hvdfm1sd__example_55959141808207_0
timestamp 1640697850
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808207  sky130_fd_pr__hvdfm1sd__example_55959141808207_1
timestamp 1640697850
transform 1 0 1224 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 1252 49 1252 49 0 FreeSans 300 0 0 0 D
flabel comment s 996 49 996 49 0 FreeSans 300 0 0 0 S
flabel comment s 740 49 740 49 0 FreeSans 300 0 0 0 D
flabel comment s 484 49 484 49 0 FreeSans 300 0 0 0 S
flabel comment s 228 49 228 49 0 FreeSans 300 0 0 0 D
flabel comment s -28 49 -28 49 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 37263422
string GDS_START 37260428
<< end >>
