magic
tech sky130A
timestamp 1619729480
<< checkpaint >>
rect -630 -630 780 2130
<< pdiff >>
rect 0 0 150 1500
use sky130_fd_io__gnd2gnd_strap  sky130_fd_io__gnd2gnd_strap_0
timestamp 1619729480
transform 1 0 0 0 1 0
box 0 0 150 1500
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 9282938
string GDS_START 9282754
<< end >>
