magic
tech sky130A
magscale 1 2
timestamp 1619729575
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 113 326 161 487
rect 281 326 329 487
rect 449 326 499 487
rect 616 326 665 487
rect 784 326 835 487
rect 953 326 1001 487
rect 23 292 1088 326
rect 23 173 57 292
rect 91 207 973 258
rect 1034 173 1088 292
rect 23 139 1088 173
rect 307 56 345 139
rect 479 56 517 139
rect 651 56 689 139
rect 823 56 861 139
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 27 360 79 527
rect 195 360 247 527
rect 363 360 415 527
rect 533 360 582 527
rect 699 360 750 527
rect 869 360 919 527
rect 1035 360 1086 527
rect 207 17 273 105
rect 379 17 445 105
rect 551 17 617 105
rect 723 17 789 105
rect 895 17 961 105
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 91 207 973 258 6 A
port 1 nsew signal input
rlabel locali s 1034 173 1088 292 6 Y
port 6 nsew signal output
rlabel locali s 953 326 1001 487 6 Y
port 6 nsew signal output
rlabel locali s 823 56 861 139 6 Y
port 6 nsew signal output
rlabel locali s 784 326 835 487 6 Y
port 6 nsew signal output
rlabel locali s 651 56 689 139 6 Y
port 6 nsew signal output
rlabel locali s 616 326 665 487 6 Y
port 6 nsew signal output
rlabel locali s 479 56 517 139 6 Y
port 6 nsew signal output
rlabel locali s 449 326 499 487 6 Y
port 6 nsew signal output
rlabel locali s 307 56 345 139 6 Y
port 6 nsew signal output
rlabel locali s 281 326 329 487 6 Y
port 6 nsew signal output
rlabel locali s 113 326 161 487 6 Y
port 6 nsew signal output
rlabel locali s 23 292 1088 326 6 Y
port 6 nsew signal output
rlabel locali s 23 173 57 292 6 Y
port 6 nsew signal output
rlabel locali s 23 139 1088 173 6 Y
port 6 nsew signal output
rlabel metal1 s 0 -48 1196 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 1234 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3682906
string GDS_START 3673716
<< end >>
