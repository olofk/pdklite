magic
tech sky130A
magscale 1 2
timestamp 1619729571
<< checkpaint >>
rect -1298 -1308 2862 1852
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1107 47 1137 177
rect 1203 47 1233 177
rect 1287 47 1317 177
rect 1371 47 1401 177
rect 1455 47 1485 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 855 297 885 497
rect 939 297 969 497
rect 1023 297 1053 497
rect 1107 297 1137 497
rect 1203 297 1233 497
rect 1287 297 1317 497
rect 1371 297 1401 497
rect 1455 297 1485 497
<< ndiff >>
rect 27 142 79 177
rect 27 108 35 142
rect 69 108 79 142
rect 27 47 79 108
rect 109 97 163 177
rect 109 63 119 97
rect 153 63 163 97
rect 109 47 163 63
rect 193 142 247 177
rect 193 108 203 142
rect 237 108 247 142
rect 193 47 247 108
rect 277 97 331 177
rect 277 63 287 97
rect 321 63 331 97
rect 277 47 331 63
rect 361 142 415 177
rect 361 108 371 142
rect 405 108 415 142
rect 361 47 415 108
rect 445 165 499 177
rect 445 131 455 165
rect 489 131 499 165
rect 445 47 499 131
rect 529 97 583 177
rect 529 63 539 97
rect 573 63 583 97
rect 529 47 583 63
rect 613 165 667 177
rect 613 131 623 165
rect 657 131 667 165
rect 613 47 667 131
rect 697 97 749 177
rect 697 63 707 97
rect 741 63 749 97
rect 697 47 749 63
rect 803 97 855 177
rect 803 63 811 97
rect 845 63 855 97
rect 803 47 855 63
rect 885 165 939 177
rect 885 131 895 165
rect 929 131 939 165
rect 885 47 939 131
rect 969 97 1023 177
rect 969 63 979 97
rect 1013 63 1023 97
rect 969 47 1023 63
rect 1053 165 1107 177
rect 1053 131 1063 165
rect 1097 131 1107 165
rect 1053 47 1107 131
rect 1137 165 1203 177
rect 1137 131 1154 165
rect 1188 131 1203 165
rect 1137 97 1203 131
rect 1137 63 1154 97
rect 1188 63 1203 97
rect 1137 47 1203 63
rect 1233 165 1287 177
rect 1233 131 1243 165
rect 1277 131 1287 165
rect 1233 47 1287 131
rect 1317 97 1371 177
rect 1317 63 1327 97
rect 1361 63 1371 97
rect 1317 47 1371 63
rect 1401 165 1455 177
rect 1401 131 1411 165
rect 1445 131 1455 165
rect 1401 47 1455 131
rect 1485 165 1537 177
rect 1485 131 1495 165
rect 1529 131 1537 165
rect 1485 97 1537 131
rect 1485 63 1495 97
rect 1529 63 1537 97
rect 1485 47 1537 63
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 417 331 451
rect 277 383 287 417
rect 321 383 331 417
rect 277 349 331 383
rect 277 315 287 349
rect 321 315 331 349
rect 277 297 331 315
rect 361 485 415 497
rect 361 451 371 485
rect 405 451 415 485
rect 361 417 415 451
rect 361 383 371 417
rect 405 383 415 417
rect 361 297 415 383
rect 445 485 499 497
rect 445 451 455 485
rect 489 451 499 485
rect 445 417 499 451
rect 445 383 455 417
rect 489 383 499 417
rect 445 349 499 383
rect 445 315 455 349
rect 489 315 499 349
rect 445 297 499 315
rect 529 485 583 497
rect 529 451 539 485
rect 573 451 583 485
rect 529 417 583 451
rect 529 383 539 417
rect 573 383 583 417
rect 529 297 583 383
rect 613 485 667 497
rect 613 451 623 485
rect 657 451 667 485
rect 613 417 667 451
rect 613 383 623 417
rect 657 383 667 417
rect 613 349 667 383
rect 613 315 623 349
rect 657 315 667 349
rect 613 297 667 315
rect 697 485 855 497
rect 697 451 707 485
rect 741 451 811 485
rect 845 451 855 485
rect 697 417 855 451
rect 697 383 707 417
rect 741 383 811 417
rect 845 383 855 417
rect 697 297 855 383
rect 885 485 939 497
rect 885 451 895 485
rect 929 451 939 485
rect 885 417 939 451
rect 885 383 895 417
rect 929 383 939 417
rect 885 349 939 383
rect 885 315 895 349
rect 929 315 939 349
rect 885 297 939 315
rect 969 485 1023 497
rect 969 451 979 485
rect 1013 451 1023 485
rect 969 417 1023 451
rect 969 383 979 417
rect 1013 383 1023 417
rect 969 297 1023 383
rect 1053 485 1107 497
rect 1053 451 1063 485
rect 1097 451 1107 485
rect 1053 417 1107 451
rect 1053 383 1063 417
rect 1097 383 1107 417
rect 1053 349 1107 383
rect 1053 315 1063 349
rect 1097 315 1107 349
rect 1053 297 1107 315
rect 1137 485 1203 497
rect 1137 451 1154 485
rect 1188 451 1203 485
rect 1137 417 1203 451
rect 1137 383 1154 417
rect 1188 383 1203 417
rect 1137 297 1203 383
rect 1233 485 1287 497
rect 1233 451 1243 485
rect 1277 451 1287 485
rect 1233 417 1287 451
rect 1233 383 1243 417
rect 1277 383 1287 417
rect 1233 349 1287 383
rect 1233 315 1243 349
rect 1277 315 1287 349
rect 1233 297 1287 315
rect 1317 485 1371 497
rect 1317 451 1327 485
rect 1361 451 1371 485
rect 1317 417 1371 451
rect 1317 383 1327 417
rect 1361 383 1371 417
rect 1317 297 1371 383
rect 1401 485 1455 497
rect 1401 451 1411 485
rect 1445 451 1455 485
rect 1401 417 1455 451
rect 1401 383 1411 417
rect 1445 383 1455 417
rect 1401 349 1455 383
rect 1401 315 1411 349
rect 1445 315 1455 349
rect 1401 297 1455 315
rect 1485 485 1537 497
rect 1485 451 1495 485
rect 1529 451 1537 485
rect 1485 417 1537 451
rect 1485 383 1495 417
rect 1529 383 1537 417
rect 1485 349 1537 383
rect 1485 315 1495 349
rect 1529 315 1537 349
rect 1485 297 1537 315
<< ndiffc >>
rect 35 108 69 142
rect 119 63 153 97
rect 203 108 237 142
rect 287 63 321 97
rect 371 108 405 142
rect 455 131 489 165
rect 539 63 573 97
rect 623 131 657 165
rect 707 63 741 97
rect 811 63 845 97
rect 895 131 929 165
rect 979 63 1013 97
rect 1063 131 1097 165
rect 1154 131 1188 165
rect 1154 63 1188 97
rect 1243 131 1277 165
rect 1327 63 1361 97
rect 1411 131 1445 165
rect 1495 131 1529 165
rect 1495 63 1529 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 203 383 237 417
rect 287 451 321 485
rect 287 383 321 417
rect 287 315 321 349
rect 371 451 405 485
rect 371 383 405 417
rect 455 451 489 485
rect 455 383 489 417
rect 455 315 489 349
rect 539 451 573 485
rect 539 383 573 417
rect 623 451 657 485
rect 623 383 657 417
rect 623 315 657 349
rect 707 451 741 485
rect 811 451 845 485
rect 707 383 741 417
rect 811 383 845 417
rect 895 451 929 485
rect 895 383 929 417
rect 895 315 929 349
rect 979 451 1013 485
rect 979 383 1013 417
rect 1063 451 1097 485
rect 1063 383 1097 417
rect 1063 315 1097 349
rect 1154 451 1188 485
rect 1154 383 1188 417
rect 1243 451 1277 485
rect 1243 383 1277 417
rect 1243 315 1277 349
rect 1327 451 1361 485
rect 1327 383 1361 417
rect 1411 451 1445 485
rect 1411 383 1445 417
rect 1411 315 1445 349
rect 1495 451 1529 485
rect 1495 383 1529 417
rect 1495 315 1529 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 855 497 885 523
rect 939 497 969 523
rect 1023 497 1053 523
rect 1107 497 1137 523
rect 1203 497 1233 523
rect 1287 497 1317 523
rect 1371 497 1401 523
rect 1455 497 1485 523
rect 79 261 109 297
rect 21 259 109 261
rect 163 259 193 297
rect 247 259 277 297
rect 331 259 361 297
rect 21 249 361 259
rect 21 215 38 249
rect 72 215 119 249
rect 153 215 203 249
rect 237 215 287 249
rect 321 215 361 249
rect 21 205 361 215
rect 21 203 109 205
rect 79 177 109 203
rect 163 177 193 205
rect 247 177 277 205
rect 331 177 361 205
rect 415 259 445 297
rect 499 259 529 297
rect 583 259 613 297
rect 667 259 697 297
rect 855 259 885 297
rect 939 259 969 297
rect 1023 259 1053 297
rect 1107 259 1137 297
rect 415 249 697 259
rect 415 215 454 249
rect 488 215 539 249
rect 573 215 623 249
rect 657 215 697 249
rect 415 205 697 215
rect 789 249 1137 259
rect 789 215 805 249
rect 839 215 895 249
rect 929 215 979 249
rect 1013 215 1063 249
rect 1097 215 1137 249
rect 789 205 1137 215
rect 415 177 445 205
rect 499 177 529 205
rect 583 177 613 205
rect 667 177 697 205
rect 855 177 885 205
rect 939 177 969 205
rect 1023 177 1053 205
rect 1107 177 1137 205
rect 1203 259 1233 297
rect 1287 259 1317 297
rect 1371 259 1401 297
rect 1455 261 1485 297
rect 1455 259 1542 261
rect 1203 249 1542 259
rect 1203 215 1309 249
rect 1343 215 1393 249
rect 1427 215 1492 249
rect 1526 215 1542 249
rect 1203 205 1542 215
rect 1203 177 1233 205
rect 1287 177 1317 205
rect 1371 177 1401 205
rect 1455 203 1542 205
rect 1455 177 1485 203
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1107 21 1137 47
rect 1203 21 1233 47
rect 1287 21 1317 47
rect 1371 21 1401 47
rect 1455 21 1485 47
<< polycont >>
rect 38 215 72 249
rect 119 215 153 249
rect 203 215 237 249
rect 287 215 321 249
rect 454 215 488 249
rect 539 215 573 249
rect 623 215 657 249
rect 805 215 839 249
rect 895 215 929 249
rect 979 215 1013 249
rect 1063 215 1097 249
rect 1309 215 1343 249
rect 1393 215 1427 249
rect 1492 215 1526 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 289 69 315
rect 103 485 169 493
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 203 485 237 527
rect 203 417 237 451
rect 203 367 237 383
rect 271 485 337 493
rect 271 451 287 485
rect 321 451 337 485
rect 271 417 337 451
rect 271 383 287 417
rect 321 383 337 417
rect 103 315 119 349
rect 153 333 169 349
rect 271 349 337 383
rect 371 485 405 527
rect 371 417 405 451
rect 371 367 405 383
rect 439 485 505 493
rect 439 451 455 485
rect 489 451 505 485
rect 439 417 505 451
rect 439 383 455 417
rect 489 383 505 417
rect 271 333 287 349
rect 153 315 287 333
rect 321 333 337 349
rect 439 349 505 383
rect 539 485 573 527
rect 539 417 573 451
rect 539 367 573 383
rect 607 485 673 493
rect 607 451 623 485
rect 657 451 673 485
rect 607 417 673 451
rect 607 383 623 417
rect 657 383 673 417
rect 439 333 455 349
rect 321 315 455 333
rect 489 333 505 349
rect 607 349 673 383
rect 707 485 845 527
rect 741 451 811 485
rect 707 417 845 451
rect 741 383 811 417
rect 707 367 845 383
rect 879 485 945 493
rect 879 451 895 485
rect 929 451 945 485
rect 879 417 945 451
rect 879 383 895 417
rect 929 383 945 417
rect 607 333 623 349
rect 489 315 623 333
rect 657 333 673 349
rect 879 349 945 383
rect 979 485 1013 527
rect 979 417 1013 451
rect 979 367 1013 383
rect 1047 485 1113 493
rect 1047 451 1063 485
rect 1097 451 1113 485
rect 1047 417 1113 451
rect 1047 383 1063 417
rect 1097 383 1113 417
rect 879 333 895 349
rect 657 315 895 333
rect 929 333 945 349
rect 1047 349 1113 383
rect 1154 485 1188 527
rect 1154 417 1188 451
rect 1154 367 1188 383
rect 1227 485 1293 493
rect 1227 451 1243 485
rect 1277 451 1293 485
rect 1227 417 1293 451
rect 1227 383 1243 417
rect 1277 383 1293 417
rect 1047 333 1063 349
rect 929 315 1063 333
rect 1097 333 1113 349
rect 1227 349 1293 383
rect 1327 485 1361 527
rect 1327 417 1361 451
rect 1327 367 1361 383
rect 1395 485 1461 493
rect 1395 451 1411 485
rect 1445 451 1461 485
rect 1395 417 1461 451
rect 1395 383 1411 417
rect 1445 383 1461 417
rect 1227 333 1243 349
rect 1097 315 1243 333
rect 1277 333 1293 349
rect 1395 349 1461 383
rect 1395 333 1411 349
rect 1277 315 1411 333
rect 1445 315 1461 349
rect 103 289 1461 315
rect 1495 485 1547 527
rect 1529 451 1547 485
rect 1495 417 1547 451
rect 1529 383 1547 417
rect 1495 349 1547 383
rect 1529 315 1547 349
rect 1495 289 1547 315
rect 21 249 340 255
rect 21 215 38 249
rect 72 215 119 249
rect 153 215 203 249
rect 237 215 287 249
rect 321 215 340 249
rect 398 249 708 255
rect 398 215 454 249
rect 488 215 539 249
rect 573 215 623 249
rect 657 215 708 249
rect 770 249 1113 255
rect 770 215 805 249
rect 839 215 895 249
rect 929 215 979 249
rect 1013 215 1063 249
rect 1097 215 1113 249
rect 1222 181 1258 289
rect 1293 249 1542 255
rect 1293 215 1309 249
rect 1343 215 1393 249
rect 1427 215 1492 249
rect 1526 215 1542 249
rect 18 142 405 181
rect 18 108 35 142
rect 69 131 203 142
rect 18 51 69 108
rect 237 131 371 142
rect 103 63 119 97
rect 153 63 169 97
rect 103 17 169 63
rect 203 51 237 108
rect 439 165 1113 181
rect 439 131 455 165
rect 489 131 623 165
rect 657 131 895 165
rect 929 131 1063 165
rect 1097 131 1113 165
rect 1154 165 1188 181
rect 1222 165 1461 181
rect 1222 131 1243 165
rect 1277 131 1411 165
rect 1445 131 1461 165
rect 1495 165 1546 181
rect 1529 131 1546 165
rect 371 97 405 108
rect 1154 97 1188 131
rect 1495 97 1546 131
rect 271 63 287 97
rect 321 63 337 97
rect 271 17 337 63
rect 371 63 539 97
rect 573 63 707 97
rect 741 63 757 97
rect 371 51 757 63
rect 795 63 811 97
rect 845 63 979 97
rect 1013 63 1154 97
rect 1188 63 1327 97
rect 1361 63 1495 97
rect 1529 63 1546 97
rect 795 51 1546 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel locali s 1500 221 1534 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1408 221 1442 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1316 221 1350 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 674 221 708 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 770 221 804 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 862 221 896 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 954 221 988 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 1046 221 1080 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 1224 221 1258 255 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 nand4_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 111390
string GDS_START 97984
string path 0.000 2.720 7.820 2.720 
<< end >>
