magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1320 -1260 1388 1391
use sky130_fd_pr__dfl1sd2__example_55959141808104  sky130_fd_pr__dfl1sd2__example_55959141808104_0
timestamp 1619729480
transform -1 0 -32 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808104  sky130_fd_pr__dfl1sd2__example_55959141808104_1
timestamp 1619729480
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 131 128 131 0 FreeSans 300 0 0 0 D
flabel comment s -60 131 -60 131 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 40051448
string GDS_START 40050330
<< end >>
