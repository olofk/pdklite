magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1260 -1260 1619 2326
<< nwell >>
rect 0 394 359 1066
<< pwell >>
rect 258 32 292 232
<< nmos >>
rect 79 32 129 232
<< pmoshvt >>
rect 89 430 139 1030
<< ndiff >>
rect 26 214 79 232
rect 26 180 34 214
rect 68 180 79 214
rect 26 146 79 180
rect 26 112 34 146
rect 68 112 79 146
rect 26 78 79 112
rect 26 44 34 78
rect 68 44 79 78
rect 26 32 79 44
rect 129 214 182 232
rect 129 180 140 214
rect 174 180 182 214
rect 129 146 182 180
rect 129 112 140 146
rect 174 112 182 146
rect 129 78 182 112
rect 129 44 140 78
rect 174 44 182 78
rect 129 32 182 44
<< pdiff >>
rect 36 1018 89 1030
rect 36 984 44 1018
rect 78 984 89 1018
rect 36 950 89 984
rect 36 916 44 950
rect 78 916 89 950
rect 36 882 89 916
rect 36 848 44 882
rect 78 848 89 882
rect 36 814 89 848
rect 36 780 44 814
rect 78 780 89 814
rect 36 746 89 780
rect 36 712 44 746
rect 78 712 89 746
rect 36 678 89 712
rect 36 644 44 678
rect 78 644 89 678
rect 36 610 89 644
rect 36 576 44 610
rect 78 576 89 610
rect 36 542 89 576
rect 36 508 44 542
rect 78 508 89 542
rect 36 430 89 508
rect 139 1018 192 1030
rect 139 984 150 1018
rect 184 984 192 1018
rect 139 950 192 984
rect 139 916 150 950
rect 184 916 192 950
rect 139 882 192 916
rect 139 848 150 882
rect 184 848 192 882
rect 139 814 192 848
rect 139 780 150 814
rect 184 780 192 814
rect 139 746 192 780
rect 139 712 150 746
rect 184 712 192 746
rect 139 678 192 712
rect 139 644 150 678
rect 184 644 192 678
rect 139 610 192 644
rect 139 576 150 610
rect 184 576 192 610
rect 139 542 192 576
rect 139 508 150 542
rect 184 508 192 542
rect 139 430 192 508
<< ndiffc >>
rect 34 180 68 214
rect 34 112 68 146
rect 34 44 68 78
rect 140 180 174 214
rect 140 112 174 146
rect 140 44 174 78
<< pdiffc >>
rect 44 984 78 1018
rect 44 916 78 950
rect 44 848 78 882
rect 44 780 78 814
rect 44 712 78 746
rect 44 644 78 678
rect 44 576 78 610
rect 44 508 78 542
rect 150 984 184 1018
rect 150 916 184 950
rect 150 848 184 882
rect 150 780 184 814
rect 150 712 184 746
rect 150 644 184 678
rect 150 576 184 610
rect 150 508 184 542
<< psubdiff >>
rect 258 208 292 232
rect 258 90 292 174
rect 258 32 292 56
<< nsubdiff >>
rect 258 937 292 999
rect 258 869 292 903
rect 258 801 292 835
rect 258 733 292 767
rect 258 665 292 699
rect 258 597 292 631
rect 258 529 292 563
rect 258 461 292 495
<< psubdiffcont >>
rect 258 174 292 208
rect 258 56 292 90
<< nsubdiffcont >>
rect 258 903 292 937
rect 258 835 292 869
rect 258 767 292 801
rect 258 699 292 733
rect 258 631 292 665
rect 258 563 292 597
rect 258 495 292 529
<< poly >>
rect 89 1030 139 1062
rect 89 398 139 430
rect 80 382 146 398
rect 80 348 96 382
rect 130 348 146 382
rect 80 314 146 348
rect 80 280 96 314
rect 130 280 146 314
rect 80 264 146 280
rect 79 232 129 264
rect 79 0 129 32
<< polycont >>
rect 96 348 130 382
rect 96 280 130 314
<< locali >>
rect 44 1018 78 1034
rect 44 950 78 984
rect 44 882 78 916
rect 44 840 78 848
rect 44 762 78 780
rect 44 684 78 712
rect 44 610 78 644
rect 44 542 78 571
rect 150 1018 184 1034
rect 150 950 184 984
rect 150 882 184 907
rect 150 814 184 830
rect 150 746 184 753
rect 150 710 184 712
rect 150 632 184 644
rect 150 554 184 576
rect 150 492 184 508
rect 258 987 292 999
rect 258 937 292 953
rect 258 869 292 873
rect 258 827 292 835
rect 258 747 292 767
rect 258 667 292 699
rect 258 597 292 631
rect 258 529 292 553
rect 258 461 292 473
rect 96 382 130 398
rect 96 314 130 348
rect 96 264 130 276
rect 34 216 68 230
rect 34 146 68 180
rect 34 78 68 112
rect 34 28 68 44
rect 140 216 174 230
rect 140 146 174 180
rect 140 78 174 112
rect 140 28 174 44
rect 258 216 292 232
rect 258 90 292 174
rect 258 32 292 44
<< viali >>
rect 44 814 78 840
rect 44 806 78 814
rect 44 746 78 762
rect 44 728 78 746
rect 44 678 78 684
rect 44 650 78 678
rect 44 576 78 605
rect 44 571 78 576
rect 44 508 78 526
rect 44 492 78 508
rect 150 984 184 1018
rect 150 916 184 941
rect 150 907 184 916
rect 150 848 184 864
rect 150 830 184 848
rect 150 780 184 787
rect 150 753 184 780
rect 150 678 184 710
rect 150 676 184 678
rect 150 610 184 632
rect 150 598 184 610
rect 150 542 184 554
rect 150 520 184 542
rect 258 953 292 987
rect 258 903 292 907
rect 258 873 292 903
rect 258 801 292 827
rect 258 793 292 801
rect 258 733 292 747
rect 258 713 292 733
rect 258 665 292 667
rect 258 633 292 665
rect 258 563 292 587
rect 258 553 292 563
rect 258 495 292 507
rect 258 473 292 495
rect 96 348 130 382
rect 96 280 130 310
rect 96 276 130 280
rect 34 214 68 216
rect 34 182 68 214
rect 34 44 68 78
rect 140 214 174 216
rect 140 182 174 214
rect 140 44 174 78
rect 258 208 292 216
rect 258 182 292 208
rect 258 56 292 78
rect 258 44 292 56
<< metal1 >>
rect 144 1018 298 1030
rect 144 984 150 1018
rect 184 987 298 1018
rect 184 984 258 987
rect 144 953 258 984
rect 292 953 298 987
rect 144 941 298 953
rect 144 907 150 941
rect 184 907 298 941
rect 144 873 258 907
rect 292 873 298 907
rect 144 864 298 873
rect 16 840 84 852
rect 16 806 44 840
rect 78 806 84 840
rect 16 762 84 806
rect 16 728 44 762
rect 78 728 84 762
rect 16 684 84 728
rect 16 650 44 684
rect 78 650 84 684
rect 16 605 84 650
rect 16 571 44 605
rect 78 571 84 605
rect 16 526 84 571
rect 16 492 44 526
rect 78 492 84 526
rect 16 480 84 492
rect 16 473 77 480
tri 77 473 84 480 nw
rect 144 830 150 864
rect 184 830 298 864
rect 144 827 298 830
rect 144 793 258 827
rect 292 793 298 827
rect 144 787 298 793
rect 144 753 150 787
rect 184 753 298 787
rect 144 747 298 753
rect 144 713 258 747
rect 292 713 298 747
rect 144 710 298 713
rect 144 676 150 710
rect 184 676 298 710
rect 144 667 298 676
rect 144 633 258 667
rect 292 633 298 667
rect 144 632 298 633
rect 144 598 150 632
rect 184 598 298 632
rect 144 587 298 598
rect 144 554 258 587
rect 144 520 150 554
rect 184 553 258 554
rect 292 553 298 587
rect 184 520 298 553
rect 144 507 298 520
rect 144 473 258 507
rect 292 473 298 507
rect 16 461 65 473
tri 65 461 77 473 nw
rect 144 461 298 473
rect 16 228 62 461
tri 62 458 65 461 nw
rect 90 382 136 394
rect 90 348 96 382
rect 130 348 136 382
rect 90 310 136 348
rect 90 276 96 310
rect 130 276 136 310
rect 90 264 136 276
tri 62 228 74 240 sw
rect 16 216 74 228
rect 16 182 34 216
rect 68 182 74 216
rect 16 78 74 182
rect 16 44 34 78
rect 68 44 74 78
rect 16 32 74 44
rect 134 216 298 228
rect 134 182 140 216
rect 174 182 258 216
rect 292 182 298 216
rect 134 78 298 182
rect 134 44 140 78
rect 174 44 258 78
rect 292 44 298 78
rect 134 32 298 44
use sky130_fd_pr__pfet_01v8__example_55959141808595  sky130_fd_pr__pfet_01v8__example_55959141808595_0
timestamp 1619729480
transform 1 0 89 0 -1 1030
box -28 0 78 267
use sky130_fd_pr__nfet_01v8__example_5595914180825  sky130_fd_pr__nfet_01v8__example_5595914180825_0
timestamp 1619729480
transform 1 0 79 0 1 32
box -28 0 78 97
<< labels >>
flabel metal1 s 106 315 124 361 3 FreeSans 200 0 0 0 IN
flabel metal1 s 179 85 234 197 3 FreeSans 200 0 0 0 VGND
flabel metal1 s 193 595 249 786 3 FreeSans 200 0 0 0 VPWR
flabel metal1 s 22 293 45 372 3 FreeSans 200 0 0 0 OUT
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 13973544
string GDS_START 13968610
<< end >>
