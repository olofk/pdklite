magic
tech sky130A
magscale 1 2
timestamp 1619729571
<< checkpaint >>
rect -1298 -1308 2034 1852
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 26 -17 60 17
<< scnmos >>
rect 81 47 111 177
rect 165 47 195 177
rect 353 47 383 177
rect 437 47 467 177
rect 543 47 573 177
rect 627 47 657 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 353 297 383 497
rect 425 297 455 497
rect 549 297 579 497
rect 621 297 651 497
<< ndiff >>
rect 29 161 81 177
rect 29 127 37 161
rect 71 127 81 161
rect 29 93 81 127
rect 29 59 37 93
rect 71 59 81 93
rect 29 47 81 59
rect 111 136 165 177
rect 111 102 121 136
rect 155 102 165 136
rect 111 47 165 102
rect 195 93 247 177
rect 195 59 205 93
rect 239 59 247 93
rect 195 47 247 59
rect 301 95 353 177
rect 301 61 309 95
rect 343 61 353 95
rect 301 47 353 61
rect 383 163 437 177
rect 383 129 393 163
rect 427 129 437 163
rect 383 47 437 129
rect 467 163 543 177
rect 467 129 494 163
rect 528 129 543 163
rect 467 95 543 129
rect 467 61 494 95
rect 528 61 543 95
rect 467 47 543 61
rect 573 89 627 177
rect 573 55 583 89
rect 617 55 627 89
rect 573 47 627 55
rect 657 163 709 177
rect 657 129 667 163
rect 701 129 709 163
rect 657 95 709 129
rect 657 61 667 95
rect 701 61 709 95
rect 657 47 709 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 477 167 497
rect 113 443 123 477
rect 157 443 167 477
rect 113 409 167 443
rect 113 375 123 409
rect 157 375 167 409
rect 113 341 167 375
rect 113 307 123 341
rect 157 307 167 341
rect 113 297 167 307
rect 197 477 353 497
rect 197 443 215 477
rect 249 443 309 477
rect 343 443 353 477
rect 197 409 353 443
rect 197 375 215 409
rect 249 375 309 409
rect 343 375 353 409
rect 197 297 353 375
rect 383 297 425 497
rect 455 477 549 497
rect 455 443 465 477
rect 499 443 549 477
rect 455 409 549 443
rect 455 375 465 409
rect 499 375 549 409
rect 455 341 549 375
rect 455 307 465 341
rect 499 307 549 341
rect 455 297 549 307
rect 579 297 621 497
rect 651 477 707 497
rect 651 443 661 477
rect 695 443 707 477
rect 651 409 707 443
rect 651 375 661 409
rect 695 375 707 409
rect 651 297 707 375
<< ndiffc >>
rect 37 127 71 161
rect 37 59 71 93
rect 121 102 155 136
rect 205 59 239 93
rect 309 61 343 95
rect 393 129 427 163
rect 494 129 528 163
rect 494 61 528 95
rect 583 55 617 89
rect 667 129 701 163
rect 667 61 701 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 443 157 477
rect 123 375 157 409
rect 123 307 157 341
rect 215 443 249 477
rect 309 443 343 477
rect 215 375 249 409
rect 309 375 343 409
rect 465 443 499 477
rect 465 375 499 409
rect 465 307 499 341
rect 661 443 695 477
rect 661 375 695 409
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 353 497 383 523
rect 425 497 455 523
rect 549 497 579 523
rect 621 497 651 523
rect 83 265 113 297
rect 167 265 197 297
rect 353 265 383 297
rect 81 249 254 265
rect 81 215 210 249
rect 244 215 254 249
rect 81 199 254 215
rect 298 249 383 265
rect 298 215 308 249
rect 342 215 383 249
rect 298 199 383 215
rect 425 265 455 297
rect 549 265 579 297
rect 425 249 479 265
rect 425 215 435 249
rect 469 215 479 249
rect 425 199 479 215
rect 521 249 579 265
rect 521 215 535 249
rect 569 215 579 249
rect 521 199 579 215
rect 621 265 651 297
rect 621 249 689 265
rect 621 215 641 249
rect 675 215 689 249
rect 621 199 689 215
rect 81 177 111 199
rect 165 177 195 199
rect 353 177 383 199
rect 437 177 467 199
rect 543 177 573 199
rect 627 177 657 199
rect 81 21 111 47
rect 165 21 195 47
rect 353 21 383 47
rect 437 21 467 47
rect 543 21 573 47
rect 627 21 657 47
<< polycont >>
rect 210 215 244 249
rect 308 215 342 249
rect 435 215 469 249
rect 535 215 569 249
rect 641 215 675 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 23 477 73 527
rect 23 443 39 477
rect 23 409 73 443
rect 23 375 39 409
rect 23 341 73 375
rect 23 307 39 341
rect 23 289 73 307
rect 118 477 161 493
rect 118 443 123 477
rect 157 443 161 477
rect 118 409 161 443
rect 118 375 123 409
rect 157 375 161 409
rect 199 477 359 527
rect 199 443 215 477
rect 249 443 309 477
rect 343 443 359 477
rect 199 409 359 443
rect 199 375 215 409
rect 249 375 309 409
rect 343 375 359 409
rect 438 477 515 493
rect 438 443 465 477
rect 499 443 515 477
rect 438 409 515 443
rect 438 375 465 409
rect 499 375 515 409
rect 118 341 161 375
rect 438 341 515 375
rect 118 307 123 341
rect 157 307 161 341
rect 37 161 71 177
rect 37 93 71 127
rect 118 136 161 307
rect 195 307 465 341
rect 499 307 515 341
rect 580 323 620 481
rect 654 477 718 527
rect 654 443 661 477
rect 695 443 718 477
rect 654 409 718 443
rect 654 375 661 409
rect 695 375 718 409
rect 654 359 718 375
rect 195 299 515 307
rect 195 249 251 299
rect 549 289 620 323
rect 549 265 585 289
rect 195 215 210 249
rect 244 215 251 249
rect 287 249 358 265
rect 287 215 308 249
rect 342 215 358 249
rect 392 249 485 265
rect 392 215 435 249
rect 469 215 485 249
rect 519 249 585 265
rect 654 255 718 323
rect 519 215 535 249
rect 569 215 585 249
rect 619 249 718 255
rect 619 215 641 249
rect 675 215 718 249
rect 195 179 251 215
rect 195 163 443 179
rect 512 165 718 173
rect 195 143 393 163
rect 118 102 121 136
rect 155 102 161 136
rect 370 129 393 143
rect 427 129 443 163
rect 478 163 718 165
rect 478 129 494 163
rect 528 139 667 163
rect 528 129 546 139
rect 118 73 161 102
rect 205 93 241 109
rect 478 95 546 129
rect 651 129 667 139
rect 701 129 718 163
rect 37 17 71 59
rect 239 59 241 93
rect 293 61 309 95
rect 343 61 494 95
rect 528 61 546 95
rect 293 59 546 61
rect 583 89 617 105
rect 205 17 241 59
rect 651 95 718 129
rect 651 61 667 95
rect 701 61 718 95
rect 651 56 718 61
rect 583 17 617 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 580 357 614 391 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 118 425 152 459 0 FreeSans 400 0 0 0 X
port 9 nsew signal output
flabel locali s 304 221 338 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 672 221 706 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 396 221 430 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel pwell s 26 -17 60 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 26 527 60 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 26 -17 60 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 26 527 60 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o22a_2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 2214766
string GDS_START 2208172
string path 0.000 0.000 18.400 0.000 
<< end >>
