magic
tech sky130A
magscale 1 2
timestamp 1619729575
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 35 -12 57 12
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
rlabel metal1 s 0 -48 368 48 8 VGND
port 1 nsew ground bidirectional abutment
rlabel pwell s 35 -12 57 12 8 VNB
port 2 nsew ground bidirectional
rlabel nwell s -38 261 406 582 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 0 496 368 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE SPACER
string FIXED_BBOX 0 0 368 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 4092970
string GDS_START 4091358
<< end >>
