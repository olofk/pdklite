magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1285 -760 1405 1761
<< labels >>
flabel comment s 145 500 145 500 0 FreeSans 300 0 0 0 D
flabel comment s -25 500 -25 500 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 3491326
string GDS_START 3490558
<< end >>
