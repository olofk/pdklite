magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1204 -1401 3122 2392
<< nwell >>
rect 818 1030 1139 1132
rect 818 598 1862 1030
<< pwell >>
rect 90 -141 600 -107
rect 905 -141 1744 -107
<< mvnmos >>
rect 111 703 211 1003
rect 267 703 367 1003
rect 423 703 523 1003
rect 579 703 679 1003
rect 96 410 396 510
rect 526 359 826 459
rect 956 359 1256 459
rect 1386 359 1686 459
<< mvpmos >>
rect 884 893 1024 1013
rect 884 717 1024 837
rect 1175 664 1275 964
rect 1331 664 1431 964
rect 1487 664 1587 964
rect 1643 664 1743 964
<< mvnnmos >>
rect 735 -33 915 167
rect 971 -33 1151 167
rect 1328 -33 1508 167
rect 1564 -33 1744 167
<< nmoslvt >>
rect 196 13 226 213
rect 282 13 312 213
rect 368 13 398 213
rect 454 13 484 213
<< ndiff >>
rect 143 195 196 213
rect 143 161 151 195
rect 185 161 196 195
rect 143 127 196 161
rect 143 93 151 127
rect 185 93 196 127
rect 143 59 196 93
rect 143 25 151 59
rect 185 25 196 59
rect 143 13 196 25
rect 226 195 282 213
rect 226 161 237 195
rect 271 161 282 195
rect 226 127 282 161
rect 226 93 237 127
rect 271 93 282 127
rect 226 59 282 93
rect 226 25 237 59
rect 271 25 282 59
rect 226 13 282 25
rect 312 195 368 213
rect 312 161 323 195
rect 357 161 368 195
rect 312 127 368 161
rect 312 93 323 127
rect 357 93 368 127
rect 312 59 368 93
rect 312 25 323 59
rect 357 25 368 59
rect 312 13 368 25
rect 398 195 454 213
rect 398 161 409 195
rect 443 161 454 195
rect 398 127 454 161
rect 398 93 409 127
rect 443 93 454 127
rect 398 59 454 93
rect 398 25 409 59
rect 443 25 454 59
rect 398 13 454 25
rect 484 195 537 213
rect 484 161 495 195
rect 529 161 537 195
rect 484 127 537 161
rect 484 93 495 127
rect 529 93 537 127
rect 484 59 537 93
rect 484 25 495 59
rect 529 25 537 59
rect 484 13 537 25
<< mvndiff >>
rect 58 991 111 1003
rect 58 957 66 991
rect 100 957 111 991
rect 58 923 111 957
rect 58 889 66 923
rect 100 889 111 923
rect 58 855 111 889
rect 58 821 66 855
rect 100 821 111 855
rect 58 787 111 821
rect 58 753 66 787
rect 100 753 111 787
rect 58 703 111 753
rect 211 991 267 1003
rect 211 957 222 991
rect 256 957 267 991
rect 211 923 267 957
rect 211 889 222 923
rect 256 889 267 923
rect 211 855 267 889
rect 211 821 222 855
rect 256 821 267 855
rect 211 787 267 821
rect 211 753 222 787
rect 256 753 267 787
rect 211 703 267 753
rect 367 991 423 1003
rect 367 957 378 991
rect 412 957 423 991
rect 367 923 423 957
rect 367 889 378 923
rect 412 889 423 923
rect 367 855 423 889
rect 367 821 378 855
rect 412 821 423 855
rect 367 787 423 821
rect 367 753 378 787
rect 412 753 423 787
rect 367 703 423 753
rect 523 991 579 1003
rect 523 957 534 991
rect 568 957 579 991
rect 523 923 579 957
rect 523 889 534 923
rect 568 889 579 923
rect 523 855 579 889
rect 523 821 534 855
rect 568 821 579 855
rect 523 787 579 821
rect 523 753 534 787
rect 568 753 579 787
rect 523 703 579 753
rect 679 991 732 1003
rect 679 957 690 991
rect 724 957 732 991
rect 679 923 732 957
rect 679 889 690 923
rect 724 889 732 923
rect 679 855 732 889
rect 679 821 690 855
rect 724 821 732 855
rect 679 787 732 821
rect 679 753 690 787
rect 724 753 732 787
rect 679 703 732 753
rect 96 555 396 563
rect 96 521 108 555
rect 142 521 176 555
rect 210 521 244 555
rect 278 521 312 555
rect 346 521 396 555
rect 96 510 396 521
rect 526 504 826 512
rect 526 470 538 504
rect 572 470 606 504
rect 640 470 674 504
rect 708 470 742 504
rect 776 470 826 504
rect 526 459 826 470
rect 956 504 1256 512
rect 956 470 968 504
rect 1002 470 1036 504
rect 1070 470 1104 504
rect 1138 470 1172 504
rect 1206 470 1256 504
rect 1386 504 1686 512
rect 956 459 1256 470
rect 96 399 396 410
rect 96 365 108 399
rect 142 365 176 399
rect 210 365 244 399
rect 278 365 312 399
rect 346 365 396 399
rect 96 357 396 365
rect 1386 470 1398 504
rect 1432 470 1466 504
rect 1500 470 1534 504
rect 1568 470 1602 504
rect 1636 470 1686 504
rect 1386 459 1686 470
rect 526 348 826 359
rect 526 314 538 348
rect 572 314 606 348
rect 640 314 674 348
rect 708 314 742 348
rect 776 314 826 348
rect 526 306 826 314
rect 956 348 1256 359
rect 956 314 968 348
rect 1002 314 1036 348
rect 1070 314 1104 348
rect 1138 314 1172 348
rect 1206 314 1256 348
rect 1386 348 1686 359
rect 956 306 1256 314
rect 1386 314 1398 348
rect 1432 314 1466 348
rect 1500 314 1534 348
rect 1568 314 1602 348
rect 1636 314 1686 348
rect 1386 306 1686 314
rect 682 149 735 167
rect 682 115 690 149
rect 724 115 735 149
rect 682 81 735 115
rect 682 47 690 81
rect 724 47 735 81
rect 682 13 735 47
rect 682 -21 690 13
rect 724 -21 735 13
rect 682 -33 735 -21
rect 915 149 971 167
rect 915 115 926 149
rect 960 115 971 149
rect 915 81 971 115
rect 915 47 926 81
rect 960 47 971 81
rect 915 13 971 47
rect 915 -21 926 13
rect 960 -21 971 13
rect 915 -33 971 -21
rect 1151 149 1204 167
rect 1151 115 1162 149
rect 1196 115 1204 149
rect 1151 81 1204 115
rect 1151 47 1162 81
rect 1196 47 1204 81
rect 1151 13 1204 47
rect 1151 -21 1162 13
rect 1196 -21 1204 13
rect 1151 -33 1204 -21
rect 1275 155 1328 167
rect 1275 121 1283 155
rect 1317 121 1328 155
rect 1275 87 1328 121
rect 1275 53 1283 87
rect 1317 53 1328 87
rect 1275 19 1328 53
rect 1275 -15 1283 19
rect 1317 -15 1328 19
rect 1275 -33 1328 -15
rect 1508 155 1564 167
rect 1508 121 1519 155
rect 1553 121 1564 155
rect 1508 87 1564 121
rect 1508 53 1519 87
rect 1553 53 1564 87
rect 1508 19 1564 53
rect 1508 -15 1519 19
rect 1553 -15 1564 19
rect 1508 -33 1564 -15
rect 1744 155 1797 167
rect 1744 121 1755 155
rect 1789 121 1797 155
rect 1744 87 1797 121
rect 1744 53 1755 87
rect 1789 53 1797 87
rect 1744 19 1797 53
rect 1744 -15 1755 19
rect 1789 -15 1797 19
rect 1744 -33 1797 -15
<< mvpdiff >>
rect 884 1058 1024 1066
rect 884 1024 896 1058
rect 930 1024 964 1058
rect 998 1024 1024 1058
rect 884 1013 1024 1024
rect 1122 952 1175 964
rect 1122 918 1130 952
rect 1164 918 1175 952
rect 884 882 1024 893
rect 884 848 896 882
rect 930 848 964 882
rect 998 848 1024 882
rect 884 837 1024 848
rect 1122 884 1175 918
rect 1122 850 1130 884
rect 1164 850 1175 884
rect 1122 816 1175 850
rect 1122 782 1130 816
rect 1164 782 1175 816
rect 1122 748 1175 782
rect 884 706 1024 717
rect 884 672 896 706
rect 930 672 964 706
rect 998 672 1024 706
rect 884 664 1024 672
rect 1122 714 1130 748
rect 1164 714 1175 748
rect 1122 664 1175 714
rect 1275 952 1331 964
rect 1275 918 1286 952
rect 1320 918 1331 952
rect 1275 884 1331 918
rect 1275 850 1286 884
rect 1320 850 1331 884
rect 1275 816 1331 850
rect 1275 782 1286 816
rect 1320 782 1331 816
rect 1275 748 1331 782
rect 1275 714 1286 748
rect 1320 714 1331 748
rect 1275 664 1331 714
rect 1431 952 1487 964
rect 1431 918 1442 952
rect 1476 918 1487 952
rect 1431 884 1487 918
rect 1431 850 1442 884
rect 1476 850 1487 884
rect 1431 816 1487 850
rect 1431 782 1442 816
rect 1476 782 1487 816
rect 1431 748 1487 782
rect 1431 714 1442 748
rect 1476 714 1487 748
rect 1431 664 1487 714
rect 1587 952 1643 964
rect 1587 918 1598 952
rect 1632 918 1643 952
rect 1587 884 1643 918
rect 1587 850 1598 884
rect 1632 850 1643 884
rect 1587 816 1643 850
rect 1587 782 1598 816
rect 1632 782 1643 816
rect 1587 748 1643 782
rect 1587 714 1598 748
rect 1632 714 1643 748
rect 1587 664 1643 714
rect 1743 952 1796 964
rect 1743 918 1754 952
rect 1788 918 1796 952
rect 1743 884 1796 918
rect 1743 850 1754 884
rect 1788 850 1796 884
rect 1743 816 1796 850
rect 1743 782 1754 816
rect 1788 782 1796 816
rect 1743 748 1796 782
rect 1743 714 1754 748
rect 1788 714 1796 748
rect 1743 664 1796 714
<< ndiffc >>
rect 151 161 185 195
rect 151 93 185 127
rect 151 25 185 59
rect 237 161 271 195
rect 237 93 271 127
rect 237 25 271 59
rect 323 161 357 195
rect 323 93 357 127
rect 323 25 357 59
rect 409 161 443 195
rect 409 93 443 127
rect 409 25 443 59
rect 495 161 529 195
rect 495 93 529 127
rect 495 25 529 59
<< mvndiffc >>
rect 66 957 100 991
rect 66 889 100 923
rect 66 821 100 855
rect 66 753 100 787
rect 222 957 256 991
rect 222 889 256 923
rect 222 821 256 855
rect 222 753 256 787
rect 378 957 412 991
rect 378 889 412 923
rect 378 821 412 855
rect 378 753 412 787
rect 534 957 568 991
rect 534 889 568 923
rect 534 821 568 855
rect 534 753 568 787
rect 690 957 724 991
rect 690 889 724 923
rect 690 821 724 855
rect 690 753 724 787
rect 108 521 142 555
rect 176 521 210 555
rect 244 521 278 555
rect 312 521 346 555
rect 538 470 572 504
rect 606 470 640 504
rect 674 470 708 504
rect 742 470 776 504
rect 968 470 1002 504
rect 1036 470 1070 504
rect 1104 470 1138 504
rect 1172 470 1206 504
rect 108 365 142 399
rect 176 365 210 399
rect 244 365 278 399
rect 312 365 346 399
rect 1398 470 1432 504
rect 1466 470 1500 504
rect 1534 470 1568 504
rect 1602 470 1636 504
rect 538 314 572 348
rect 606 314 640 348
rect 674 314 708 348
rect 742 314 776 348
rect 968 314 1002 348
rect 1036 314 1070 348
rect 1104 314 1138 348
rect 1172 314 1206 348
rect 1398 314 1432 348
rect 1466 314 1500 348
rect 1534 314 1568 348
rect 1602 314 1636 348
rect 690 115 724 149
rect 690 47 724 81
rect 690 -21 724 13
rect 926 115 960 149
rect 926 47 960 81
rect 926 -21 960 13
rect 1162 115 1196 149
rect 1162 47 1196 81
rect 1162 -21 1196 13
rect 1283 121 1317 155
rect 1283 53 1317 87
rect 1283 -15 1317 19
rect 1519 121 1553 155
rect 1519 53 1553 87
rect 1519 -15 1553 19
rect 1755 121 1789 155
rect 1755 53 1789 87
rect 1755 -15 1789 19
<< mvpdiffc >>
rect 896 1024 930 1058
rect 964 1024 998 1058
rect 1130 918 1164 952
rect 896 848 930 882
rect 964 848 998 882
rect 1130 850 1164 884
rect 1130 782 1164 816
rect 896 672 930 706
rect 964 672 998 706
rect 1130 714 1164 748
rect 1286 918 1320 952
rect 1286 850 1320 884
rect 1286 782 1320 816
rect 1286 714 1320 748
rect 1442 918 1476 952
rect 1442 850 1476 884
rect 1442 782 1476 816
rect 1442 714 1476 748
rect 1598 918 1632 952
rect 1598 850 1632 884
rect 1598 782 1632 816
rect 1598 714 1632 748
rect 1754 918 1788 952
rect 1754 850 1788 884
rect 1754 782 1788 816
rect 1754 714 1788 748
<< psubdiff >>
rect 90 -141 114 -107
rect 148 -141 186 -107
rect 220 -141 258 -107
rect 292 -141 329 -107
rect 363 -141 400 -107
rect 434 -141 471 -107
rect 505 -141 542 -107
rect 576 -141 600 -107
<< mvpsubdiff >>
rect 905 -141 929 -107
rect 963 -141 998 -107
rect 1032 -141 1067 -107
rect 1101 -141 1136 -107
rect 1170 -141 1205 -107
rect 1239 -141 1274 -107
rect 1308 -141 1343 -107
rect 1377 -141 1412 -107
rect 1446 -141 1481 -107
rect 1515 -141 1550 -107
rect 1584 -141 1618 -107
rect 1652 -141 1686 -107
rect 1720 -141 1744 -107
<< psubdiffcont >>
rect 114 -141 148 -107
rect 186 -141 220 -107
rect 258 -141 292 -107
rect 329 -141 363 -107
rect 400 -141 434 -107
rect 471 -141 505 -107
rect 542 -141 576 -107
<< mvpsubdiffcont >>
rect 929 -141 963 -107
rect 998 -141 1032 -107
rect 1067 -141 1101 -107
rect 1136 -141 1170 -107
rect 1205 -141 1239 -107
rect 1274 -141 1308 -107
rect 1343 -141 1377 -107
rect 1412 -141 1446 -107
rect 1481 -141 1515 -107
rect 1550 -141 1584 -107
rect 1618 -141 1652 -107
rect 1686 -141 1720 -107
<< poly >>
rect 111 1003 211 1035
rect 267 1003 367 1035
rect 423 1003 523 1035
rect 579 1003 679 1035
rect 786 1013 852 1022
rect 786 1006 884 1013
rect 786 972 802 1006
rect 836 972 884 1006
rect 786 938 884 972
rect 786 904 802 938
rect 836 904 884 938
rect 786 893 884 904
rect 1024 893 1056 1013
rect 1175 964 1275 996
rect 1331 964 1431 996
rect 1487 964 1587 996
rect 1643 964 1743 996
rect 786 888 852 893
rect 786 837 852 842
rect 786 826 884 837
rect 786 792 802 826
rect 836 792 884 826
rect 786 758 884 792
rect 786 724 802 758
rect 836 724 884 758
rect 786 717 884 724
rect 1024 717 1056 837
rect 786 708 852 717
rect 111 671 211 703
rect 267 671 367 703
rect 423 671 523 703
rect 111 655 523 671
rect 111 621 127 655
rect 161 621 196 655
rect 230 621 265 655
rect 299 621 334 655
rect 368 621 403 655
rect 437 621 473 655
rect 507 621 523 655
rect 111 605 523 621
rect 579 671 679 703
rect 579 655 713 671
rect 579 621 595 655
rect 629 621 663 655
rect 697 621 713 655
rect 579 605 713 621
rect 1175 632 1275 664
rect 1331 632 1431 664
rect 1487 632 1587 664
rect 1175 616 1587 632
rect 1175 582 1191 616
rect 1225 582 1261 616
rect 1295 582 1330 616
rect 1364 582 1399 616
rect 1433 582 1468 616
rect 1502 582 1537 616
rect 1571 582 1587 616
rect 1175 566 1587 582
rect 1643 632 1743 664
rect 1643 616 1778 632
rect 1643 582 1659 616
rect 1693 582 1728 616
rect 1762 582 1778 616
rect 1643 566 1778 582
rect 64 410 96 510
rect 396 494 494 510
rect 396 460 444 494
rect 478 460 494 494
rect 396 459 494 460
rect 858 494 924 510
rect 858 460 874 494
rect 908 460 924 494
rect 858 459 924 460
rect 1288 461 1354 477
rect 1288 459 1304 461
rect 396 410 526 459
rect 428 409 526 410
rect 428 375 444 409
rect 478 375 526 409
rect 428 359 526 375
rect 826 409 956 459
rect 826 375 874 409
rect 908 375 956 409
rect 826 359 956 375
rect 1256 427 1304 459
rect 1338 459 1354 461
rect 1338 427 1386 459
rect 1256 393 1386 427
rect 1256 359 1304 393
rect 1338 359 1386 393
rect 1686 359 1718 459
rect 1288 343 1354 359
rect 178 289 312 305
rect 178 255 194 289
rect 228 255 262 289
rect 296 255 312 289
rect 178 239 312 255
rect 362 289 496 305
rect 362 255 378 289
rect 412 255 446 289
rect 480 255 496 289
rect 362 239 496 255
rect 735 243 1744 259
rect 196 213 226 239
rect 282 213 312 239
rect 368 213 398 239
rect 454 213 484 239
rect 735 209 1232 243
rect 1266 209 1309 243
rect 1343 209 1386 243
rect 1420 209 1463 243
rect 1497 209 1540 243
rect 1574 209 1617 243
rect 1651 209 1694 243
rect 1728 209 1744 243
rect 735 193 1744 209
rect 735 167 915 193
rect 971 167 1151 193
rect 1328 167 1508 193
rect 1564 167 1744 193
rect 196 -19 226 13
rect 282 -19 312 13
rect 368 -19 398 13
rect 454 -19 484 13
rect 735 -65 915 -33
rect 971 -65 1151 -33
rect 1328 -65 1508 -33
rect 1564 -65 1744 -33
<< polycont >>
rect 802 972 836 1006
rect 802 904 836 938
rect 802 792 836 826
rect 802 724 836 758
rect 127 621 161 655
rect 196 621 230 655
rect 265 621 299 655
rect 334 621 368 655
rect 403 621 437 655
rect 473 621 507 655
rect 595 621 629 655
rect 663 621 697 655
rect 1191 582 1225 616
rect 1261 582 1295 616
rect 1330 582 1364 616
rect 1399 582 1433 616
rect 1468 582 1502 616
rect 1537 582 1571 616
rect 1659 582 1693 616
rect 1728 582 1762 616
rect 444 460 478 494
rect 874 460 908 494
rect 444 375 478 409
rect 874 375 908 409
rect 1304 427 1338 461
rect 1304 359 1338 393
rect 194 255 228 289
rect 262 255 296 289
rect 378 255 412 289
rect 446 255 480 289
rect 1232 209 1266 243
rect 1309 209 1343 243
rect 1386 209 1420 243
rect 1463 209 1497 243
rect 1540 209 1574 243
rect 1617 209 1651 243
rect 1694 209 1728 243
<< locali >>
rect 914 1058 952 1059
rect 930 1025 952 1058
rect 880 1024 896 1025
rect 930 1024 964 1025
rect 998 1024 1014 1058
rect 66 1005 100 1007
rect 66 933 100 957
rect 66 855 100 889
rect 66 787 100 821
rect 222 991 256 1007
rect 222 923 256 957
rect 222 855 256 889
rect 222 787 256 821
rect 66 737 100 753
rect 219 753 222 771
rect 378 1005 412 1007
rect 378 933 412 957
rect 378 855 412 889
rect 378 787 412 821
rect 256 753 257 771
rect 219 737 257 753
rect 534 991 568 1007
rect 534 923 568 957
rect 534 855 568 889
rect 534 787 568 821
rect 657 1005 724 1007
rect 691 991 724 1005
rect 802 1006 836 1022
rect 657 957 690 971
rect 657 933 724 957
rect 836 972 870 975
rect 832 941 870 972
rect 691 923 724 933
rect 657 889 690 899
rect 657 855 724 889
rect 802 938 836 941
rect 802 888 836 904
rect 1130 911 1164 918
rect 657 821 690 855
rect 880 848 896 882
rect 930 848 949 882
rect 998 848 1021 882
rect 657 787 724 821
rect 378 737 412 753
rect 568 753 575 771
rect 537 737 575 753
rect 657 753 690 787
rect 657 737 724 753
rect 802 829 836 842
rect 802 758 836 792
rect 802 708 836 723
rect 1130 816 1164 850
rect 1130 748 1164 782
rect 880 672 883 706
rect 930 672 955 706
rect 998 672 1014 706
rect 1130 698 1164 714
rect 1286 952 1320 968
rect 1286 884 1320 918
rect 1286 816 1320 850
rect 1286 748 1320 749
rect 1286 711 1320 714
rect 1442 911 1476 918
rect 1442 816 1476 850
rect 1442 748 1476 782
rect 1442 698 1476 714
rect 1598 952 1632 968
rect 1598 884 1632 918
rect 1598 816 1632 850
rect 1598 748 1632 749
rect 1598 711 1632 714
rect 1754 911 1788 918
rect 1754 816 1788 850
rect 1754 748 1788 782
rect 1754 698 1788 714
rect 111 621 123 655
rect 161 621 196 655
rect 246 621 265 655
rect 299 621 300 655
rect 368 621 388 655
rect 437 621 473 655
rect 510 621 523 655
rect 579 621 591 655
rect 629 621 663 655
rect 697 621 713 655
rect 1175 582 1187 616
rect 1225 582 1261 616
rect 1310 582 1330 616
rect 1364 582 1365 616
rect 1433 582 1453 616
rect 1502 582 1537 616
rect 1575 582 1587 616
rect 1643 582 1659 616
rect 1693 582 1728 616
rect 1762 610 1778 616
rect 1767 582 1778 610
rect 142 521 165 555
rect 210 521 240 555
rect 278 521 312 555
rect 348 521 362 555
rect 1733 538 1767 576
rect 444 494 478 510
rect 406 442 444 476
rect 522 470 538 504
rect 572 470 606 504
rect 640 470 674 504
rect 720 470 742 504
rect 874 494 908 510
rect 444 409 478 442
rect 142 365 165 399
rect 210 365 240 399
rect 278 365 312 399
rect 348 365 362 399
rect 444 359 478 375
rect 952 470 968 504
rect 1002 470 1036 504
rect 1082 470 1104 504
rect 1155 470 1172 504
rect 874 425 908 460
rect 1304 461 1338 477
rect 1382 470 1398 504
rect 1447 470 1466 504
rect 1522 470 1534 504
rect 1597 470 1602 504
rect 1636 470 1637 504
rect 1304 425 1338 427
rect 908 391 946 425
rect 1302 393 1340 425
rect 1302 391 1304 393
rect 874 359 908 375
rect 1338 391 1340 393
rect 522 314 538 348
rect 572 314 606 348
rect 640 314 674 348
rect 723 314 742 348
rect 952 314 968 348
rect 1003 314 1036 348
rect 1078 314 1104 348
rect 1153 314 1172 348
rect 1304 343 1338 359
rect 1382 314 1398 348
rect 1447 314 1466 348
rect 1522 314 1534 348
rect 1597 314 1602 348
rect 1636 314 1637 348
rect 178 289 199 301
rect 233 289 271 301
rect 178 255 194 289
rect 233 267 262 289
rect 305 267 312 301
rect 228 255 262 267
rect 296 255 312 267
rect 362 255 378 289
rect 414 255 446 289
rect 486 255 496 289
rect 724 220 762 254
rect 1106 220 1144 254
rect 151 195 185 211
rect 151 127 185 161
rect 151 59 185 93
rect 151 -27 185 11
rect 237 195 271 211
rect 237 127 271 140
rect 237 59 271 68
rect 237 9 271 25
rect 323 195 357 211
rect 323 127 357 161
rect 323 59 357 93
rect 151 -77 185 -61
rect 323 -37 357 1
rect 409 195 443 211
rect 409 127 443 161
rect 409 59 443 93
rect 409 -29 443 9
rect 495 195 601 211
rect 529 161 601 195
rect 495 127 601 161
rect 529 98 601 127
rect 529 64 567 98
rect 495 59 601 64
rect 529 25 601 59
rect 323 -77 357 -71
rect 495 -107 601 25
rect 690 149 752 220
rect 1116 165 1178 220
rect 1216 209 1232 243
rect 1266 209 1307 243
rect 1343 209 1382 243
rect 1420 209 1456 243
rect 1497 209 1530 243
rect 1574 209 1604 243
rect 1651 209 1678 243
rect 1728 209 1744 243
rect 1283 167 1317 171
rect 724 115 752 149
rect 690 81 752 115
rect 724 47 752 81
rect 690 13 752 47
rect 926 149 960 165
rect 926 81 960 115
rect 926 33 960 47
rect 1116 149 1196 165
rect 1116 115 1162 149
rect 1307 155 1345 167
rect 1317 133 1345 155
rect 1519 155 1553 171
rect 1755 167 1789 171
rect 1116 81 1196 115
rect 1116 47 1162 81
rect 724 -21 752 13
rect 931 13 969 33
rect 960 -1 969 13
rect 1116 13 1196 47
rect 690 -37 752 -21
rect 926 -37 960 -21
rect 1116 -21 1162 13
rect 1116 -37 1196 -21
rect 1283 87 1317 121
rect 1717 133 1755 167
rect 1519 104 1553 121
rect 1497 87 1535 104
rect 1497 70 1519 87
rect 1755 87 1789 121
rect 1283 19 1317 53
rect 1283 -31 1317 -15
rect 1519 19 1553 53
rect 1519 -31 1553 -15
rect 1755 19 1789 53
rect 1755 -31 1789 -15
rect 90 -141 114 -107
rect 148 -141 186 -107
rect 220 -141 258 -107
rect 292 -141 329 -107
rect 363 -141 400 -107
rect 434 -141 471 -107
rect 505 -141 542 -107
rect 576 -141 600 -107
rect 905 -141 929 -107
rect 963 -141 998 -107
rect 1032 -141 1067 -107
rect 1101 -141 1136 -107
rect 1170 -141 1205 -107
rect 1239 -141 1274 -107
rect 1308 -141 1343 -107
rect 1377 -141 1412 -107
rect 1446 -141 1481 -107
rect 1515 -141 1550 -107
rect 1584 -141 1618 -107
rect 1652 -141 1686 -107
rect 1720 -141 1744 -107
<< viali >>
rect 880 1058 914 1059
rect 952 1058 986 1059
rect 880 1025 896 1058
rect 896 1025 914 1058
rect 952 1025 964 1058
rect 964 1025 986 1058
rect 66 991 100 1005
rect 66 971 100 991
rect 66 923 100 933
rect 66 899 100 923
rect 185 737 219 771
rect 378 991 412 1005
rect 378 971 412 991
rect 378 923 412 933
rect 378 899 412 923
rect 257 737 291 771
rect 657 991 691 1005
rect 657 971 690 991
rect 690 971 691 991
rect 798 972 802 975
rect 802 972 832 975
rect 798 941 832 972
rect 870 941 904 975
rect 1130 952 1164 983
rect 1130 949 1164 952
rect 657 923 691 933
rect 657 899 690 923
rect 690 899 691 923
rect 1130 884 1164 911
rect 949 848 964 882
rect 964 848 983 882
rect 1021 848 1055 882
rect 1130 877 1164 884
rect 503 753 534 771
rect 534 753 537 771
rect 503 737 537 753
rect 575 737 609 771
rect 802 826 836 829
rect 802 795 836 826
rect 802 724 836 757
rect 802 723 836 724
rect 883 672 896 706
rect 896 672 917 706
rect 955 672 964 706
rect 964 672 989 706
rect 1286 782 1320 783
rect 1286 749 1320 782
rect 1286 677 1320 711
rect 1442 952 1476 983
rect 1442 949 1476 952
rect 1442 884 1476 911
rect 1442 877 1476 884
rect 1598 782 1632 783
rect 1598 749 1632 782
rect 1598 677 1632 711
rect 1754 952 1788 983
rect 1754 949 1788 952
rect 1754 884 1788 911
rect 1754 877 1788 884
rect 123 621 127 655
rect 127 621 157 655
rect 212 621 230 655
rect 230 621 246 655
rect 300 621 334 655
rect 388 621 403 655
rect 403 621 422 655
rect 476 621 507 655
rect 507 621 510 655
rect 591 621 595 655
rect 595 621 625 655
rect 663 621 697 655
rect 1187 582 1191 616
rect 1191 582 1221 616
rect 1276 582 1295 616
rect 1295 582 1310 616
rect 1365 582 1399 616
rect 1453 582 1468 616
rect 1468 582 1487 616
rect 1541 582 1571 616
rect 1571 582 1575 616
rect 1733 582 1762 610
rect 1762 582 1767 610
rect 1733 576 1767 582
rect 90 521 108 555
rect 108 521 124 555
rect 165 521 176 555
rect 176 521 199 555
rect 240 521 244 555
rect 244 521 274 555
rect 314 521 346 555
rect 346 521 348 555
rect 372 442 406 476
rect 444 460 478 476
rect 686 470 708 504
rect 708 470 720 504
rect 758 470 776 504
rect 776 470 792 504
rect 1733 504 1767 538
rect 444 442 478 460
rect 90 365 108 399
rect 108 365 124 399
rect 165 365 176 399
rect 176 365 199 399
rect 240 365 244 399
rect 244 365 274 399
rect 314 365 346 399
rect 346 365 348 399
rect 1048 470 1070 504
rect 1070 470 1082 504
rect 1121 470 1138 504
rect 1138 470 1155 504
rect 1193 470 1206 504
rect 1206 470 1227 504
rect 1413 470 1432 504
rect 1432 470 1447 504
rect 1488 470 1500 504
rect 1500 470 1522 504
rect 1563 470 1568 504
rect 1568 470 1597 504
rect 1637 470 1671 504
rect 874 409 908 425
rect 874 391 908 409
rect 946 391 980 425
rect 1268 391 1302 425
rect 1340 391 1374 425
rect 689 314 708 348
rect 708 314 723 348
rect 761 314 776 348
rect 776 314 795 348
rect 969 314 1002 348
rect 1002 314 1003 348
rect 1044 314 1070 348
rect 1070 314 1078 348
rect 1119 314 1138 348
rect 1138 314 1153 348
rect 1193 314 1206 348
rect 1206 314 1227 348
rect 1413 314 1432 348
rect 1432 314 1447 348
rect 1488 314 1500 348
rect 1500 314 1522 348
rect 1563 314 1568 348
rect 1568 314 1597 348
rect 1637 314 1671 348
rect 199 289 233 301
rect 271 289 305 301
rect 199 267 228 289
rect 228 267 233 289
rect 271 267 296 289
rect 296 267 305 289
rect 380 255 412 289
rect 412 255 414 289
rect 452 255 480 289
rect 480 255 486 289
rect 690 220 724 254
rect 762 220 796 254
rect 1072 220 1106 254
rect 1144 220 1178 254
rect 151 25 185 45
rect 151 11 185 25
rect 237 161 271 174
rect 237 140 271 161
rect 237 93 271 102
rect 237 68 271 93
rect 323 25 357 35
rect 151 -61 185 -27
rect 323 1 357 25
rect 323 -71 357 -37
rect 409 25 443 43
rect 409 9 443 25
rect 409 -63 443 -29
rect 495 93 529 98
rect 495 64 529 93
rect 567 64 601 98
rect 1307 209 1309 243
rect 1309 209 1341 243
rect 1382 209 1386 243
rect 1386 209 1416 243
rect 1456 209 1463 243
rect 1463 209 1490 243
rect 1530 209 1540 243
rect 1540 209 1564 243
rect 1604 209 1617 243
rect 1617 209 1638 243
rect 1678 209 1694 243
rect 1694 209 1712 243
rect 1273 155 1307 167
rect 1273 133 1283 155
rect 1283 133 1307 155
rect 1345 133 1379 167
rect 897 13 931 33
rect 897 -1 926 13
rect 926 -1 931 13
rect 969 -1 1003 33
rect 1683 133 1717 167
rect 1755 155 1789 167
rect 1755 133 1789 155
rect 1463 70 1497 104
rect 1535 87 1569 104
rect 1535 70 1553 87
rect 1553 70 1569 87
<< metal1 >>
tri 734 1059 740 1065 se
rect 740 1059 998 1065
tri 725 1050 734 1059 se
rect 734 1050 880 1059
rect 725 1026 880 1050
rect 725 1025 783 1026
tri 783 1025 784 1026 nw
tri 861 1025 862 1026 ne
rect 862 1025 880 1026
rect 914 1025 952 1059
rect 986 1025 998 1059
rect 60 1005 697 1017
rect 60 971 66 1005
rect 100 971 378 1005
rect 412 971 657 1005
rect 691 971 697 1005
rect 60 933 697 971
rect 60 899 66 933
rect 100 905 378 933
rect 100 899 106 905
rect 60 887 106 899
rect 372 899 378 905
rect 412 905 657 933
rect 412 899 418 905
rect 372 887 418 899
rect 651 899 657 905
rect 691 899 697 933
rect 651 887 697 899
rect 725 848 758 1025
tri 758 1000 783 1025 nw
tri 862 1019 868 1025 ne
rect 868 1019 998 1025
tri 1105 1000 1122 1017 se
rect 1122 1000 1824 1076
tri 1100 995 1105 1000 se
rect 1105 995 1824 1000
tri 1088 983 1100 995 se
rect 1100 983 1824 995
tri 1086 981 1088 983 se
rect 1088 981 1130 983
rect 786 975 916 981
rect 786 941 798 975
rect 832 941 870 975
rect 904 941 916 975
tri 1071 966 1086 981 se
rect 1086 966 1130 981
rect 786 935 916 941
tri 844 925 854 935 ne
rect 854 925 906 935
tri 906 925 916 935 nw
rect 952 949 1130 966
rect 1164 949 1442 983
rect 1476 949 1754 983
rect 1788 949 1824 983
tri 948 925 952 929 se
rect 952 925 1824 949
tri 854 911 868 925 ne
rect 868 911 906 925
tri 868 908 871 911 ne
tri 758 848 775 865 sw
rect 725 841 775 848
tri 775 841 782 848 sw
rect 725 829 842 841
tri 694 795 725 826 se
rect 725 795 802 829
rect 836 795 842 829
tri 682 783 694 795 se
rect 694 783 842 795
rect 172 771 842 783
rect 172 737 185 771
rect 219 737 257 771
rect 291 737 503 771
rect 537 737 575 771
rect 609 757 842 771
rect 609 737 802 757
rect 172 731 802 737
tri 755 723 763 731 ne
rect 763 723 802 731
rect 836 723 842 757
tri 763 711 775 723 ne
rect 775 711 842 723
tri 775 706 780 711 ne
rect 780 706 842 711
tri 780 691 795 706 ne
rect 111 661 223 667
rect 111 655 522 661
rect 111 621 123 655
rect 157 621 212 655
rect 246 621 300 655
rect 334 621 388 655
rect 422 621 476 655
rect 510 621 522 655
rect 111 615 522 621
rect 579 655 709 661
rect 579 621 591 655
rect 625 621 663 655
rect 697 621 709 655
rect 579 615 709 621
rect 56 555 643 561
rect 56 521 90 555
rect 124 521 165 555
rect 199 521 240 555
rect 274 521 314 555
rect 348 544 643 555
tri 643 544 660 561 sw
rect 348 538 660 544
tri 660 538 666 544 sw
tri 789 538 795 544 se
rect 795 538 842 706
rect 871 795 906 911
tri 937 914 948 925 se
rect 948 914 1824 925
rect 937 911 1824 914
rect 937 882 1130 911
rect 937 848 949 882
rect 983 848 1021 882
rect 1055 877 1130 882
rect 1164 877 1442 911
rect 1476 877 1754 911
rect 1788 877 1824 911
rect 1055 865 1824 877
rect 1055 848 1067 865
rect 937 842 1067 848
tri 1067 842 1090 865 nw
tri 906 795 933 822 sw
rect 871 783 1842 795
rect 871 749 1286 783
rect 1320 749 1598 783
rect 1632 749 1842 783
rect 871 711 1842 749
rect 871 706 1286 711
rect 871 672 883 706
rect 917 672 955 706
rect 989 677 1286 706
rect 1320 677 1598 711
rect 1632 677 1842 711
rect 989 672 1842 677
rect 871 666 1842 672
rect 1280 665 1326 666
rect 1592 665 1713 666
tri 1713 665 1714 666 nw
tri 1605 661 1609 665 ne
rect 1609 661 1683 665
tri 1609 633 1637 661 ne
rect 1175 616 1587 622
rect 1175 582 1187 616
rect 1221 582 1276 616
rect 1310 582 1365 616
rect 1399 582 1453 616
rect 1487 582 1541 616
rect 1575 582 1587 616
rect 1175 576 1587 582
tri 1631 538 1637 544 se
rect 1637 538 1683 661
tri 1683 635 1713 665 nw
rect 348 521 666 538
rect 56 515 666 521
tri 623 510 628 515 ne
rect 628 510 666 515
tri 666 510 694 538 sw
tri 761 510 789 538 se
rect 789 510 842 538
tri 1605 512 1631 538 se
rect 1631 512 1683 538
tri 628 504 634 510 ne
rect 634 504 842 510
tri 634 495 643 504 ne
rect 643 495 686 504
tri 643 482 656 495 ne
rect 656 482 686 495
rect 56 476 614 482
rect 56 442 372 476
rect 406 442 444 476
rect 478 473 614 476
tri 614 473 623 482 sw
tri 656 473 665 482 ne
rect 665 473 686 482
rect 478 470 623 473
tri 623 470 626 473 sw
tri 665 470 668 473 ne
rect 668 470 686 473
rect 720 470 758 504
rect 792 470 842 504
rect 478 464 626 470
tri 626 464 632 470 sw
tri 668 464 674 470 ne
rect 674 464 842 470
rect 1036 504 1683 512
rect 1036 470 1048 504
rect 1082 470 1121 504
rect 1155 470 1193 504
rect 1227 470 1413 504
rect 1447 470 1488 504
rect 1522 470 1563 504
rect 1597 470 1637 504
rect 1671 470 1683 504
rect 1036 466 1683 470
rect 1036 464 1239 466
rect 1401 464 1683 466
rect 1727 610 1773 622
rect 1727 576 1733 610
rect 1767 576 1773 610
rect 1727 538 1773 576
rect 1727 504 1733 538
rect 1767 504 1773 538
rect 478 442 632 464
rect 56 436 632 442
tri 594 431 599 436 ne
rect 599 431 632 436
tri 632 431 665 464 sw
tri 1710 431 1727 448 se
rect 1727 431 1773 504
tri 599 425 605 431 ne
rect 605 428 1773 431
rect 605 425 1730 428
tri 605 416 614 425 ne
rect 614 416 874 425
tri 614 405 625 416 ne
rect 625 405 874 416
rect 56 399 565 405
rect 56 365 90 399
rect 124 365 165 399
rect 199 365 240 399
rect 274 365 314 399
rect 348 391 565 399
tri 565 391 579 405 sw
tri 625 391 639 405 ne
rect 639 391 874 405
rect 908 391 946 425
rect 980 391 1268 425
rect 1302 391 1340 425
rect 1374 391 1730 425
rect 348 385 579 391
tri 579 385 585 391 sw
tri 639 385 645 391 ne
rect 645 385 1730 391
tri 1730 385 1773 428 nw
rect 348 365 585 385
rect 56 359 585 365
tri 545 354 550 359 ne
rect 550 354 585 359
tri 585 354 616 385 sw
tri 550 348 556 354 ne
rect 556 348 824 354
tri 556 339 565 348 ne
rect 565 339 689 348
tri 565 314 590 339 ne
rect 590 314 689 339
rect 723 314 761 348
rect 795 314 824 348
tri 590 308 596 314 ne
rect 596 308 824 314
rect 956 348 1687 355
rect 956 314 969 348
rect 1003 314 1044 348
rect 1078 314 1119 348
rect 1153 314 1193 348
rect 1227 314 1413 348
rect 1447 314 1488 348
rect 1522 314 1563 348
rect 1597 314 1637 348
rect 1671 314 1687 348
rect 956 309 1687 314
rect 957 308 1294 309
tri 1294 308 1295 309 nw
rect 1401 308 1683 309
tri 643 307 644 308 ne
rect 644 307 824 308
rect 187 301 317 307
rect 187 267 199 301
rect 233 267 271 301
rect 305 267 317 301
tri 644 295 656 307 ne
rect 656 295 824 307
rect 187 261 317 267
rect 368 289 498 295
rect 368 255 380 289
rect 414 255 452 289
rect 486 255 498 289
tri 656 287 664 295 ne
rect 664 287 824 295
tri 1198 287 1219 308 ne
rect 1219 287 1266 308
tri 664 274 677 287 ne
rect 677 280 824 287
tri 824 280 831 287 sw
tri 1219 280 1226 287 ne
rect 368 249 498 255
rect 677 260 831 280
tri 831 260 851 280 sw
rect 677 254 1190 260
rect 677 220 690 254
rect 724 220 762 254
rect 796 220 1072 254
rect 1106 220 1144 254
rect 1178 220 1190 254
rect 677 214 1190 220
rect 231 182 277 186
rect 1226 182 1266 287
tri 1266 280 1294 308 nw
rect 1295 243 1724 249
rect 1295 209 1307 243
rect 1341 209 1382 243
rect 1416 209 1456 243
rect 1490 209 1530 243
rect 1564 209 1604 243
rect 1638 209 1678 243
rect 1712 209 1724 243
rect 1295 203 1724 209
tri 1266 182 1276 192 sw
rect 231 174 1028 182
rect 231 140 237 174
rect 271 167 1028 174
tri 1028 167 1043 182 sw
rect 1226 173 1276 182
tri 1276 173 1285 182 sw
rect 1226 167 1801 173
rect 271 150 1043 167
rect 271 140 277 150
rect 231 102 277 140
tri 1014 137 1027 150 ne
rect 1027 137 1043 150
tri 1043 137 1073 167 sw
tri 1027 136 1028 137 ne
rect 1028 136 1073 137
tri 1028 133 1031 136 ne
rect 1031 133 1073 136
tri 1073 133 1077 137 sw
rect 1226 133 1273 167
rect 1307 133 1345 167
rect 1379 139 1683 167
rect 1379 133 1419 139
tri 1419 133 1425 139 nw
tri 1615 133 1621 139 ne
rect 1621 133 1683 139
rect 1717 133 1755 167
rect 1789 133 1801 167
tri 1031 107 1057 133 ne
rect 1057 110 1077 133
tri 1077 110 1100 133 sw
rect 1226 127 1413 133
tri 1413 127 1419 133 nw
tri 1621 127 1627 133 ne
rect 1627 127 1801 133
rect 1057 107 1100 110
rect 231 68 237 102
rect 271 68 277 102
tri 136 48 145 57 se
rect 145 48 191 57
rect 231 56 277 68
rect 483 55 489 107
rect 541 55 553 107
rect 605 104 611 107
tri 1057 104 1060 107 ne
rect 1060 104 1100 107
tri 1100 104 1106 110 sw
tri 1445 104 1451 110 se
rect 1451 104 1581 110
rect 605 58 613 104
tri 1060 91 1073 104 ne
rect 1073 91 1106 104
tri 1106 91 1119 104 sw
tri 1432 91 1445 104 se
rect 1445 91 1463 104
tri 1073 70 1094 91 ne
rect 1094 70 1463 91
rect 1497 70 1535 104
rect 1569 70 1581 104
tri 1094 59 1105 70 ne
rect 1105 64 1581 70
rect 1105 59 1456 64
tri 1456 59 1461 64 nw
rect 605 55 611 58
tri 133 45 136 48 se
rect 136 47 191 48
tri 191 47 192 48 sw
rect 136 45 192 47
tri 124 36 133 45 se
rect 133 36 151 45
rect 68 11 151 36
rect 185 43 192 45
tri 192 43 196 47 sw
tri 313 43 317 47 se
rect 317 43 363 47
rect 185 35 196 43
tri 196 35 204 43 sw
tri 305 35 313 43 se
rect 313 35 363 43
rect 185 26 204 35
tri 204 26 213 35 sw
tri 296 26 305 35 se
rect 305 26 323 35
rect 185 11 323 26
rect 68 1 323 11
rect 357 1 363 35
rect 68 -27 363 1
rect 68 -61 151 -27
rect 185 -37 363 -27
rect 185 -61 323 -37
rect 68 -71 323 -61
rect 357 -71 363 -37
rect 68 -83 363 -71
rect 403 43 449 55
rect 403 9 409 43
rect 443 11 449 43
tri 759 36 762 39 se
rect 762 36 1015 39
tri 756 33 759 36 se
rect 759 33 1015 36
tri 734 11 756 33 se
rect 756 11 897 33
rect 443 9 897 11
rect 403 -1 897 9
rect 931 -1 969 33
rect 1003 -1 1015 33
rect 403 -7 1015 -1
rect 403 -29 754 -7
rect 403 -63 409 -29
rect 443 -35 754 -29
tri 754 -35 782 -7 nw
rect 443 -63 449 -35
rect 403 -75 449 -63
<< via1 >>
rect 489 98 541 107
rect 489 64 495 98
rect 495 64 529 98
rect 529 64 541 98
rect 489 55 541 64
rect 553 98 605 107
rect 553 64 567 98
rect 567 64 601 98
rect 601 64 605 98
rect 553 55 605 64
<< metal2 >>
rect 483 55 489 107
rect 541 55 553 107
rect 605 55 611 107
use sky130_fd_pr__nfet_01v8__example_55959141808498  sky130_fd_pr__nfet_01v8__example_55959141808498_0
timestamp 1619729480
transform -1 0 484 0 1 13
box -28 0 144 97
use sky130_fd_pr__nfet_01v8__example_55959141808498  sky130_fd_pr__nfet_01v8__example_55959141808498_1
timestamp 1619729480
transform -1 0 312 0 1 13
box -28 0 144 97
use sky130_fd_pr__nfet_01v8__example_55959141808497  sky130_fd_pr__nfet_01v8__example_55959141808497_0
timestamp 1619729480
transform -1 0 1151 0 1 -33
box -28 0 444 97
use sky130_fd_pr__nfet_01v8__example_55959141808496  sky130_fd_pr__nfet_01v8__example_55959141808496_0
timestamp 1619729480
transform -1 0 1744 0 -1 167
box -28 0 444 97
use sky130_fd_pr__nfet_01v8__example_55959141808495  sky130_fd_pr__nfet_01v8__example_55959141808495_0
timestamp 1619729480
transform 0 1 526 -1 0 459
box -28 0 128 131
use sky130_fd_pr__nfet_01v8__example_55959141808495  sky130_fd_pr__nfet_01v8__example_55959141808495_1
timestamp 1619729480
transform 0 1 956 -1 0 459
box -28 0 128 131
use sky130_fd_pr__nfet_01v8__example_55959141808495  sky130_fd_pr__nfet_01v8__example_55959141808495_2
timestamp 1619729480
transform 0 1 1386 -1 0 459
box -28 0 128 131
use sky130_fd_pr__nfet_01v8__example_55959141808495  sky130_fd_pr__nfet_01v8__example_55959141808495_3
timestamp 1619729480
transform 0 1 96 -1 0 510
box -28 0 128 131
use sky130_fd_pr__nfet_01v8__example_55959141808494  sky130_fd_pr__nfet_01v8__example_55959141808494_0
timestamp 1619729480
transform -1 0 679 0 -1 1003
box -28 0 128 131
use sky130_fd_pr__nfet_01v8__example_55959141808493  sky130_fd_pr__nfet_01v8__example_55959141808493_0
timestamp 1619729480
transform -1 0 523 0 -1 1003
box -28 0 440 131
use sky130_fd_pr__pfet_01v8__example_55959141808492  sky130_fd_pr__pfet_01v8__example_55959141808492_0
timestamp 1619729480
transform 0 1 884 -1 0 837
box -28 0 148 63
use sky130_fd_pr__pfet_01v8__example_55959141808492  sky130_fd_pr__pfet_01v8__example_55959141808492_1
timestamp 1619729480
transform 0 1 884 1 0 893
box -28 0 148 63
use sky130_fd_pr__pfet_01v8__example_55959141808490  sky130_fd_pr__pfet_01v8__example_55959141808490_0
timestamp 1619729480
transform 1 0 1175 0 -1 964
box -28 0 440 131
use sky130_fd_pr__pfet_01v8__example_55959141808489  sky130_fd_pr__pfet_01v8__example_55959141808489_0
timestamp 1619729480
transform 1 0 1643 0 -1 964
box -28 0 128 131
<< labels >>
flabel metal1 s 726 733 754 773 3 FreeSans 280 180 0 0 OUT_H
flabel metal1 s 1309 587 1337 615 3 FreeSans 280 0 0 0 RST2_H_N
flabel metal1 s 73 961 101 989 3 FreeSans 280 0 0 0 VGND
flabel metal1 s 1800 666 1828 795 3 FreeSans 280 180 0 0 OUT_H_N
flabel metal1 s 1626 212 1654 240 3 FreeSans 280 0 0 0 VPWR_LV
flabel metal1 s 159 447 187 475 3 FreeSans 280 0 0 0 RST_H_N
flabel metal1 s 232 266 260 294 3 FreeSans 280 0 0 0 IN
flabel metal1 s 411 -18 439 10 3 FreeSans 280 0 0 0 IN_B
flabel metal1 s 73 -17 101 11 3 FreeSans 280 0 0 0 VGND
flabel metal1 s 1505 998 1505 998 3 FreeSans 280 0 0 0 VPWR_HV
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 48487398
string GDS_START 48462034
<< end >>
