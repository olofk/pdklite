magic
tech sky130A
magscale 1 2
timestamp 1640697850
use sky130_fd_pr__hvdfl1sd__example_5595914180851  sky130_fd_pr__hvdfl1sd__example_5595914180851_0
timestamp 1640697850
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_5595914180851  sky130_fd_pr__hvdfl1sd__example_5595914180851_1
timestamp 1640697850
transform 1 0 1600 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 1628 471 1628 471 0 FreeSans 300 0 0 0 D
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 11344032
string GDS_START 11342978
<< end >>
