magic
tech sky130A
magscale 1 2
timestamp 1640697980
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 21 1887 203
rect 30 -17 64 21
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 119 359 161 527
rect 279 427 329 527
rect 447 427 497 527
rect 615 427 665 527
rect 783 323 833 425
rect 949 323 993 425
rect 277 289 715 323
rect 277 257 311 289
rect 20 215 311 257
rect 345 215 615 255
rect 649 215 715 289
rect 749 283 993 323
rect 1231 359 1273 527
rect 1391 359 1441 527
rect 749 181 783 283
rect 1189 215 1464 255
rect 1519 215 1809 255
rect 35 17 69 179
rect 203 17 237 111
rect 355 145 1009 181
rect 355 129 599 145
rect 707 17 741 111
rect 775 55 841 145
rect 875 17 909 111
rect 943 55 1009 145
rect 1043 17 1181 111
rect 1315 17 1349 111
rect 1483 17 1517 111
rect 1651 17 1685 111
rect 1819 17 1853 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< obsli1 >>
rect 17 325 85 493
rect 195 393 243 493
rect 363 393 413 493
rect 531 393 581 493
rect 699 459 1093 493
rect 699 393 749 459
rect 195 359 749 393
rect 195 325 243 359
rect 17 291 243 325
rect 867 359 915 459
rect 1027 291 1093 459
rect 1131 325 1197 493
rect 1308 325 1356 493
rect 1475 459 1862 493
rect 1475 325 1525 459
rect 1131 291 1525 325
rect 1559 325 1609 425
rect 1643 359 1693 459
rect 1727 325 1777 425
rect 1812 359 1862 459
rect 1559 291 1915 325
rect 817 215 1145 249
rect 1111 181 1145 215
rect 1843 181 1915 291
rect 103 145 321 181
rect 103 51 169 145
rect 271 95 321 145
rect 1111 147 1915 181
rect 271 51 673 95
rect 1215 145 1785 147
rect 1215 51 1281 145
rect 1383 51 1449 145
rect 1551 51 1617 145
rect 1719 51 1785 145
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
rlabel locali s 1189 215 1464 255 6 A1_N
port 1 nsew signal input
rlabel locali s 1519 215 1809 255 6 A2_N
port 2 nsew signal input
rlabel locali s 649 215 715 289 6 B1
port 3 nsew signal input
rlabel locali s 20 215 311 257 6 B1
port 3 nsew signal input
rlabel locali s 277 257 311 289 6 B1
port 3 nsew signal input
rlabel locali s 277 289 715 323 6 B1
port 3 nsew signal input
rlabel locali s 345 215 615 255 6 B2
port 4 nsew signal input
rlabel metal1 s 0 -48 1932 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1869 -17 1903 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1777 -17 1811 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1685 -17 1719 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1593 -17 1627 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1501 -17 1535 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1409 -17 1443 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1317 -17 1351 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1225 -17 1259 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1133 -17 1167 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1041 -17 1075 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 949 -17 983 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 857 -17 891 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 765 -17 799 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 673 -17 707 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 581 -17 615 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 489 -17 523 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 397 -17 431 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 305 -17 339 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 213 -17 247 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 121 -17 155 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 29 -17 63 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1932 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1819 17 1853 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1651 17 1685 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1483 17 1517 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1315 17 1349 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1043 17 1181 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 875 17 909 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 707 17 741 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 203 17 237 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 35 17 69 179 6 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 1887 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1970 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1869 527 1903 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1777 527 1811 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1685 527 1719 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1593 527 1627 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1501 527 1535 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1409 527 1443 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1317 527 1351 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1225 527 1259 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1133 527 1167 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1041 527 1075 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 949 527 983 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 857 527 891 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 765 527 799 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 673 527 707 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 581 527 615 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 489 527 523 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 397 527 431 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 305 527 339 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 213 527 247 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 121 527 155 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 29 527 63 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1391 359 1441 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1231 359 1273 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 615 427 665 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 447 427 497 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 279 427 329 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 119 359 161 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1932 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 943 55 1009 145 6 Y
port 9 nsew signal output
rlabel locali s 775 55 841 145 6 Y
port 9 nsew signal output
rlabel locali s 355 129 599 145 6 Y
port 9 nsew signal output
rlabel locali s 355 145 1009 181 6 Y
port 9 nsew signal output
rlabel locali s 749 181 783 283 6 Y
port 9 nsew signal output
rlabel locali s 749 283 993 323 6 Y
port 9 nsew signal output
rlabel locali s 949 323 993 425 6 Y
port 9 nsew signal output
rlabel locali s 783 323 833 425 6 Y
port 9 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3972394
string GDS_START 3958152
<< end >>
