magic
tech sky130A
magscale 1 2
timestamp 1640697980
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 7 21 1463 203
rect 29 -17 63 21
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 33 289 83 527
rect 201 425 251 527
rect 713 425 757 527
rect 885 425 933 527
rect 369 391 419 425
rect 537 391 587 425
rect 1387 425 1443 527
rect 369 357 783 391
rect 1051 391 1101 425
rect 1219 391 1269 425
rect 1051 357 1455 391
rect 749 323 783 357
rect 230 289 715 323
rect 749 289 825 323
rect 230 255 283 289
rect 17 215 283 255
rect 337 215 619 255
rect 655 249 715 289
rect 655 215 721 249
rect 125 17 159 111
rect 293 17 327 111
rect 461 17 495 111
rect 629 17 663 111
rect 791 164 825 289
rect 859 289 1387 323
rect 859 199 988 289
rect 1022 215 1292 255
rect 1343 199 1387 289
rect 1421 164 1455 357
rect 791 129 1455 164
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< obsli1 >>
rect 117 391 167 493
rect 285 459 679 493
rect 285 391 335 459
rect 453 425 503 459
rect 621 425 679 459
rect 791 425 851 493
rect 967 459 1353 493
rect 117 357 335 391
rect 817 391 851 425
rect 967 391 1017 459
rect 1135 425 1185 459
rect 1303 427 1353 459
rect 817 357 1017 391
rect 117 289 167 357
rect 25 147 757 181
rect 25 145 259 147
rect 25 51 91 145
rect 193 51 259 145
rect 361 145 595 147
rect 361 51 427 145
rect 529 51 595 145
rect 697 95 757 147
rect 697 51 1449 95
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
rlabel locali s 655 215 721 249 6 A1
port 1 nsew signal input
rlabel locali s 655 249 715 289 6 A1
port 1 nsew signal input
rlabel locali s 17 215 283 255 6 A1
port 1 nsew signal input
rlabel locali s 230 255 283 289 6 A1
port 1 nsew signal input
rlabel locali s 230 289 715 323 6 A1
port 1 nsew signal input
rlabel locali s 337 215 619 255 6 A2
port 2 nsew signal input
rlabel locali s 1343 199 1387 289 6 B1
port 3 nsew signal input
rlabel locali s 859 199 988 289 6 B1
port 3 nsew signal input
rlabel locali s 859 289 1387 323 6 B1
port 3 nsew signal input
rlabel locali s 1022 215 1292 255 6 B2
port 4 nsew signal input
rlabel metal1 s 0 -48 1472 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1409 -17 1443 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1317 -17 1351 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1225 -17 1259 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1133 -17 1167 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1041 -17 1075 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 949 -17 983 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 857 -17 891 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 765 -17 799 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 673 -17 707 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 581 -17 615 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 489 -17 523 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 397 -17 431 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 305 -17 339 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 213 -17 247 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 121 -17 155 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 29 -17 63 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1472 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 629 17 663 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 461 17 495 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 293 17 327 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 125 17 159 111 6 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 7 21 1463 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1510 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1472 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1409 527 1443 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1317 527 1351 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1225 527 1259 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1133 527 1167 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1041 527 1075 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 949 527 983 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 857 527 891 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 765 527 799 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 673 527 707 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 581 527 615 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 489 527 523 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 397 527 431 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 305 527 339 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 213 527 247 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 121 527 155 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 29 527 63 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1387 425 1443 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 885 425 933 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 713 425 757 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 201 425 251 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 33 289 83 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1472 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 791 129 1455 164 6 Y
port 9 nsew signal output
rlabel locali s 1421 164 1455 357 6 Y
port 9 nsew signal output
rlabel locali s 791 164 825 289 6 Y
port 9 nsew signal output
rlabel locali s 749 289 825 323 6 Y
port 9 nsew signal output
rlabel locali s 749 323 783 357 6 Y
port 9 nsew signal output
rlabel locali s 1051 357 1455 391 6 Y
port 9 nsew signal output
rlabel locali s 369 357 783 391 6 Y
port 9 nsew signal output
rlabel locali s 1219 391 1269 425 6 Y
port 9 nsew signal output
rlabel locali s 1051 391 1101 425 6 Y
port 9 nsew signal output
rlabel locali s 537 391 587 425 6 Y
port 9 nsew signal output
rlabel locali s 369 391 419 425 6 Y
port 9 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1417224
string GDS_START 1406620
<< end >>
