magic
tech sky130A
magscale 1 2
timestamp 1640697980
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 1 21 2203 203
rect 30 -17 64 21
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 119 357 153 527
rect 287 357 321 527
rect 455 367 489 527
rect 623 367 657 527
rect 791 367 825 527
rect 859 323 925 493
rect 959 367 993 527
rect 1027 323 1093 493
rect 1127 367 1161 527
rect 1195 323 1261 493
rect 1295 367 1329 527
rect 1363 323 1429 493
rect 1463 367 1497 527
rect 1531 323 1597 493
rect 1631 367 1665 527
rect 1699 323 1765 493
rect 1799 367 1833 527
rect 1867 323 1933 493
rect 1967 367 2001 527
rect 2035 323 2101 493
rect 2135 367 2169 527
rect 859 289 2191 323
rect 18 215 253 255
rect 2136 181 2191 289
rect 859 147 2191 181
rect 119 17 153 113
rect 287 17 321 113
rect 455 17 489 113
rect 623 17 657 113
rect 791 17 825 113
rect 859 52 925 147
rect 859 51 909 52
rect 959 17 993 113
rect 1027 52 1093 147
rect 1043 51 1077 52
rect 1127 17 1161 113
rect 1195 52 1261 147
rect 1211 51 1245 52
rect 1295 17 1329 113
rect 1363 52 1429 147
rect 1463 17 1497 113
rect 1531 52 1597 147
rect 1631 17 1665 113
rect 1699 52 1765 147
rect 1799 17 1833 113
rect 1867 52 1933 147
rect 1967 17 2001 113
rect 2035 52 2101 147
rect 2135 17 2169 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< obsli1 >>
rect 19 323 85 493
rect 187 323 253 493
rect 355 323 421 493
rect 523 323 589 493
rect 691 323 757 493
rect 19 289 321 323
rect 355 289 825 323
rect 287 255 321 289
rect 790 255 825 289
rect 287 215 749 255
rect 790 215 2102 255
rect 287 181 321 215
rect 790 181 825 215
rect 19 147 321 181
rect 355 147 825 181
rect 19 52 85 147
rect 187 52 253 147
rect 355 52 421 147
rect 523 52 589 147
rect 691 52 757 147
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
rlabel locali s 18 215 253 255 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 2208 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 2145 -17 2179 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 2053 -17 2087 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 1961 -17 1995 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 1869 -17 1903 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 1777 -17 1811 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 1685 -17 1719 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 1593 -17 1627 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 1501 -17 1535 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 1409 -17 1443 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 1317 -17 1351 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 1225 -17 1259 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 1133 -17 1167 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 1041 -17 1075 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 949 -17 983 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 857 -17 891 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 765 -17 799 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 673 -17 707 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 581 -17 615 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 489 -17 523 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 397 -17 431 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 305 -17 339 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 213 -17 247 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 121 -17 155 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel viali s 29 -17 63 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 0 -17 2208 17 8 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 2135 17 2169 113 6 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 1967 17 2001 113 6 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 1799 17 1833 113 6 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 1631 17 1665 113 6 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 1463 17 1497 113 6 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 1295 17 1329 113 6 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 1127 17 1161 113 6 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 959 17 993 113 6 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 791 17 825 113 6 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 623 17 657 113 6 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 455 17 489 113 6 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 287 17 321 113 6 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 119 17 153 113 6 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 2203 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 2246 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 2208 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 2145 527 2179 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 2053 527 2087 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1961 527 1995 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1869 527 1903 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1777 527 1811 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1685 527 1719 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1593 527 1627 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1501 527 1535 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1409 527 1443 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1317 527 1351 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1225 527 1259 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1133 527 1167 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1041 527 1075 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 949 527 983 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 857 527 891 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 765 527 799 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 673 527 707 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 581 527 615 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 489 527 523 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 397 527 431 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 305 527 339 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 213 527 247 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 121 527 155 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 29 527 63 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 2135 367 2169 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1967 367 2001 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1799 367 1833 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1631 367 1665 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1463 367 1497 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1295 367 1329 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1127 367 1161 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 959 367 993 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 791 367 825 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 623 367 657 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 455 367 489 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 287 357 321 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 119 357 153 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 2208 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1211 51 1245 52 6 Y
port 6 nsew signal output
rlabel locali s 1043 51 1077 52 6 Y
port 6 nsew signal output
rlabel locali s 859 51 909 52 6 Y
port 6 nsew signal output
rlabel locali s 2035 52 2101 147 6 Y
port 6 nsew signal output
rlabel locali s 1867 52 1933 147 6 Y
port 6 nsew signal output
rlabel locali s 1699 52 1765 147 6 Y
port 6 nsew signal output
rlabel locali s 1531 52 1597 147 6 Y
port 6 nsew signal output
rlabel locali s 1363 52 1429 147 6 Y
port 6 nsew signal output
rlabel locali s 1195 52 1261 147 6 Y
port 6 nsew signal output
rlabel locali s 1027 52 1093 147 6 Y
port 6 nsew signal output
rlabel locali s 859 52 925 147 6 Y
port 6 nsew signal output
rlabel locali s 859 147 2191 181 6 Y
port 6 nsew signal output
rlabel locali s 2136 181 2191 289 6 Y
port 6 nsew signal output
rlabel locali s 859 289 2191 323 6 Y
port 6 nsew signal output
rlabel locali s 2035 323 2101 493 6 Y
port 6 nsew signal output
rlabel locali s 1867 323 1933 493 6 Y
port 6 nsew signal output
rlabel locali s 1699 323 1765 493 6 Y
port 6 nsew signal output
rlabel locali s 1531 323 1597 493 6 Y
port 6 nsew signal output
rlabel locali s 1363 323 1429 493 6 Y
port 6 nsew signal output
rlabel locali s 1195 323 1261 493 6 Y
port 6 nsew signal output
rlabel locali s 1027 323 1093 493 6 Y
port 6 nsew signal output
rlabel locali s 859 323 925 493 6 Y
port 6 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2208 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3223662
string GDS_START 3206836
<< end >>
