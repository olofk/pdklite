magic
tech sky130A
magscale 1 2
timestamp 1619729575
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 29 -17 63 17
<< locali >>
rect 100 202 166 325
rect 200 319 482 353
rect 200 157 247 319
rect 849 319 1078 353
rect 849 255 884 319
rect 805 202 884 255
rect 918 202 991 272
rect 1044 258 1078 319
rect 1044 211 1140 258
rect 200 123 468 157
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 21 421 110 493
rect 144 455 210 527
rect 316 455 382 527
rect 487 455 554 527
rect 611 442 813 476
rect 847 455 913 527
rect 1015 455 1081 527
rect 21 387 574 421
rect 21 359 113 387
rect 21 168 66 359
rect 21 51 108 168
rect 540 305 574 387
rect 611 339 645 442
rect 777 421 813 442
rect 777 387 1165 421
rect 540 271 661 305
rect 281 237 506 265
rect 281 199 562 237
rect 599 199 661 271
rect 528 160 562 199
rect 695 168 729 361
rect 777 289 813 387
rect 1114 292 1165 387
rect 528 157 602 160
rect 695 157 993 168
rect 528 134 993 157
rect 528 123 729 134
rect 142 17 210 89
rect 316 17 382 89
rect 503 17 657 89
rect 695 51 729 123
rect 771 17 837 89
rect 937 81 993 134
rect 1109 17 1165 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 918 202 991 272 6 A1
port 1 nsew signal input
rlabel locali s 1044 258 1078 319 6 A2
port 2 nsew signal input
rlabel locali s 1044 211 1140 258 6 A2
port 2 nsew signal input
rlabel locali s 849 319 1078 353 6 A2
port 2 nsew signal input
rlabel locali s 849 255 884 319 6 A2
port 2 nsew signal input
rlabel locali s 805 202 884 255 6 A2
port 2 nsew signal input
rlabel locali s 100 202 166 325 6 B1_N
port 3 nsew signal input
rlabel locali s 200 319 482 353 6 X
port 8 nsew signal output
rlabel locali s 200 157 247 319 6 X
port 8 nsew signal output
rlabel locali s 200 123 468 157 6 X
port 8 nsew signal output
rlabel metal1 s 0 -48 1196 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1234 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2637762
string GDS_START 2629514
<< end >>
