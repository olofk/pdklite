magic
tech sky130A
magscale 1 2
timestamp 1640697850
<< metal3 >>
rect 120 2304 4900 2306
rect 120 2240 126 2304
rect 190 2240 208 2304
rect 272 2240 290 2304
rect 354 2240 372 2304
rect 436 2240 454 2304
rect 518 2240 536 2304
rect 600 2240 618 2304
rect 682 2240 699 2304
rect 763 2240 780 2304
rect 844 2240 861 2304
rect 925 2240 942 2304
rect 1006 2240 1023 2304
rect 1087 2240 1104 2304
rect 1168 2240 1185 2304
rect 1249 2240 1266 2304
rect 1330 2240 1347 2304
rect 1411 2240 1428 2304
rect 1492 2240 1509 2304
rect 1573 2240 1590 2304
rect 1654 2240 1671 2304
rect 1735 2240 1752 2304
rect 1816 2240 1833 2304
rect 1897 2240 1914 2304
rect 1978 2240 1995 2304
rect 2059 2240 2076 2304
rect 2140 2240 2157 2304
rect 2221 2240 2238 2304
rect 2302 2240 2319 2304
rect 2383 2240 2400 2304
rect 2464 2240 2481 2304
rect 2545 2240 2562 2304
rect 2626 2240 2643 2304
rect 2707 2240 2724 2304
rect 2788 2240 2805 2304
rect 2869 2240 2886 2304
rect 2950 2240 2967 2304
rect 3031 2240 3048 2304
rect 3112 2240 3129 2304
rect 3193 2240 3210 2304
rect 3274 2240 3291 2304
rect 3355 2240 3372 2304
rect 3436 2240 3453 2304
rect 3517 2240 3534 2304
rect 3598 2240 3615 2304
rect 3679 2240 3696 2304
rect 3760 2240 3777 2304
rect 3841 2240 3858 2304
rect 3922 2240 3939 2304
rect 4003 2240 4020 2304
rect 4084 2240 4101 2304
rect 4165 2240 4182 2304
rect 4246 2240 4263 2304
rect 4327 2240 4344 2304
rect 4408 2240 4425 2304
rect 4489 2240 4506 2304
rect 4570 2240 4587 2304
rect 4651 2240 4668 2304
rect 4732 2240 4749 2304
rect 4813 2240 4830 2304
rect 4894 2240 4900 2304
rect 120 2218 4900 2240
rect 120 2154 126 2218
rect 190 2154 208 2218
rect 272 2154 290 2218
rect 354 2154 372 2218
rect 436 2154 454 2218
rect 518 2154 536 2218
rect 600 2154 618 2218
rect 682 2154 699 2218
rect 763 2154 780 2218
rect 844 2154 861 2218
rect 925 2154 942 2218
rect 1006 2154 1023 2218
rect 1087 2154 1104 2218
rect 1168 2154 1185 2218
rect 1249 2154 1266 2218
rect 1330 2154 1347 2218
rect 1411 2154 1428 2218
rect 1492 2154 1509 2218
rect 1573 2154 1590 2218
rect 1654 2154 1671 2218
rect 1735 2154 1752 2218
rect 1816 2154 1833 2218
rect 1897 2154 1914 2218
rect 1978 2154 1995 2218
rect 2059 2154 2076 2218
rect 2140 2154 2157 2218
rect 2221 2154 2238 2218
rect 2302 2154 2319 2218
rect 2383 2154 2400 2218
rect 2464 2154 2481 2218
rect 2545 2154 2562 2218
rect 2626 2154 2643 2218
rect 2707 2154 2724 2218
rect 2788 2154 2805 2218
rect 2869 2154 2886 2218
rect 2950 2154 2967 2218
rect 3031 2154 3048 2218
rect 3112 2154 3129 2218
rect 3193 2154 3210 2218
rect 3274 2154 3291 2218
rect 3355 2154 3372 2218
rect 3436 2154 3453 2218
rect 3517 2154 3534 2218
rect 3598 2154 3615 2218
rect 3679 2154 3696 2218
rect 3760 2154 3777 2218
rect 3841 2154 3858 2218
rect 3922 2154 3939 2218
rect 4003 2154 4020 2218
rect 4084 2154 4101 2218
rect 4165 2154 4182 2218
rect 4246 2154 4263 2218
rect 4327 2154 4344 2218
rect 4408 2154 4425 2218
rect 4489 2154 4506 2218
rect 4570 2154 4587 2218
rect 4651 2154 4668 2218
rect 4732 2154 4749 2218
rect 4813 2154 4830 2218
rect 4894 2154 4900 2218
rect 120 2132 4900 2154
rect 120 2068 126 2132
rect 190 2068 208 2132
rect 272 2068 290 2132
rect 354 2068 372 2132
rect 436 2068 454 2132
rect 518 2068 536 2132
rect 600 2068 618 2132
rect 682 2068 699 2132
rect 763 2068 780 2132
rect 844 2068 861 2132
rect 925 2068 942 2132
rect 1006 2068 1023 2132
rect 1087 2068 1104 2132
rect 1168 2068 1185 2132
rect 1249 2068 1266 2132
rect 1330 2068 1347 2132
rect 1411 2068 1428 2132
rect 1492 2068 1509 2132
rect 1573 2068 1590 2132
rect 1654 2068 1671 2132
rect 1735 2068 1752 2132
rect 1816 2068 1833 2132
rect 1897 2068 1914 2132
rect 1978 2068 1995 2132
rect 2059 2068 2076 2132
rect 2140 2068 2157 2132
rect 2221 2068 2238 2132
rect 2302 2068 2319 2132
rect 2383 2068 2400 2132
rect 2464 2068 2481 2132
rect 2545 2068 2562 2132
rect 2626 2068 2643 2132
rect 2707 2068 2724 2132
rect 2788 2068 2805 2132
rect 2869 2068 2886 2132
rect 2950 2068 2967 2132
rect 3031 2068 3048 2132
rect 3112 2068 3129 2132
rect 3193 2068 3210 2132
rect 3274 2068 3291 2132
rect 3355 2068 3372 2132
rect 3436 2068 3453 2132
rect 3517 2068 3534 2132
rect 3598 2068 3615 2132
rect 3679 2068 3696 2132
rect 3760 2068 3777 2132
rect 3841 2068 3858 2132
rect 3922 2068 3939 2132
rect 4003 2068 4020 2132
rect 4084 2068 4101 2132
rect 4165 2068 4182 2132
rect 4246 2068 4263 2132
rect 4327 2068 4344 2132
rect 4408 2068 4425 2132
rect 4489 2068 4506 2132
rect 4570 2068 4587 2132
rect 4651 2068 4668 2132
rect 4732 2068 4749 2132
rect 4813 2068 4830 2132
rect 4894 2068 4900 2132
rect 120 2046 4900 2068
rect 120 1982 126 2046
rect 190 1982 208 2046
rect 272 1982 290 2046
rect 354 1982 372 2046
rect 436 1982 454 2046
rect 518 1982 536 2046
rect 600 1982 618 2046
rect 682 1982 699 2046
rect 763 1982 780 2046
rect 844 1982 861 2046
rect 925 1982 942 2046
rect 1006 1982 1023 2046
rect 1087 1982 1104 2046
rect 1168 1982 1185 2046
rect 1249 1982 1266 2046
rect 1330 1982 1347 2046
rect 1411 1982 1428 2046
rect 1492 1982 1509 2046
rect 1573 1982 1590 2046
rect 1654 1982 1671 2046
rect 1735 1982 1752 2046
rect 1816 1982 1833 2046
rect 1897 1982 1914 2046
rect 1978 1982 1995 2046
rect 2059 1982 2076 2046
rect 2140 1982 2157 2046
rect 2221 1982 2238 2046
rect 2302 1982 2319 2046
rect 2383 1982 2400 2046
rect 2464 1982 2481 2046
rect 2545 1982 2562 2046
rect 2626 1982 2643 2046
rect 2707 1982 2724 2046
rect 2788 1982 2805 2046
rect 2869 1982 2886 2046
rect 2950 1982 2967 2046
rect 3031 1982 3048 2046
rect 3112 1982 3129 2046
rect 3193 1982 3210 2046
rect 3274 1982 3291 2046
rect 3355 1982 3372 2046
rect 3436 1982 3453 2046
rect 3517 1982 3534 2046
rect 3598 1982 3615 2046
rect 3679 1982 3696 2046
rect 3760 1982 3777 2046
rect 3841 1982 3858 2046
rect 3922 1982 3939 2046
rect 4003 1982 4020 2046
rect 4084 1982 4101 2046
rect 4165 1982 4182 2046
rect 4246 1982 4263 2046
rect 4327 1982 4344 2046
rect 4408 1982 4425 2046
rect 4489 1982 4506 2046
rect 4570 1982 4587 2046
rect 4651 1982 4668 2046
rect 4732 1982 4749 2046
rect 4813 1982 4830 2046
rect 4894 1982 4900 2046
rect 120 1960 4900 1982
rect 120 1896 126 1960
rect 190 1896 208 1960
rect 272 1896 290 1960
rect 354 1896 372 1960
rect 436 1896 454 1960
rect 518 1896 536 1960
rect 600 1896 618 1960
rect 682 1896 699 1960
rect 763 1896 780 1960
rect 844 1896 861 1960
rect 925 1896 942 1960
rect 1006 1896 1023 1960
rect 1087 1896 1104 1960
rect 1168 1896 1185 1960
rect 1249 1896 1266 1960
rect 1330 1896 1347 1960
rect 1411 1896 1428 1960
rect 1492 1896 1509 1960
rect 1573 1896 1590 1960
rect 1654 1896 1671 1960
rect 1735 1896 1752 1960
rect 1816 1896 1833 1960
rect 1897 1896 1914 1960
rect 1978 1896 1995 1960
rect 2059 1896 2076 1960
rect 2140 1896 2157 1960
rect 2221 1896 2238 1960
rect 2302 1896 2319 1960
rect 2383 1896 2400 1960
rect 2464 1896 2481 1960
rect 2545 1896 2562 1960
rect 2626 1896 2643 1960
rect 2707 1896 2724 1960
rect 2788 1896 2805 1960
rect 2869 1896 2886 1960
rect 2950 1896 2967 1960
rect 3031 1896 3048 1960
rect 3112 1896 3129 1960
rect 3193 1896 3210 1960
rect 3274 1896 3291 1960
rect 3355 1896 3372 1960
rect 3436 1896 3453 1960
rect 3517 1896 3534 1960
rect 3598 1896 3615 1960
rect 3679 1896 3696 1960
rect 3760 1896 3777 1960
rect 3841 1896 3858 1960
rect 3922 1896 3939 1960
rect 4003 1896 4020 1960
rect 4084 1896 4101 1960
rect 4165 1896 4182 1960
rect 4246 1896 4263 1960
rect 4327 1896 4344 1960
rect 4408 1896 4425 1960
rect 4489 1896 4506 1960
rect 4570 1896 4587 1960
rect 4651 1896 4668 1960
rect 4732 1896 4749 1960
rect 4813 1896 4830 1960
rect 4894 1896 4900 1960
rect 120 1874 4900 1896
rect 120 1810 126 1874
rect 190 1810 208 1874
rect 272 1810 290 1874
rect 354 1810 372 1874
rect 436 1810 454 1874
rect 518 1810 536 1874
rect 600 1810 618 1874
rect 682 1810 699 1874
rect 763 1810 780 1874
rect 844 1810 861 1874
rect 925 1810 942 1874
rect 1006 1810 1023 1874
rect 1087 1810 1104 1874
rect 1168 1810 1185 1874
rect 1249 1810 1266 1874
rect 1330 1810 1347 1874
rect 1411 1810 1428 1874
rect 1492 1810 1509 1874
rect 1573 1810 1590 1874
rect 1654 1810 1671 1874
rect 1735 1810 1752 1874
rect 1816 1810 1833 1874
rect 1897 1810 1914 1874
rect 1978 1810 1995 1874
rect 2059 1810 2076 1874
rect 2140 1810 2157 1874
rect 2221 1810 2238 1874
rect 2302 1810 2319 1874
rect 2383 1810 2400 1874
rect 2464 1810 2481 1874
rect 2545 1810 2562 1874
rect 2626 1810 2643 1874
rect 2707 1810 2724 1874
rect 2788 1810 2805 1874
rect 2869 1810 2886 1874
rect 2950 1810 2967 1874
rect 3031 1810 3048 1874
rect 3112 1810 3129 1874
rect 3193 1810 3210 1874
rect 3274 1810 3291 1874
rect 3355 1810 3372 1874
rect 3436 1810 3453 1874
rect 3517 1810 3534 1874
rect 3598 1810 3615 1874
rect 3679 1810 3696 1874
rect 3760 1810 3777 1874
rect 3841 1810 3858 1874
rect 3922 1810 3939 1874
rect 4003 1810 4020 1874
rect 4084 1810 4101 1874
rect 4165 1810 4182 1874
rect 4246 1810 4263 1874
rect 4327 1810 4344 1874
rect 4408 1810 4425 1874
rect 4489 1810 4506 1874
rect 4570 1810 4587 1874
rect 4651 1810 4668 1874
rect 4732 1810 4749 1874
rect 4813 1810 4830 1874
rect 4894 1810 4900 1874
rect 120 1788 4900 1810
rect 120 1724 126 1788
rect 190 1724 208 1788
rect 272 1724 290 1788
rect 354 1724 372 1788
rect 436 1724 454 1788
rect 518 1724 536 1788
rect 600 1724 618 1788
rect 682 1724 699 1788
rect 763 1724 780 1788
rect 844 1724 861 1788
rect 925 1724 942 1788
rect 1006 1724 1023 1788
rect 1087 1724 1104 1788
rect 1168 1724 1185 1788
rect 1249 1724 1266 1788
rect 1330 1724 1347 1788
rect 1411 1724 1428 1788
rect 1492 1724 1509 1788
rect 1573 1724 1590 1788
rect 1654 1724 1671 1788
rect 1735 1724 1752 1788
rect 1816 1724 1833 1788
rect 1897 1724 1914 1788
rect 1978 1724 1995 1788
rect 2059 1724 2076 1788
rect 2140 1724 2157 1788
rect 2221 1724 2238 1788
rect 2302 1724 2319 1788
rect 2383 1724 2400 1788
rect 2464 1724 2481 1788
rect 2545 1724 2562 1788
rect 2626 1724 2643 1788
rect 2707 1724 2724 1788
rect 2788 1724 2805 1788
rect 2869 1724 2886 1788
rect 2950 1724 2967 1788
rect 3031 1724 3048 1788
rect 3112 1724 3129 1788
rect 3193 1724 3210 1788
rect 3274 1724 3291 1788
rect 3355 1724 3372 1788
rect 3436 1724 3453 1788
rect 3517 1724 3534 1788
rect 3598 1724 3615 1788
rect 3679 1724 3696 1788
rect 3760 1724 3777 1788
rect 3841 1724 3858 1788
rect 3922 1724 3939 1788
rect 4003 1724 4020 1788
rect 4084 1724 4101 1788
rect 4165 1724 4182 1788
rect 4246 1724 4263 1788
rect 4327 1724 4344 1788
rect 4408 1724 4425 1788
rect 4489 1724 4506 1788
rect 4570 1724 4587 1788
rect 4651 1724 4668 1788
rect 4732 1724 4749 1788
rect 4813 1724 4830 1788
rect 4894 1724 4900 1788
rect 120 1702 4900 1724
rect 120 1638 126 1702
rect 190 1638 208 1702
rect 272 1638 290 1702
rect 354 1638 372 1702
rect 436 1638 454 1702
rect 518 1638 536 1702
rect 600 1638 618 1702
rect 682 1638 699 1702
rect 763 1638 780 1702
rect 844 1638 861 1702
rect 925 1638 942 1702
rect 1006 1638 1023 1702
rect 1087 1638 1104 1702
rect 1168 1638 1185 1702
rect 1249 1638 1266 1702
rect 1330 1638 1347 1702
rect 1411 1638 1428 1702
rect 1492 1638 1509 1702
rect 1573 1638 1590 1702
rect 1654 1638 1671 1702
rect 1735 1638 1752 1702
rect 1816 1638 1833 1702
rect 1897 1638 1914 1702
rect 1978 1638 1995 1702
rect 2059 1638 2076 1702
rect 2140 1638 2157 1702
rect 2221 1638 2238 1702
rect 2302 1638 2319 1702
rect 2383 1638 2400 1702
rect 2464 1638 2481 1702
rect 2545 1638 2562 1702
rect 2626 1638 2643 1702
rect 2707 1638 2724 1702
rect 2788 1638 2805 1702
rect 2869 1638 2886 1702
rect 2950 1638 2967 1702
rect 3031 1638 3048 1702
rect 3112 1638 3129 1702
rect 3193 1638 3210 1702
rect 3274 1638 3291 1702
rect 3355 1638 3372 1702
rect 3436 1638 3453 1702
rect 3517 1638 3534 1702
rect 3598 1638 3615 1702
rect 3679 1638 3696 1702
rect 3760 1638 3777 1702
rect 3841 1638 3858 1702
rect 3922 1638 3939 1702
rect 4003 1638 4020 1702
rect 4084 1638 4101 1702
rect 4165 1638 4182 1702
rect 4246 1638 4263 1702
rect 4327 1638 4344 1702
rect 4408 1638 4425 1702
rect 4489 1638 4506 1702
rect 4570 1638 4587 1702
rect 4651 1638 4668 1702
rect 4732 1638 4749 1702
rect 4813 1638 4830 1702
rect 4894 1638 4900 1702
rect 120 1616 4900 1638
rect 120 1552 126 1616
rect 190 1552 208 1616
rect 272 1552 290 1616
rect 354 1552 372 1616
rect 436 1552 454 1616
rect 518 1552 536 1616
rect 600 1552 618 1616
rect 682 1552 699 1616
rect 763 1552 780 1616
rect 844 1552 861 1616
rect 925 1552 942 1616
rect 1006 1552 1023 1616
rect 1087 1552 1104 1616
rect 1168 1552 1185 1616
rect 1249 1552 1266 1616
rect 1330 1552 1347 1616
rect 1411 1552 1428 1616
rect 1492 1552 1509 1616
rect 1573 1552 1590 1616
rect 1654 1552 1671 1616
rect 1735 1552 1752 1616
rect 1816 1552 1833 1616
rect 1897 1552 1914 1616
rect 1978 1552 1995 1616
rect 2059 1552 2076 1616
rect 2140 1552 2157 1616
rect 2221 1552 2238 1616
rect 2302 1552 2319 1616
rect 2383 1552 2400 1616
rect 2464 1552 2481 1616
rect 2545 1552 2562 1616
rect 2626 1552 2643 1616
rect 2707 1552 2724 1616
rect 2788 1552 2805 1616
rect 2869 1552 2886 1616
rect 2950 1552 2967 1616
rect 3031 1552 3048 1616
rect 3112 1552 3129 1616
rect 3193 1552 3210 1616
rect 3274 1552 3291 1616
rect 3355 1552 3372 1616
rect 3436 1552 3453 1616
rect 3517 1552 3534 1616
rect 3598 1552 3615 1616
rect 3679 1552 3696 1616
rect 3760 1552 3777 1616
rect 3841 1552 3858 1616
rect 3922 1552 3939 1616
rect 4003 1552 4020 1616
rect 4084 1552 4101 1616
rect 4165 1552 4182 1616
rect 4246 1552 4263 1616
rect 4327 1552 4344 1616
rect 4408 1552 4425 1616
rect 4489 1552 4506 1616
rect 4570 1552 4587 1616
rect 4651 1552 4668 1616
rect 4732 1552 4749 1616
rect 4813 1552 4830 1616
rect 4894 1552 4900 1616
rect 120 1530 4900 1552
rect 120 1466 126 1530
rect 190 1466 208 1530
rect 272 1466 290 1530
rect 354 1466 372 1530
rect 436 1466 454 1530
rect 518 1466 536 1530
rect 600 1466 618 1530
rect 682 1466 699 1530
rect 763 1466 780 1530
rect 844 1466 861 1530
rect 925 1466 942 1530
rect 1006 1466 1023 1530
rect 1087 1466 1104 1530
rect 1168 1466 1185 1530
rect 1249 1466 1266 1530
rect 1330 1466 1347 1530
rect 1411 1466 1428 1530
rect 1492 1466 1509 1530
rect 1573 1466 1590 1530
rect 1654 1466 1671 1530
rect 1735 1466 1752 1530
rect 1816 1466 1833 1530
rect 1897 1466 1914 1530
rect 1978 1466 1995 1530
rect 2059 1466 2076 1530
rect 2140 1466 2157 1530
rect 2221 1466 2238 1530
rect 2302 1466 2319 1530
rect 2383 1466 2400 1530
rect 2464 1466 2481 1530
rect 2545 1466 2562 1530
rect 2626 1466 2643 1530
rect 2707 1466 2724 1530
rect 2788 1466 2805 1530
rect 2869 1466 2886 1530
rect 2950 1466 2967 1530
rect 3031 1466 3048 1530
rect 3112 1466 3129 1530
rect 3193 1466 3210 1530
rect 3274 1466 3291 1530
rect 3355 1466 3372 1530
rect 3436 1466 3453 1530
rect 3517 1466 3534 1530
rect 3598 1466 3615 1530
rect 3679 1466 3696 1530
rect 3760 1466 3777 1530
rect 3841 1466 3858 1530
rect 3922 1466 3939 1530
rect 4003 1466 4020 1530
rect 4084 1466 4101 1530
rect 4165 1466 4182 1530
rect 4246 1466 4263 1530
rect 4327 1466 4344 1530
rect 4408 1466 4425 1530
rect 4489 1466 4506 1530
rect 4570 1466 4587 1530
rect 4651 1466 4668 1530
rect 4732 1466 4749 1530
rect 4813 1466 4830 1530
rect 4894 1466 4900 1530
rect 120 1444 4900 1466
rect 120 1380 126 1444
rect 190 1380 208 1444
rect 272 1380 290 1444
rect 354 1380 372 1444
rect 436 1380 454 1444
rect 518 1380 536 1444
rect 600 1380 618 1444
rect 682 1380 699 1444
rect 763 1380 780 1444
rect 844 1380 861 1444
rect 925 1380 942 1444
rect 1006 1380 1023 1444
rect 1087 1380 1104 1444
rect 1168 1380 1185 1444
rect 1249 1380 1266 1444
rect 1330 1380 1347 1444
rect 1411 1380 1428 1444
rect 1492 1380 1509 1444
rect 1573 1380 1590 1444
rect 1654 1380 1671 1444
rect 1735 1380 1752 1444
rect 1816 1380 1833 1444
rect 1897 1380 1914 1444
rect 1978 1380 1995 1444
rect 2059 1380 2076 1444
rect 2140 1380 2157 1444
rect 2221 1380 2238 1444
rect 2302 1380 2319 1444
rect 2383 1380 2400 1444
rect 2464 1380 2481 1444
rect 2545 1380 2562 1444
rect 2626 1380 2643 1444
rect 2707 1380 2724 1444
rect 2788 1380 2805 1444
rect 2869 1380 2886 1444
rect 2950 1380 2967 1444
rect 3031 1380 3048 1444
rect 3112 1380 3129 1444
rect 3193 1380 3210 1444
rect 3274 1380 3291 1444
rect 3355 1380 3372 1444
rect 3436 1380 3453 1444
rect 3517 1380 3534 1444
rect 3598 1380 3615 1444
rect 3679 1380 3696 1444
rect 3760 1380 3777 1444
rect 3841 1380 3858 1444
rect 3922 1380 3939 1444
rect 4003 1380 4020 1444
rect 4084 1380 4101 1444
rect 4165 1380 4182 1444
rect 4246 1380 4263 1444
rect 4327 1380 4344 1444
rect 4408 1380 4425 1444
rect 4489 1380 4506 1444
rect 4570 1380 4587 1444
rect 4651 1380 4668 1444
rect 4732 1380 4749 1444
rect 4813 1380 4830 1444
rect 4894 1380 4900 1444
rect 120 1378 4900 1380
rect 10151 2304 14931 2306
rect 10151 2240 10157 2304
rect 10221 2240 10239 2304
rect 10303 2240 10321 2304
rect 10385 2240 10403 2304
rect 10467 2240 10485 2304
rect 10549 2240 10567 2304
rect 10631 2240 10649 2304
rect 10713 2240 10730 2304
rect 10794 2240 10811 2304
rect 10875 2240 10892 2304
rect 10956 2240 10973 2304
rect 11037 2240 11054 2304
rect 11118 2240 11135 2304
rect 11199 2240 11216 2304
rect 11280 2240 11297 2304
rect 11361 2240 11378 2304
rect 11442 2240 11459 2304
rect 11523 2240 11540 2304
rect 11604 2240 11621 2304
rect 11685 2240 11702 2304
rect 11766 2240 11783 2304
rect 11847 2240 11864 2304
rect 11928 2240 11945 2304
rect 12009 2240 12026 2304
rect 12090 2240 12107 2304
rect 12171 2240 12188 2304
rect 12252 2240 12269 2304
rect 12333 2240 12350 2304
rect 12414 2240 12431 2304
rect 12495 2240 12512 2304
rect 12576 2240 12593 2304
rect 12657 2240 12674 2304
rect 12738 2240 12755 2304
rect 12819 2240 12836 2304
rect 12900 2240 12917 2304
rect 12981 2240 12998 2304
rect 13062 2240 13079 2304
rect 13143 2240 13160 2304
rect 13224 2240 13241 2304
rect 13305 2240 13322 2304
rect 13386 2240 13403 2304
rect 13467 2240 13484 2304
rect 13548 2240 13565 2304
rect 13629 2240 13646 2304
rect 13710 2240 13727 2304
rect 13791 2240 13808 2304
rect 13872 2240 13889 2304
rect 13953 2240 13970 2304
rect 14034 2240 14051 2304
rect 14115 2240 14132 2304
rect 14196 2240 14213 2304
rect 14277 2240 14294 2304
rect 14358 2240 14375 2304
rect 14439 2240 14456 2304
rect 14520 2240 14537 2304
rect 14601 2240 14618 2304
rect 14682 2240 14699 2304
rect 14763 2240 14780 2304
rect 14844 2240 14861 2304
rect 14925 2240 14931 2304
rect 10151 2218 14931 2240
rect 10151 2154 10157 2218
rect 10221 2154 10239 2218
rect 10303 2154 10321 2218
rect 10385 2154 10403 2218
rect 10467 2154 10485 2218
rect 10549 2154 10567 2218
rect 10631 2154 10649 2218
rect 10713 2154 10730 2218
rect 10794 2154 10811 2218
rect 10875 2154 10892 2218
rect 10956 2154 10973 2218
rect 11037 2154 11054 2218
rect 11118 2154 11135 2218
rect 11199 2154 11216 2218
rect 11280 2154 11297 2218
rect 11361 2154 11378 2218
rect 11442 2154 11459 2218
rect 11523 2154 11540 2218
rect 11604 2154 11621 2218
rect 11685 2154 11702 2218
rect 11766 2154 11783 2218
rect 11847 2154 11864 2218
rect 11928 2154 11945 2218
rect 12009 2154 12026 2218
rect 12090 2154 12107 2218
rect 12171 2154 12188 2218
rect 12252 2154 12269 2218
rect 12333 2154 12350 2218
rect 12414 2154 12431 2218
rect 12495 2154 12512 2218
rect 12576 2154 12593 2218
rect 12657 2154 12674 2218
rect 12738 2154 12755 2218
rect 12819 2154 12836 2218
rect 12900 2154 12917 2218
rect 12981 2154 12998 2218
rect 13062 2154 13079 2218
rect 13143 2154 13160 2218
rect 13224 2154 13241 2218
rect 13305 2154 13322 2218
rect 13386 2154 13403 2218
rect 13467 2154 13484 2218
rect 13548 2154 13565 2218
rect 13629 2154 13646 2218
rect 13710 2154 13727 2218
rect 13791 2154 13808 2218
rect 13872 2154 13889 2218
rect 13953 2154 13970 2218
rect 14034 2154 14051 2218
rect 14115 2154 14132 2218
rect 14196 2154 14213 2218
rect 14277 2154 14294 2218
rect 14358 2154 14375 2218
rect 14439 2154 14456 2218
rect 14520 2154 14537 2218
rect 14601 2154 14618 2218
rect 14682 2154 14699 2218
rect 14763 2154 14780 2218
rect 14844 2154 14861 2218
rect 14925 2154 14931 2218
rect 10151 2132 14931 2154
rect 10151 2068 10157 2132
rect 10221 2068 10239 2132
rect 10303 2068 10321 2132
rect 10385 2068 10403 2132
rect 10467 2068 10485 2132
rect 10549 2068 10567 2132
rect 10631 2068 10649 2132
rect 10713 2068 10730 2132
rect 10794 2068 10811 2132
rect 10875 2068 10892 2132
rect 10956 2068 10973 2132
rect 11037 2068 11054 2132
rect 11118 2068 11135 2132
rect 11199 2068 11216 2132
rect 11280 2068 11297 2132
rect 11361 2068 11378 2132
rect 11442 2068 11459 2132
rect 11523 2068 11540 2132
rect 11604 2068 11621 2132
rect 11685 2068 11702 2132
rect 11766 2068 11783 2132
rect 11847 2068 11864 2132
rect 11928 2068 11945 2132
rect 12009 2068 12026 2132
rect 12090 2068 12107 2132
rect 12171 2068 12188 2132
rect 12252 2068 12269 2132
rect 12333 2068 12350 2132
rect 12414 2068 12431 2132
rect 12495 2068 12512 2132
rect 12576 2068 12593 2132
rect 12657 2068 12674 2132
rect 12738 2068 12755 2132
rect 12819 2068 12836 2132
rect 12900 2068 12917 2132
rect 12981 2068 12998 2132
rect 13062 2068 13079 2132
rect 13143 2068 13160 2132
rect 13224 2068 13241 2132
rect 13305 2068 13322 2132
rect 13386 2068 13403 2132
rect 13467 2068 13484 2132
rect 13548 2068 13565 2132
rect 13629 2068 13646 2132
rect 13710 2068 13727 2132
rect 13791 2068 13808 2132
rect 13872 2068 13889 2132
rect 13953 2068 13970 2132
rect 14034 2068 14051 2132
rect 14115 2068 14132 2132
rect 14196 2068 14213 2132
rect 14277 2068 14294 2132
rect 14358 2068 14375 2132
rect 14439 2068 14456 2132
rect 14520 2068 14537 2132
rect 14601 2068 14618 2132
rect 14682 2068 14699 2132
rect 14763 2068 14780 2132
rect 14844 2068 14861 2132
rect 14925 2068 14931 2132
rect 10151 2046 14931 2068
rect 10151 1982 10157 2046
rect 10221 1982 10239 2046
rect 10303 1982 10321 2046
rect 10385 1982 10403 2046
rect 10467 1982 10485 2046
rect 10549 1982 10567 2046
rect 10631 1982 10649 2046
rect 10713 1982 10730 2046
rect 10794 1982 10811 2046
rect 10875 1982 10892 2046
rect 10956 1982 10973 2046
rect 11037 1982 11054 2046
rect 11118 1982 11135 2046
rect 11199 1982 11216 2046
rect 11280 1982 11297 2046
rect 11361 1982 11378 2046
rect 11442 1982 11459 2046
rect 11523 1982 11540 2046
rect 11604 1982 11621 2046
rect 11685 1982 11702 2046
rect 11766 1982 11783 2046
rect 11847 1982 11864 2046
rect 11928 1982 11945 2046
rect 12009 1982 12026 2046
rect 12090 1982 12107 2046
rect 12171 1982 12188 2046
rect 12252 1982 12269 2046
rect 12333 1982 12350 2046
rect 12414 1982 12431 2046
rect 12495 1982 12512 2046
rect 12576 1982 12593 2046
rect 12657 1982 12674 2046
rect 12738 1982 12755 2046
rect 12819 1982 12836 2046
rect 12900 1982 12917 2046
rect 12981 1982 12998 2046
rect 13062 1982 13079 2046
rect 13143 1982 13160 2046
rect 13224 1982 13241 2046
rect 13305 1982 13322 2046
rect 13386 1982 13403 2046
rect 13467 1982 13484 2046
rect 13548 1982 13565 2046
rect 13629 1982 13646 2046
rect 13710 1982 13727 2046
rect 13791 1982 13808 2046
rect 13872 1982 13889 2046
rect 13953 1982 13970 2046
rect 14034 1982 14051 2046
rect 14115 1982 14132 2046
rect 14196 1982 14213 2046
rect 14277 1982 14294 2046
rect 14358 1982 14375 2046
rect 14439 1982 14456 2046
rect 14520 1982 14537 2046
rect 14601 1982 14618 2046
rect 14682 1982 14699 2046
rect 14763 1982 14780 2046
rect 14844 1982 14861 2046
rect 14925 1982 14931 2046
rect 10151 1960 14931 1982
rect 10151 1896 10157 1960
rect 10221 1896 10239 1960
rect 10303 1896 10321 1960
rect 10385 1896 10403 1960
rect 10467 1896 10485 1960
rect 10549 1896 10567 1960
rect 10631 1896 10649 1960
rect 10713 1896 10730 1960
rect 10794 1896 10811 1960
rect 10875 1896 10892 1960
rect 10956 1896 10973 1960
rect 11037 1896 11054 1960
rect 11118 1896 11135 1960
rect 11199 1896 11216 1960
rect 11280 1896 11297 1960
rect 11361 1896 11378 1960
rect 11442 1896 11459 1960
rect 11523 1896 11540 1960
rect 11604 1896 11621 1960
rect 11685 1896 11702 1960
rect 11766 1896 11783 1960
rect 11847 1896 11864 1960
rect 11928 1896 11945 1960
rect 12009 1896 12026 1960
rect 12090 1896 12107 1960
rect 12171 1896 12188 1960
rect 12252 1896 12269 1960
rect 12333 1896 12350 1960
rect 12414 1896 12431 1960
rect 12495 1896 12512 1960
rect 12576 1896 12593 1960
rect 12657 1896 12674 1960
rect 12738 1896 12755 1960
rect 12819 1896 12836 1960
rect 12900 1896 12917 1960
rect 12981 1896 12998 1960
rect 13062 1896 13079 1960
rect 13143 1896 13160 1960
rect 13224 1896 13241 1960
rect 13305 1896 13322 1960
rect 13386 1896 13403 1960
rect 13467 1896 13484 1960
rect 13548 1896 13565 1960
rect 13629 1896 13646 1960
rect 13710 1896 13727 1960
rect 13791 1896 13808 1960
rect 13872 1896 13889 1960
rect 13953 1896 13970 1960
rect 14034 1896 14051 1960
rect 14115 1896 14132 1960
rect 14196 1896 14213 1960
rect 14277 1896 14294 1960
rect 14358 1896 14375 1960
rect 14439 1896 14456 1960
rect 14520 1896 14537 1960
rect 14601 1896 14618 1960
rect 14682 1896 14699 1960
rect 14763 1896 14780 1960
rect 14844 1896 14861 1960
rect 14925 1896 14931 1960
rect 10151 1874 14931 1896
rect 10151 1810 10157 1874
rect 10221 1810 10239 1874
rect 10303 1810 10321 1874
rect 10385 1810 10403 1874
rect 10467 1810 10485 1874
rect 10549 1810 10567 1874
rect 10631 1810 10649 1874
rect 10713 1810 10730 1874
rect 10794 1810 10811 1874
rect 10875 1810 10892 1874
rect 10956 1810 10973 1874
rect 11037 1810 11054 1874
rect 11118 1810 11135 1874
rect 11199 1810 11216 1874
rect 11280 1810 11297 1874
rect 11361 1810 11378 1874
rect 11442 1810 11459 1874
rect 11523 1810 11540 1874
rect 11604 1810 11621 1874
rect 11685 1810 11702 1874
rect 11766 1810 11783 1874
rect 11847 1810 11864 1874
rect 11928 1810 11945 1874
rect 12009 1810 12026 1874
rect 12090 1810 12107 1874
rect 12171 1810 12188 1874
rect 12252 1810 12269 1874
rect 12333 1810 12350 1874
rect 12414 1810 12431 1874
rect 12495 1810 12512 1874
rect 12576 1810 12593 1874
rect 12657 1810 12674 1874
rect 12738 1810 12755 1874
rect 12819 1810 12836 1874
rect 12900 1810 12917 1874
rect 12981 1810 12998 1874
rect 13062 1810 13079 1874
rect 13143 1810 13160 1874
rect 13224 1810 13241 1874
rect 13305 1810 13322 1874
rect 13386 1810 13403 1874
rect 13467 1810 13484 1874
rect 13548 1810 13565 1874
rect 13629 1810 13646 1874
rect 13710 1810 13727 1874
rect 13791 1810 13808 1874
rect 13872 1810 13889 1874
rect 13953 1810 13970 1874
rect 14034 1810 14051 1874
rect 14115 1810 14132 1874
rect 14196 1810 14213 1874
rect 14277 1810 14294 1874
rect 14358 1810 14375 1874
rect 14439 1810 14456 1874
rect 14520 1810 14537 1874
rect 14601 1810 14618 1874
rect 14682 1810 14699 1874
rect 14763 1810 14780 1874
rect 14844 1810 14861 1874
rect 14925 1810 14931 1874
rect 10151 1788 14931 1810
rect 10151 1724 10157 1788
rect 10221 1724 10239 1788
rect 10303 1724 10321 1788
rect 10385 1724 10403 1788
rect 10467 1724 10485 1788
rect 10549 1724 10567 1788
rect 10631 1724 10649 1788
rect 10713 1724 10730 1788
rect 10794 1724 10811 1788
rect 10875 1724 10892 1788
rect 10956 1724 10973 1788
rect 11037 1724 11054 1788
rect 11118 1724 11135 1788
rect 11199 1724 11216 1788
rect 11280 1724 11297 1788
rect 11361 1724 11378 1788
rect 11442 1724 11459 1788
rect 11523 1724 11540 1788
rect 11604 1724 11621 1788
rect 11685 1724 11702 1788
rect 11766 1724 11783 1788
rect 11847 1724 11864 1788
rect 11928 1724 11945 1788
rect 12009 1724 12026 1788
rect 12090 1724 12107 1788
rect 12171 1724 12188 1788
rect 12252 1724 12269 1788
rect 12333 1724 12350 1788
rect 12414 1724 12431 1788
rect 12495 1724 12512 1788
rect 12576 1724 12593 1788
rect 12657 1724 12674 1788
rect 12738 1724 12755 1788
rect 12819 1724 12836 1788
rect 12900 1724 12917 1788
rect 12981 1724 12998 1788
rect 13062 1724 13079 1788
rect 13143 1724 13160 1788
rect 13224 1724 13241 1788
rect 13305 1724 13322 1788
rect 13386 1724 13403 1788
rect 13467 1724 13484 1788
rect 13548 1724 13565 1788
rect 13629 1724 13646 1788
rect 13710 1724 13727 1788
rect 13791 1724 13808 1788
rect 13872 1724 13889 1788
rect 13953 1724 13970 1788
rect 14034 1724 14051 1788
rect 14115 1724 14132 1788
rect 14196 1724 14213 1788
rect 14277 1724 14294 1788
rect 14358 1724 14375 1788
rect 14439 1724 14456 1788
rect 14520 1724 14537 1788
rect 14601 1724 14618 1788
rect 14682 1724 14699 1788
rect 14763 1724 14780 1788
rect 14844 1724 14861 1788
rect 14925 1724 14931 1788
rect 10151 1702 14931 1724
rect 10151 1638 10157 1702
rect 10221 1638 10239 1702
rect 10303 1638 10321 1702
rect 10385 1638 10403 1702
rect 10467 1638 10485 1702
rect 10549 1638 10567 1702
rect 10631 1638 10649 1702
rect 10713 1638 10730 1702
rect 10794 1638 10811 1702
rect 10875 1638 10892 1702
rect 10956 1638 10973 1702
rect 11037 1638 11054 1702
rect 11118 1638 11135 1702
rect 11199 1638 11216 1702
rect 11280 1638 11297 1702
rect 11361 1638 11378 1702
rect 11442 1638 11459 1702
rect 11523 1638 11540 1702
rect 11604 1638 11621 1702
rect 11685 1638 11702 1702
rect 11766 1638 11783 1702
rect 11847 1638 11864 1702
rect 11928 1638 11945 1702
rect 12009 1638 12026 1702
rect 12090 1638 12107 1702
rect 12171 1638 12188 1702
rect 12252 1638 12269 1702
rect 12333 1638 12350 1702
rect 12414 1638 12431 1702
rect 12495 1638 12512 1702
rect 12576 1638 12593 1702
rect 12657 1638 12674 1702
rect 12738 1638 12755 1702
rect 12819 1638 12836 1702
rect 12900 1638 12917 1702
rect 12981 1638 12998 1702
rect 13062 1638 13079 1702
rect 13143 1638 13160 1702
rect 13224 1638 13241 1702
rect 13305 1638 13322 1702
rect 13386 1638 13403 1702
rect 13467 1638 13484 1702
rect 13548 1638 13565 1702
rect 13629 1638 13646 1702
rect 13710 1638 13727 1702
rect 13791 1638 13808 1702
rect 13872 1638 13889 1702
rect 13953 1638 13970 1702
rect 14034 1638 14051 1702
rect 14115 1638 14132 1702
rect 14196 1638 14213 1702
rect 14277 1638 14294 1702
rect 14358 1638 14375 1702
rect 14439 1638 14456 1702
rect 14520 1638 14537 1702
rect 14601 1638 14618 1702
rect 14682 1638 14699 1702
rect 14763 1638 14780 1702
rect 14844 1638 14861 1702
rect 14925 1638 14931 1702
rect 10151 1616 14931 1638
rect 10151 1552 10157 1616
rect 10221 1552 10239 1616
rect 10303 1552 10321 1616
rect 10385 1552 10403 1616
rect 10467 1552 10485 1616
rect 10549 1552 10567 1616
rect 10631 1552 10649 1616
rect 10713 1552 10730 1616
rect 10794 1552 10811 1616
rect 10875 1552 10892 1616
rect 10956 1552 10973 1616
rect 11037 1552 11054 1616
rect 11118 1552 11135 1616
rect 11199 1552 11216 1616
rect 11280 1552 11297 1616
rect 11361 1552 11378 1616
rect 11442 1552 11459 1616
rect 11523 1552 11540 1616
rect 11604 1552 11621 1616
rect 11685 1552 11702 1616
rect 11766 1552 11783 1616
rect 11847 1552 11864 1616
rect 11928 1552 11945 1616
rect 12009 1552 12026 1616
rect 12090 1552 12107 1616
rect 12171 1552 12188 1616
rect 12252 1552 12269 1616
rect 12333 1552 12350 1616
rect 12414 1552 12431 1616
rect 12495 1552 12512 1616
rect 12576 1552 12593 1616
rect 12657 1552 12674 1616
rect 12738 1552 12755 1616
rect 12819 1552 12836 1616
rect 12900 1552 12917 1616
rect 12981 1552 12998 1616
rect 13062 1552 13079 1616
rect 13143 1552 13160 1616
rect 13224 1552 13241 1616
rect 13305 1552 13322 1616
rect 13386 1552 13403 1616
rect 13467 1552 13484 1616
rect 13548 1552 13565 1616
rect 13629 1552 13646 1616
rect 13710 1552 13727 1616
rect 13791 1552 13808 1616
rect 13872 1552 13889 1616
rect 13953 1552 13970 1616
rect 14034 1552 14051 1616
rect 14115 1552 14132 1616
rect 14196 1552 14213 1616
rect 14277 1552 14294 1616
rect 14358 1552 14375 1616
rect 14439 1552 14456 1616
rect 14520 1552 14537 1616
rect 14601 1552 14618 1616
rect 14682 1552 14699 1616
rect 14763 1552 14780 1616
rect 14844 1552 14861 1616
rect 14925 1552 14931 1616
rect 10151 1530 14931 1552
rect 10151 1466 10157 1530
rect 10221 1466 10239 1530
rect 10303 1466 10321 1530
rect 10385 1466 10403 1530
rect 10467 1466 10485 1530
rect 10549 1466 10567 1530
rect 10631 1466 10649 1530
rect 10713 1466 10730 1530
rect 10794 1466 10811 1530
rect 10875 1466 10892 1530
rect 10956 1466 10973 1530
rect 11037 1466 11054 1530
rect 11118 1466 11135 1530
rect 11199 1466 11216 1530
rect 11280 1466 11297 1530
rect 11361 1466 11378 1530
rect 11442 1466 11459 1530
rect 11523 1466 11540 1530
rect 11604 1466 11621 1530
rect 11685 1466 11702 1530
rect 11766 1466 11783 1530
rect 11847 1466 11864 1530
rect 11928 1466 11945 1530
rect 12009 1466 12026 1530
rect 12090 1466 12107 1530
rect 12171 1466 12188 1530
rect 12252 1466 12269 1530
rect 12333 1466 12350 1530
rect 12414 1466 12431 1530
rect 12495 1466 12512 1530
rect 12576 1466 12593 1530
rect 12657 1466 12674 1530
rect 12738 1466 12755 1530
rect 12819 1466 12836 1530
rect 12900 1466 12917 1530
rect 12981 1466 12998 1530
rect 13062 1466 13079 1530
rect 13143 1466 13160 1530
rect 13224 1466 13241 1530
rect 13305 1466 13322 1530
rect 13386 1466 13403 1530
rect 13467 1466 13484 1530
rect 13548 1466 13565 1530
rect 13629 1466 13646 1530
rect 13710 1466 13727 1530
rect 13791 1466 13808 1530
rect 13872 1466 13889 1530
rect 13953 1466 13970 1530
rect 14034 1466 14051 1530
rect 14115 1466 14132 1530
rect 14196 1466 14213 1530
rect 14277 1466 14294 1530
rect 14358 1466 14375 1530
rect 14439 1466 14456 1530
rect 14520 1466 14537 1530
rect 14601 1466 14618 1530
rect 14682 1466 14699 1530
rect 14763 1466 14780 1530
rect 14844 1466 14861 1530
rect 14925 1466 14931 1530
rect 10151 1444 14931 1466
rect 10151 1380 10157 1444
rect 10221 1380 10239 1444
rect 10303 1380 10321 1444
rect 10385 1380 10403 1444
rect 10467 1380 10485 1444
rect 10549 1380 10567 1444
rect 10631 1380 10649 1444
rect 10713 1380 10730 1444
rect 10794 1380 10811 1444
rect 10875 1380 10892 1444
rect 10956 1380 10973 1444
rect 11037 1380 11054 1444
rect 11118 1380 11135 1444
rect 11199 1380 11216 1444
rect 11280 1380 11297 1444
rect 11361 1380 11378 1444
rect 11442 1380 11459 1444
rect 11523 1380 11540 1444
rect 11604 1380 11621 1444
rect 11685 1380 11702 1444
rect 11766 1380 11783 1444
rect 11847 1380 11864 1444
rect 11928 1380 11945 1444
rect 12009 1380 12026 1444
rect 12090 1380 12107 1444
rect 12171 1380 12188 1444
rect 12252 1380 12269 1444
rect 12333 1380 12350 1444
rect 12414 1380 12431 1444
rect 12495 1380 12512 1444
rect 12576 1380 12593 1444
rect 12657 1380 12674 1444
rect 12738 1380 12755 1444
rect 12819 1380 12836 1444
rect 12900 1380 12917 1444
rect 12981 1380 12998 1444
rect 13062 1380 13079 1444
rect 13143 1380 13160 1444
rect 13224 1380 13241 1444
rect 13305 1380 13322 1444
rect 13386 1380 13403 1444
rect 13467 1380 13484 1444
rect 13548 1380 13565 1444
rect 13629 1380 13646 1444
rect 13710 1380 13727 1444
rect 13791 1380 13808 1444
rect 13872 1380 13889 1444
rect 13953 1380 13970 1444
rect 14034 1380 14051 1444
rect 14115 1380 14132 1444
rect 14196 1380 14213 1444
rect 14277 1380 14294 1444
rect 14358 1380 14375 1444
rect 14439 1380 14456 1444
rect 14520 1380 14537 1444
rect 14601 1380 14618 1444
rect 14682 1380 14699 1444
rect 14763 1380 14780 1444
rect 14844 1380 14861 1444
rect 14925 1380 14931 1444
rect 10151 1378 14931 1380
<< via3 >>
rect 126 2240 190 2304
rect 208 2240 272 2304
rect 290 2240 354 2304
rect 372 2240 436 2304
rect 454 2240 518 2304
rect 536 2240 600 2304
rect 618 2240 682 2304
rect 699 2240 763 2304
rect 780 2240 844 2304
rect 861 2240 925 2304
rect 942 2240 1006 2304
rect 1023 2240 1087 2304
rect 1104 2240 1168 2304
rect 1185 2240 1249 2304
rect 1266 2240 1330 2304
rect 1347 2240 1411 2304
rect 1428 2240 1492 2304
rect 1509 2240 1573 2304
rect 1590 2240 1654 2304
rect 1671 2240 1735 2304
rect 1752 2240 1816 2304
rect 1833 2240 1897 2304
rect 1914 2240 1978 2304
rect 1995 2240 2059 2304
rect 2076 2240 2140 2304
rect 2157 2240 2221 2304
rect 2238 2240 2302 2304
rect 2319 2240 2383 2304
rect 2400 2240 2464 2304
rect 2481 2240 2545 2304
rect 2562 2240 2626 2304
rect 2643 2240 2707 2304
rect 2724 2240 2788 2304
rect 2805 2240 2869 2304
rect 2886 2240 2950 2304
rect 2967 2240 3031 2304
rect 3048 2240 3112 2304
rect 3129 2240 3193 2304
rect 3210 2240 3274 2304
rect 3291 2240 3355 2304
rect 3372 2240 3436 2304
rect 3453 2240 3517 2304
rect 3534 2240 3598 2304
rect 3615 2240 3679 2304
rect 3696 2240 3760 2304
rect 3777 2240 3841 2304
rect 3858 2240 3922 2304
rect 3939 2240 4003 2304
rect 4020 2240 4084 2304
rect 4101 2240 4165 2304
rect 4182 2240 4246 2304
rect 4263 2240 4327 2304
rect 4344 2240 4408 2304
rect 4425 2240 4489 2304
rect 4506 2240 4570 2304
rect 4587 2240 4651 2304
rect 4668 2240 4732 2304
rect 4749 2240 4813 2304
rect 4830 2240 4894 2304
rect 126 2154 190 2218
rect 208 2154 272 2218
rect 290 2154 354 2218
rect 372 2154 436 2218
rect 454 2154 518 2218
rect 536 2154 600 2218
rect 618 2154 682 2218
rect 699 2154 763 2218
rect 780 2154 844 2218
rect 861 2154 925 2218
rect 942 2154 1006 2218
rect 1023 2154 1087 2218
rect 1104 2154 1168 2218
rect 1185 2154 1249 2218
rect 1266 2154 1330 2218
rect 1347 2154 1411 2218
rect 1428 2154 1492 2218
rect 1509 2154 1573 2218
rect 1590 2154 1654 2218
rect 1671 2154 1735 2218
rect 1752 2154 1816 2218
rect 1833 2154 1897 2218
rect 1914 2154 1978 2218
rect 1995 2154 2059 2218
rect 2076 2154 2140 2218
rect 2157 2154 2221 2218
rect 2238 2154 2302 2218
rect 2319 2154 2383 2218
rect 2400 2154 2464 2218
rect 2481 2154 2545 2218
rect 2562 2154 2626 2218
rect 2643 2154 2707 2218
rect 2724 2154 2788 2218
rect 2805 2154 2869 2218
rect 2886 2154 2950 2218
rect 2967 2154 3031 2218
rect 3048 2154 3112 2218
rect 3129 2154 3193 2218
rect 3210 2154 3274 2218
rect 3291 2154 3355 2218
rect 3372 2154 3436 2218
rect 3453 2154 3517 2218
rect 3534 2154 3598 2218
rect 3615 2154 3679 2218
rect 3696 2154 3760 2218
rect 3777 2154 3841 2218
rect 3858 2154 3922 2218
rect 3939 2154 4003 2218
rect 4020 2154 4084 2218
rect 4101 2154 4165 2218
rect 4182 2154 4246 2218
rect 4263 2154 4327 2218
rect 4344 2154 4408 2218
rect 4425 2154 4489 2218
rect 4506 2154 4570 2218
rect 4587 2154 4651 2218
rect 4668 2154 4732 2218
rect 4749 2154 4813 2218
rect 4830 2154 4894 2218
rect 126 2068 190 2132
rect 208 2068 272 2132
rect 290 2068 354 2132
rect 372 2068 436 2132
rect 454 2068 518 2132
rect 536 2068 600 2132
rect 618 2068 682 2132
rect 699 2068 763 2132
rect 780 2068 844 2132
rect 861 2068 925 2132
rect 942 2068 1006 2132
rect 1023 2068 1087 2132
rect 1104 2068 1168 2132
rect 1185 2068 1249 2132
rect 1266 2068 1330 2132
rect 1347 2068 1411 2132
rect 1428 2068 1492 2132
rect 1509 2068 1573 2132
rect 1590 2068 1654 2132
rect 1671 2068 1735 2132
rect 1752 2068 1816 2132
rect 1833 2068 1897 2132
rect 1914 2068 1978 2132
rect 1995 2068 2059 2132
rect 2076 2068 2140 2132
rect 2157 2068 2221 2132
rect 2238 2068 2302 2132
rect 2319 2068 2383 2132
rect 2400 2068 2464 2132
rect 2481 2068 2545 2132
rect 2562 2068 2626 2132
rect 2643 2068 2707 2132
rect 2724 2068 2788 2132
rect 2805 2068 2869 2132
rect 2886 2068 2950 2132
rect 2967 2068 3031 2132
rect 3048 2068 3112 2132
rect 3129 2068 3193 2132
rect 3210 2068 3274 2132
rect 3291 2068 3355 2132
rect 3372 2068 3436 2132
rect 3453 2068 3517 2132
rect 3534 2068 3598 2132
rect 3615 2068 3679 2132
rect 3696 2068 3760 2132
rect 3777 2068 3841 2132
rect 3858 2068 3922 2132
rect 3939 2068 4003 2132
rect 4020 2068 4084 2132
rect 4101 2068 4165 2132
rect 4182 2068 4246 2132
rect 4263 2068 4327 2132
rect 4344 2068 4408 2132
rect 4425 2068 4489 2132
rect 4506 2068 4570 2132
rect 4587 2068 4651 2132
rect 4668 2068 4732 2132
rect 4749 2068 4813 2132
rect 4830 2068 4894 2132
rect 126 1982 190 2046
rect 208 1982 272 2046
rect 290 1982 354 2046
rect 372 1982 436 2046
rect 454 1982 518 2046
rect 536 1982 600 2046
rect 618 1982 682 2046
rect 699 1982 763 2046
rect 780 1982 844 2046
rect 861 1982 925 2046
rect 942 1982 1006 2046
rect 1023 1982 1087 2046
rect 1104 1982 1168 2046
rect 1185 1982 1249 2046
rect 1266 1982 1330 2046
rect 1347 1982 1411 2046
rect 1428 1982 1492 2046
rect 1509 1982 1573 2046
rect 1590 1982 1654 2046
rect 1671 1982 1735 2046
rect 1752 1982 1816 2046
rect 1833 1982 1897 2046
rect 1914 1982 1978 2046
rect 1995 1982 2059 2046
rect 2076 1982 2140 2046
rect 2157 1982 2221 2046
rect 2238 1982 2302 2046
rect 2319 1982 2383 2046
rect 2400 1982 2464 2046
rect 2481 1982 2545 2046
rect 2562 1982 2626 2046
rect 2643 1982 2707 2046
rect 2724 1982 2788 2046
rect 2805 1982 2869 2046
rect 2886 1982 2950 2046
rect 2967 1982 3031 2046
rect 3048 1982 3112 2046
rect 3129 1982 3193 2046
rect 3210 1982 3274 2046
rect 3291 1982 3355 2046
rect 3372 1982 3436 2046
rect 3453 1982 3517 2046
rect 3534 1982 3598 2046
rect 3615 1982 3679 2046
rect 3696 1982 3760 2046
rect 3777 1982 3841 2046
rect 3858 1982 3922 2046
rect 3939 1982 4003 2046
rect 4020 1982 4084 2046
rect 4101 1982 4165 2046
rect 4182 1982 4246 2046
rect 4263 1982 4327 2046
rect 4344 1982 4408 2046
rect 4425 1982 4489 2046
rect 4506 1982 4570 2046
rect 4587 1982 4651 2046
rect 4668 1982 4732 2046
rect 4749 1982 4813 2046
rect 4830 1982 4894 2046
rect 126 1896 190 1960
rect 208 1896 272 1960
rect 290 1896 354 1960
rect 372 1896 436 1960
rect 454 1896 518 1960
rect 536 1896 600 1960
rect 618 1896 682 1960
rect 699 1896 763 1960
rect 780 1896 844 1960
rect 861 1896 925 1960
rect 942 1896 1006 1960
rect 1023 1896 1087 1960
rect 1104 1896 1168 1960
rect 1185 1896 1249 1960
rect 1266 1896 1330 1960
rect 1347 1896 1411 1960
rect 1428 1896 1492 1960
rect 1509 1896 1573 1960
rect 1590 1896 1654 1960
rect 1671 1896 1735 1960
rect 1752 1896 1816 1960
rect 1833 1896 1897 1960
rect 1914 1896 1978 1960
rect 1995 1896 2059 1960
rect 2076 1896 2140 1960
rect 2157 1896 2221 1960
rect 2238 1896 2302 1960
rect 2319 1896 2383 1960
rect 2400 1896 2464 1960
rect 2481 1896 2545 1960
rect 2562 1896 2626 1960
rect 2643 1896 2707 1960
rect 2724 1896 2788 1960
rect 2805 1896 2869 1960
rect 2886 1896 2950 1960
rect 2967 1896 3031 1960
rect 3048 1896 3112 1960
rect 3129 1896 3193 1960
rect 3210 1896 3274 1960
rect 3291 1896 3355 1960
rect 3372 1896 3436 1960
rect 3453 1896 3517 1960
rect 3534 1896 3598 1960
rect 3615 1896 3679 1960
rect 3696 1896 3760 1960
rect 3777 1896 3841 1960
rect 3858 1896 3922 1960
rect 3939 1896 4003 1960
rect 4020 1896 4084 1960
rect 4101 1896 4165 1960
rect 4182 1896 4246 1960
rect 4263 1896 4327 1960
rect 4344 1896 4408 1960
rect 4425 1896 4489 1960
rect 4506 1896 4570 1960
rect 4587 1896 4651 1960
rect 4668 1896 4732 1960
rect 4749 1896 4813 1960
rect 4830 1896 4894 1960
rect 126 1810 190 1874
rect 208 1810 272 1874
rect 290 1810 354 1874
rect 372 1810 436 1874
rect 454 1810 518 1874
rect 536 1810 600 1874
rect 618 1810 682 1874
rect 699 1810 763 1874
rect 780 1810 844 1874
rect 861 1810 925 1874
rect 942 1810 1006 1874
rect 1023 1810 1087 1874
rect 1104 1810 1168 1874
rect 1185 1810 1249 1874
rect 1266 1810 1330 1874
rect 1347 1810 1411 1874
rect 1428 1810 1492 1874
rect 1509 1810 1573 1874
rect 1590 1810 1654 1874
rect 1671 1810 1735 1874
rect 1752 1810 1816 1874
rect 1833 1810 1897 1874
rect 1914 1810 1978 1874
rect 1995 1810 2059 1874
rect 2076 1810 2140 1874
rect 2157 1810 2221 1874
rect 2238 1810 2302 1874
rect 2319 1810 2383 1874
rect 2400 1810 2464 1874
rect 2481 1810 2545 1874
rect 2562 1810 2626 1874
rect 2643 1810 2707 1874
rect 2724 1810 2788 1874
rect 2805 1810 2869 1874
rect 2886 1810 2950 1874
rect 2967 1810 3031 1874
rect 3048 1810 3112 1874
rect 3129 1810 3193 1874
rect 3210 1810 3274 1874
rect 3291 1810 3355 1874
rect 3372 1810 3436 1874
rect 3453 1810 3517 1874
rect 3534 1810 3598 1874
rect 3615 1810 3679 1874
rect 3696 1810 3760 1874
rect 3777 1810 3841 1874
rect 3858 1810 3922 1874
rect 3939 1810 4003 1874
rect 4020 1810 4084 1874
rect 4101 1810 4165 1874
rect 4182 1810 4246 1874
rect 4263 1810 4327 1874
rect 4344 1810 4408 1874
rect 4425 1810 4489 1874
rect 4506 1810 4570 1874
rect 4587 1810 4651 1874
rect 4668 1810 4732 1874
rect 4749 1810 4813 1874
rect 4830 1810 4894 1874
rect 126 1724 190 1788
rect 208 1724 272 1788
rect 290 1724 354 1788
rect 372 1724 436 1788
rect 454 1724 518 1788
rect 536 1724 600 1788
rect 618 1724 682 1788
rect 699 1724 763 1788
rect 780 1724 844 1788
rect 861 1724 925 1788
rect 942 1724 1006 1788
rect 1023 1724 1087 1788
rect 1104 1724 1168 1788
rect 1185 1724 1249 1788
rect 1266 1724 1330 1788
rect 1347 1724 1411 1788
rect 1428 1724 1492 1788
rect 1509 1724 1573 1788
rect 1590 1724 1654 1788
rect 1671 1724 1735 1788
rect 1752 1724 1816 1788
rect 1833 1724 1897 1788
rect 1914 1724 1978 1788
rect 1995 1724 2059 1788
rect 2076 1724 2140 1788
rect 2157 1724 2221 1788
rect 2238 1724 2302 1788
rect 2319 1724 2383 1788
rect 2400 1724 2464 1788
rect 2481 1724 2545 1788
rect 2562 1724 2626 1788
rect 2643 1724 2707 1788
rect 2724 1724 2788 1788
rect 2805 1724 2869 1788
rect 2886 1724 2950 1788
rect 2967 1724 3031 1788
rect 3048 1724 3112 1788
rect 3129 1724 3193 1788
rect 3210 1724 3274 1788
rect 3291 1724 3355 1788
rect 3372 1724 3436 1788
rect 3453 1724 3517 1788
rect 3534 1724 3598 1788
rect 3615 1724 3679 1788
rect 3696 1724 3760 1788
rect 3777 1724 3841 1788
rect 3858 1724 3922 1788
rect 3939 1724 4003 1788
rect 4020 1724 4084 1788
rect 4101 1724 4165 1788
rect 4182 1724 4246 1788
rect 4263 1724 4327 1788
rect 4344 1724 4408 1788
rect 4425 1724 4489 1788
rect 4506 1724 4570 1788
rect 4587 1724 4651 1788
rect 4668 1724 4732 1788
rect 4749 1724 4813 1788
rect 4830 1724 4894 1788
rect 126 1638 190 1702
rect 208 1638 272 1702
rect 290 1638 354 1702
rect 372 1638 436 1702
rect 454 1638 518 1702
rect 536 1638 600 1702
rect 618 1638 682 1702
rect 699 1638 763 1702
rect 780 1638 844 1702
rect 861 1638 925 1702
rect 942 1638 1006 1702
rect 1023 1638 1087 1702
rect 1104 1638 1168 1702
rect 1185 1638 1249 1702
rect 1266 1638 1330 1702
rect 1347 1638 1411 1702
rect 1428 1638 1492 1702
rect 1509 1638 1573 1702
rect 1590 1638 1654 1702
rect 1671 1638 1735 1702
rect 1752 1638 1816 1702
rect 1833 1638 1897 1702
rect 1914 1638 1978 1702
rect 1995 1638 2059 1702
rect 2076 1638 2140 1702
rect 2157 1638 2221 1702
rect 2238 1638 2302 1702
rect 2319 1638 2383 1702
rect 2400 1638 2464 1702
rect 2481 1638 2545 1702
rect 2562 1638 2626 1702
rect 2643 1638 2707 1702
rect 2724 1638 2788 1702
rect 2805 1638 2869 1702
rect 2886 1638 2950 1702
rect 2967 1638 3031 1702
rect 3048 1638 3112 1702
rect 3129 1638 3193 1702
rect 3210 1638 3274 1702
rect 3291 1638 3355 1702
rect 3372 1638 3436 1702
rect 3453 1638 3517 1702
rect 3534 1638 3598 1702
rect 3615 1638 3679 1702
rect 3696 1638 3760 1702
rect 3777 1638 3841 1702
rect 3858 1638 3922 1702
rect 3939 1638 4003 1702
rect 4020 1638 4084 1702
rect 4101 1638 4165 1702
rect 4182 1638 4246 1702
rect 4263 1638 4327 1702
rect 4344 1638 4408 1702
rect 4425 1638 4489 1702
rect 4506 1638 4570 1702
rect 4587 1638 4651 1702
rect 4668 1638 4732 1702
rect 4749 1638 4813 1702
rect 4830 1638 4894 1702
rect 126 1552 190 1616
rect 208 1552 272 1616
rect 290 1552 354 1616
rect 372 1552 436 1616
rect 454 1552 518 1616
rect 536 1552 600 1616
rect 618 1552 682 1616
rect 699 1552 763 1616
rect 780 1552 844 1616
rect 861 1552 925 1616
rect 942 1552 1006 1616
rect 1023 1552 1087 1616
rect 1104 1552 1168 1616
rect 1185 1552 1249 1616
rect 1266 1552 1330 1616
rect 1347 1552 1411 1616
rect 1428 1552 1492 1616
rect 1509 1552 1573 1616
rect 1590 1552 1654 1616
rect 1671 1552 1735 1616
rect 1752 1552 1816 1616
rect 1833 1552 1897 1616
rect 1914 1552 1978 1616
rect 1995 1552 2059 1616
rect 2076 1552 2140 1616
rect 2157 1552 2221 1616
rect 2238 1552 2302 1616
rect 2319 1552 2383 1616
rect 2400 1552 2464 1616
rect 2481 1552 2545 1616
rect 2562 1552 2626 1616
rect 2643 1552 2707 1616
rect 2724 1552 2788 1616
rect 2805 1552 2869 1616
rect 2886 1552 2950 1616
rect 2967 1552 3031 1616
rect 3048 1552 3112 1616
rect 3129 1552 3193 1616
rect 3210 1552 3274 1616
rect 3291 1552 3355 1616
rect 3372 1552 3436 1616
rect 3453 1552 3517 1616
rect 3534 1552 3598 1616
rect 3615 1552 3679 1616
rect 3696 1552 3760 1616
rect 3777 1552 3841 1616
rect 3858 1552 3922 1616
rect 3939 1552 4003 1616
rect 4020 1552 4084 1616
rect 4101 1552 4165 1616
rect 4182 1552 4246 1616
rect 4263 1552 4327 1616
rect 4344 1552 4408 1616
rect 4425 1552 4489 1616
rect 4506 1552 4570 1616
rect 4587 1552 4651 1616
rect 4668 1552 4732 1616
rect 4749 1552 4813 1616
rect 4830 1552 4894 1616
rect 126 1466 190 1530
rect 208 1466 272 1530
rect 290 1466 354 1530
rect 372 1466 436 1530
rect 454 1466 518 1530
rect 536 1466 600 1530
rect 618 1466 682 1530
rect 699 1466 763 1530
rect 780 1466 844 1530
rect 861 1466 925 1530
rect 942 1466 1006 1530
rect 1023 1466 1087 1530
rect 1104 1466 1168 1530
rect 1185 1466 1249 1530
rect 1266 1466 1330 1530
rect 1347 1466 1411 1530
rect 1428 1466 1492 1530
rect 1509 1466 1573 1530
rect 1590 1466 1654 1530
rect 1671 1466 1735 1530
rect 1752 1466 1816 1530
rect 1833 1466 1897 1530
rect 1914 1466 1978 1530
rect 1995 1466 2059 1530
rect 2076 1466 2140 1530
rect 2157 1466 2221 1530
rect 2238 1466 2302 1530
rect 2319 1466 2383 1530
rect 2400 1466 2464 1530
rect 2481 1466 2545 1530
rect 2562 1466 2626 1530
rect 2643 1466 2707 1530
rect 2724 1466 2788 1530
rect 2805 1466 2869 1530
rect 2886 1466 2950 1530
rect 2967 1466 3031 1530
rect 3048 1466 3112 1530
rect 3129 1466 3193 1530
rect 3210 1466 3274 1530
rect 3291 1466 3355 1530
rect 3372 1466 3436 1530
rect 3453 1466 3517 1530
rect 3534 1466 3598 1530
rect 3615 1466 3679 1530
rect 3696 1466 3760 1530
rect 3777 1466 3841 1530
rect 3858 1466 3922 1530
rect 3939 1466 4003 1530
rect 4020 1466 4084 1530
rect 4101 1466 4165 1530
rect 4182 1466 4246 1530
rect 4263 1466 4327 1530
rect 4344 1466 4408 1530
rect 4425 1466 4489 1530
rect 4506 1466 4570 1530
rect 4587 1466 4651 1530
rect 4668 1466 4732 1530
rect 4749 1466 4813 1530
rect 4830 1466 4894 1530
rect 126 1380 190 1444
rect 208 1380 272 1444
rect 290 1380 354 1444
rect 372 1380 436 1444
rect 454 1380 518 1444
rect 536 1380 600 1444
rect 618 1380 682 1444
rect 699 1380 763 1444
rect 780 1380 844 1444
rect 861 1380 925 1444
rect 942 1380 1006 1444
rect 1023 1380 1087 1444
rect 1104 1380 1168 1444
rect 1185 1380 1249 1444
rect 1266 1380 1330 1444
rect 1347 1380 1411 1444
rect 1428 1380 1492 1444
rect 1509 1380 1573 1444
rect 1590 1380 1654 1444
rect 1671 1380 1735 1444
rect 1752 1380 1816 1444
rect 1833 1380 1897 1444
rect 1914 1380 1978 1444
rect 1995 1380 2059 1444
rect 2076 1380 2140 1444
rect 2157 1380 2221 1444
rect 2238 1380 2302 1444
rect 2319 1380 2383 1444
rect 2400 1380 2464 1444
rect 2481 1380 2545 1444
rect 2562 1380 2626 1444
rect 2643 1380 2707 1444
rect 2724 1380 2788 1444
rect 2805 1380 2869 1444
rect 2886 1380 2950 1444
rect 2967 1380 3031 1444
rect 3048 1380 3112 1444
rect 3129 1380 3193 1444
rect 3210 1380 3274 1444
rect 3291 1380 3355 1444
rect 3372 1380 3436 1444
rect 3453 1380 3517 1444
rect 3534 1380 3598 1444
rect 3615 1380 3679 1444
rect 3696 1380 3760 1444
rect 3777 1380 3841 1444
rect 3858 1380 3922 1444
rect 3939 1380 4003 1444
rect 4020 1380 4084 1444
rect 4101 1380 4165 1444
rect 4182 1380 4246 1444
rect 4263 1380 4327 1444
rect 4344 1380 4408 1444
rect 4425 1380 4489 1444
rect 4506 1380 4570 1444
rect 4587 1380 4651 1444
rect 4668 1380 4732 1444
rect 4749 1380 4813 1444
rect 4830 1380 4894 1444
rect 10157 2240 10221 2304
rect 10239 2240 10303 2304
rect 10321 2240 10385 2304
rect 10403 2240 10467 2304
rect 10485 2240 10549 2304
rect 10567 2240 10631 2304
rect 10649 2240 10713 2304
rect 10730 2240 10794 2304
rect 10811 2240 10875 2304
rect 10892 2240 10956 2304
rect 10973 2240 11037 2304
rect 11054 2240 11118 2304
rect 11135 2240 11199 2304
rect 11216 2240 11280 2304
rect 11297 2240 11361 2304
rect 11378 2240 11442 2304
rect 11459 2240 11523 2304
rect 11540 2240 11604 2304
rect 11621 2240 11685 2304
rect 11702 2240 11766 2304
rect 11783 2240 11847 2304
rect 11864 2240 11928 2304
rect 11945 2240 12009 2304
rect 12026 2240 12090 2304
rect 12107 2240 12171 2304
rect 12188 2240 12252 2304
rect 12269 2240 12333 2304
rect 12350 2240 12414 2304
rect 12431 2240 12495 2304
rect 12512 2240 12576 2304
rect 12593 2240 12657 2304
rect 12674 2240 12738 2304
rect 12755 2240 12819 2304
rect 12836 2240 12900 2304
rect 12917 2240 12981 2304
rect 12998 2240 13062 2304
rect 13079 2240 13143 2304
rect 13160 2240 13224 2304
rect 13241 2240 13305 2304
rect 13322 2240 13386 2304
rect 13403 2240 13467 2304
rect 13484 2240 13548 2304
rect 13565 2240 13629 2304
rect 13646 2240 13710 2304
rect 13727 2240 13791 2304
rect 13808 2240 13872 2304
rect 13889 2240 13953 2304
rect 13970 2240 14034 2304
rect 14051 2240 14115 2304
rect 14132 2240 14196 2304
rect 14213 2240 14277 2304
rect 14294 2240 14358 2304
rect 14375 2240 14439 2304
rect 14456 2240 14520 2304
rect 14537 2240 14601 2304
rect 14618 2240 14682 2304
rect 14699 2240 14763 2304
rect 14780 2240 14844 2304
rect 14861 2240 14925 2304
rect 10157 2154 10221 2218
rect 10239 2154 10303 2218
rect 10321 2154 10385 2218
rect 10403 2154 10467 2218
rect 10485 2154 10549 2218
rect 10567 2154 10631 2218
rect 10649 2154 10713 2218
rect 10730 2154 10794 2218
rect 10811 2154 10875 2218
rect 10892 2154 10956 2218
rect 10973 2154 11037 2218
rect 11054 2154 11118 2218
rect 11135 2154 11199 2218
rect 11216 2154 11280 2218
rect 11297 2154 11361 2218
rect 11378 2154 11442 2218
rect 11459 2154 11523 2218
rect 11540 2154 11604 2218
rect 11621 2154 11685 2218
rect 11702 2154 11766 2218
rect 11783 2154 11847 2218
rect 11864 2154 11928 2218
rect 11945 2154 12009 2218
rect 12026 2154 12090 2218
rect 12107 2154 12171 2218
rect 12188 2154 12252 2218
rect 12269 2154 12333 2218
rect 12350 2154 12414 2218
rect 12431 2154 12495 2218
rect 12512 2154 12576 2218
rect 12593 2154 12657 2218
rect 12674 2154 12738 2218
rect 12755 2154 12819 2218
rect 12836 2154 12900 2218
rect 12917 2154 12981 2218
rect 12998 2154 13062 2218
rect 13079 2154 13143 2218
rect 13160 2154 13224 2218
rect 13241 2154 13305 2218
rect 13322 2154 13386 2218
rect 13403 2154 13467 2218
rect 13484 2154 13548 2218
rect 13565 2154 13629 2218
rect 13646 2154 13710 2218
rect 13727 2154 13791 2218
rect 13808 2154 13872 2218
rect 13889 2154 13953 2218
rect 13970 2154 14034 2218
rect 14051 2154 14115 2218
rect 14132 2154 14196 2218
rect 14213 2154 14277 2218
rect 14294 2154 14358 2218
rect 14375 2154 14439 2218
rect 14456 2154 14520 2218
rect 14537 2154 14601 2218
rect 14618 2154 14682 2218
rect 14699 2154 14763 2218
rect 14780 2154 14844 2218
rect 14861 2154 14925 2218
rect 10157 2068 10221 2132
rect 10239 2068 10303 2132
rect 10321 2068 10385 2132
rect 10403 2068 10467 2132
rect 10485 2068 10549 2132
rect 10567 2068 10631 2132
rect 10649 2068 10713 2132
rect 10730 2068 10794 2132
rect 10811 2068 10875 2132
rect 10892 2068 10956 2132
rect 10973 2068 11037 2132
rect 11054 2068 11118 2132
rect 11135 2068 11199 2132
rect 11216 2068 11280 2132
rect 11297 2068 11361 2132
rect 11378 2068 11442 2132
rect 11459 2068 11523 2132
rect 11540 2068 11604 2132
rect 11621 2068 11685 2132
rect 11702 2068 11766 2132
rect 11783 2068 11847 2132
rect 11864 2068 11928 2132
rect 11945 2068 12009 2132
rect 12026 2068 12090 2132
rect 12107 2068 12171 2132
rect 12188 2068 12252 2132
rect 12269 2068 12333 2132
rect 12350 2068 12414 2132
rect 12431 2068 12495 2132
rect 12512 2068 12576 2132
rect 12593 2068 12657 2132
rect 12674 2068 12738 2132
rect 12755 2068 12819 2132
rect 12836 2068 12900 2132
rect 12917 2068 12981 2132
rect 12998 2068 13062 2132
rect 13079 2068 13143 2132
rect 13160 2068 13224 2132
rect 13241 2068 13305 2132
rect 13322 2068 13386 2132
rect 13403 2068 13467 2132
rect 13484 2068 13548 2132
rect 13565 2068 13629 2132
rect 13646 2068 13710 2132
rect 13727 2068 13791 2132
rect 13808 2068 13872 2132
rect 13889 2068 13953 2132
rect 13970 2068 14034 2132
rect 14051 2068 14115 2132
rect 14132 2068 14196 2132
rect 14213 2068 14277 2132
rect 14294 2068 14358 2132
rect 14375 2068 14439 2132
rect 14456 2068 14520 2132
rect 14537 2068 14601 2132
rect 14618 2068 14682 2132
rect 14699 2068 14763 2132
rect 14780 2068 14844 2132
rect 14861 2068 14925 2132
rect 10157 1982 10221 2046
rect 10239 1982 10303 2046
rect 10321 1982 10385 2046
rect 10403 1982 10467 2046
rect 10485 1982 10549 2046
rect 10567 1982 10631 2046
rect 10649 1982 10713 2046
rect 10730 1982 10794 2046
rect 10811 1982 10875 2046
rect 10892 1982 10956 2046
rect 10973 1982 11037 2046
rect 11054 1982 11118 2046
rect 11135 1982 11199 2046
rect 11216 1982 11280 2046
rect 11297 1982 11361 2046
rect 11378 1982 11442 2046
rect 11459 1982 11523 2046
rect 11540 1982 11604 2046
rect 11621 1982 11685 2046
rect 11702 1982 11766 2046
rect 11783 1982 11847 2046
rect 11864 1982 11928 2046
rect 11945 1982 12009 2046
rect 12026 1982 12090 2046
rect 12107 1982 12171 2046
rect 12188 1982 12252 2046
rect 12269 1982 12333 2046
rect 12350 1982 12414 2046
rect 12431 1982 12495 2046
rect 12512 1982 12576 2046
rect 12593 1982 12657 2046
rect 12674 1982 12738 2046
rect 12755 1982 12819 2046
rect 12836 1982 12900 2046
rect 12917 1982 12981 2046
rect 12998 1982 13062 2046
rect 13079 1982 13143 2046
rect 13160 1982 13224 2046
rect 13241 1982 13305 2046
rect 13322 1982 13386 2046
rect 13403 1982 13467 2046
rect 13484 1982 13548 2046
rect 13565 1982 13629 2046
rect 13646 1982 13710 2046
rect 13727 1982 13791 2046
rect 13808 1982 13872 2046
rect 13889 1982 13953 2046
rect 13970 1982 14034 2046
rect 14051 1982 14115 2046
rect 14132 1982 14196 2046
rect 14213 1982 14277 2046
rect 14294 1982 14358 2046
rect 14375 1982 14439 2046
rect 14456 1982 14520 2046
rect 14537 1982 14601 2046
rect 14618 1982 14682 2046
rect 14699 1982 14763 2046
rect 14780 1982 14844 2046
rect 14861 1982 14925 2046
rect 10157 1896 10221 1960
rect 10239 1896 10303 1960
rect 10321 1896 10385 1960
rect 10403 1896 10467 1960
rect 10485 1896 10549 1960
rect 10567 1896 10631 1960
rect 10649 1896 10713 1960
rect 10730 1896 10794 1960
rect 10811 1896 10875 1960
rect 10892 1896 10956 1960
rect 10973 1896 11037 1960
rect 11054 1896 11118 1960
rect 11135 1896 11199 1960
rect 11216 1896 11280 1960
rect 11297 1896 11361 1960
rect 11378 1896 11442 1960
rect 11459 1896 11523 1960
rect 11540 1896 11604 1960
rect 11621 1896 11685 1960
rect 11702 1896 11766 1960
rect 11783 1896 11847 1960
rect 11864 1896 11928 1960
rect 11945 1896 12009 1960
rect 12026 1896 12090 1960
rect 12107 1896 12171 1960
rect 12188 1896 12252 1960
rect 12269 1896 12333 1960
rect 12350 1896 12414 1960
rect 12431 1896 12495 1960
rect 12512 1896 12576 1960
rect 12593 1896 12657 1960
rect 12674 1896 12738 1960
rect 12755 1896 12819 1960
rect 12836 1896 12900 1960
rect 12917 1896 12981 1960
rect 12998 1896 13062 1960
rect 13079 1896 13143 1960
rect 13160 1896 13224 1960
rect 13241 1896 13305 1960
rect 13322 1896 13386 1960
rect 13403 1896 13467 1960
rect 13484 1896 13548 1960
rect 13565 1896 13629 1960
rect 13646 1896 13710 1960
rect 13727 1896 13791 1960
rect 13808 1896 13872 1960
rect 13889 1896 13953 1960
rect 13970 1896 14034 1960
rect 14051 1896 14115 1960
rect 14132 1896 14196 1960
rect 14213 1896 14277 1960
rect 14294 1896 14358 1960
rect 14375 1896 14439 1960
rect 14456 1896 14520 1960
rect 14537 1896 14601 1960
rect 14618 1896 14682 1960
rect 14699 1896 14763 1960
rect 14780 1896 14844 1960
rect 14861 1896 14925 1960
rect 10157 1810 10221 1874
rect 10239 1810 10303 1874
rect 10321 1810 10385 1874
rect 10403 1810 10467 1874
rect 10485 1810 10549 1874
rect 10567 1810 10631 1874
rect 10649 1810 10713 1874
rect 10730 1810 10794 1874
rect 10811 1810 10875 1874
rect 10892 1810 10956 1874
rect 10973 1810 11037 1874
rect 11054 1810 11118 1874
rect 11135 1810 11199 1874
rect 11216 1810 11280 1874
rect 11297 1810 11361 1874
rect 11378 1810 11442 1874
rect 11459 1810 11523 1874
rect 11540 1810 11604 1874
rect 11621 1810 11685 1874
rect 11702 1810 11766 1874
rect 11783 1810 11847 1874
rect 11864 1810 11928 1874
rect 11945 1810 12009 1874
rect 12026 1810 12090 1874
rect 12107 1810 12171 1874
rect 12188 1810 12252 1874
rect 12269 1810 12333 1874
rect 12350 1810 12414 1874
rect 12431 1810 12495 1874
rect 12512 1810 12576 1874
rect 12593 1810 12657 1874
rect 12674 1810 12738 1874
rect 12755 1810 12819 1874
rect 12836 1810 12900 1874
rect 12917 1810 12981 1874
rect 12998 1810 13062 1874
rect 13079 1810 13143 1874
rect 13160 1810 13224 1874
rect 13241 1810 13305 1874
rect 13322 1810 13386 1874
rect 13403 1810 13467 1874
rect 13484 1810 13548 1874
rect 13565 1810 13629 1874
rect 13646 1810 13710 1874
rect 13727 1810 13791 1874
rect 13808 1810 13872 1874
rect 13889 1810 13953 1874
rect 13970 1810 14034 1874
rect 14051 1810 14115 1874
rect 14132 1810 14196 1874
rect 14213 1810 14277 1874
rect 14294 1810 14358 1874
rect 14375 1810 14439 1874
rect 14456 1810 14520 1874
rect 14537 1810 14601 1874
rect 14618 1810 14682 1874
rect 14699 1810 14763 1874
rect 14780 1810 14844 1874
rect 14861 1810 14925 1874
rect 10157 1724 10221 1788
rect 10239 1724 10303 1788
rect 10321 1724 10385 1788
rect 10403 1724 10467 1788
rect 10485 1724 10549 1788
rect 10567 1724 10631 1788
rect 10649 1724 10713 1788
rect 10730 1724 10794 1788
rect 10811 1724 10875 1788
rect 10892 1724 10956 1788
rect 10973 1724 11037 1788
rect 11054 1724 11118 1788
rect 11135 1724 11199 1788
rect 11216 1724 11280 1788
rect 11297 1724 11361 1788
rect 11378 1724 11442 1788
rect 11459 1724 11523 1788
rect 11540 1724 11604 1788
rect 11621 1724 11685 1788
rect 11702 1724 11766 1788
rect 11783 1724 11847 1788
rect 11864 1724 11928 1788
rect 11945 1724 12009 1788
rect 12026 1724 12090 1788
rect 12107 1724 12171 1788
rect 12188 1724 12252 1788
rect 12269 1724 12333 1788
rect 12350 1724 12414 1788
rect 12431 1724 12495 1788
rect 12512 1724 12576 1788
rect 12593 1724 12657 1788
rect 12674 1724 12738 1788
rect 12755 1724 12819 1788
rect 12836 1724 12900 1788
rect 12917 1724 12981 1788
rect 12998 1724 13062 1788
rect 13079 1724 13143 1788
rect 13160 1724 13224 1788
rect 13241 1724 13305 1788
rect 13322 1724 13386 1788
rect 13403 1724 13467 1788
rect 13484 1724 13548 1788
rect 13565 1724 13629 1788
rect 13646 1724 13710 1788
rect 13727 1724 13791 1788
rect 13808 1724 13872 1788
rect 13889 1724 13953 1788
rect 13970 1724 14034 1788
rect 14051 1724 14115 1788
rect 14132 1724 14196 1788
rect 14213 1724 14277 1788
rect 14294 1724 14358 1788
rect 14375 1724 14439 1788
rect 14456 1724 14520 1788
rect 14537 1724 14601 1788
rect 14618 1724 14682 1788
rect 14699 1724 14763 1788
rect 14780 1724 14844 1788
rect 14861 1724 14925 1788
rect 10157 1638 10221 1702
rect 10239 1638 10303 1702
rect 10321 1638 10385 1702
rect 10403 1638 10467 1702
rect 10485 1638 10549 1702
rect 10567 1638 10631 1702
rect 10649 1638 10713 1702
rect 10730 1638 10794 1702
rect 10811 1638 10875 1702
rect 10892 1638 10956 1702
rect 10973 1638 11037 1702
rect 11054 1638 11118 1702
rect 11135 1638 11199 1702
rect 11216 1638 11280 1702
rect 11297 1638 11361 1702
rect 11378 1638 11442 1702
rect 11459 1638 11523 1702
rect 11540 1638 11604 1702
rect 11621 1638 11685 1702
rect 11702 1638 11766 1702
rect 11783 1638 11847 1702
rect 11864 1638 11928 1702
rect 11945 1638 12009 1702
rect 12026 1638 12090 1702
rect 12107 1638 12171 1702
rect 12188 1638 12252 1702
rect 12269 1638 12333 1702
rect 12350 1638 12414 1702
rect 12431 1638 12495 1702
rect 12512 1638 12576 1702
rect 12593 1638 12657 1702
rect 12674 1638 12738 1702
rect 12755 1638 12819 1702
rect 12836 1638 12900 1702
rect 12917 1638 12981 1702
rect 12998 1638 13062 1702
rect 13079 1638 13143 1702
rect 13160 1638 13224 1702
rect 13241 1638 13305 1702
rect 13322 1638 13386 1702
rect 13403 1638 13467 1702
rect 13484 1638 13548 1702
rect 13565 1638 13629 1702
rect 13646 1638 13710 1702
rect 13727 1638 13791 1702
rect 13808 1638 13872 1702
rect 13889 1638 13953 1702
rect 13970 1638 14034 1702
rect 14051 1638 14115 1702
rect 14132 1638 14196 1702
rect 14213 1638 14277 1702
rect 14294 1638 14358 1702
rect 14375 1638 14439 1702
rect 14456 1638 14520 1702
rect 14537 1638 14601 1702
rect 14618 1638 14682 1702
rect 14699 1638 14763 1702
rect 14780 1638 14844 1702
rect 14861 1638 14925 1702
rect 10157 1552 10221 1616
rect 10239 1552 10303 1616
rect 10321 1552 10385 1616
rect 10403 1552 10467 1616
rect 10485 1552 10549 1616
rect 10567 1552 10631 1616
rect 10649 1552 10713 1616
rect 10730 1552 10794 1616
rect 10811 1552 10875 1616
rect 10892 1552 10956 1616
rect 10973 1552 11037 1616
rect 11054 1552 11118 1616
rect 11135 1552 11199 1616
rect 11216 1552 11280 1616
rect 11297 1552 11361 1616
rect 11378 1552 11442 1616
rect 11459 1552 11523 1616
rect 11540 1552 11604 1616
rect 11621 1552 11685 1616
rect 11702 1552 11766 1616
rect 11783 1552 11847 1616
rect 11864 1552 11928 1616
rect 11945 1552 12009 1616
rect 12026 1552 12090 1616
rect 12107 1552 12171 1616
rect 12188 1552 12252 1616
rect 12269 1552 12333 1616
rect 12350 1552 12414 1616
rect 12431 1552 12495 1616
rect 12512 1552 12576 1616
rect 12593 1552 12657 1616
rect 12674 1552 12738 1616
rect 12755 1552 12819 1616
rect 12836 1552 12900 1616
rect 12917 1552 12981 1616
rect 12998 1552 13062 1616
rect 13079 1552 13143 1616
rect 13160 1552 13224 1616
rect 13241 1552 13305 1616
rect 13322 1552 13386 1616
rect 13403 1552 13467 1616
rect 13484 1552 13548 1616
rect 13565 1552 13629 1616
rect 13646 1552 13710 1616
rect 13727 1552 13791 1616
rect 13808 1552 13872 1616
rect 13889 1552 13953 1616
rect 13970 1552 14034 1616
rect 14051 1552 14115 1616
rect 14132 1552 14196 1616
rect 14213 1552 14277 1616
rect 14294 1552 14358 1616
rect 14375 1552 14439 1616
rect 14456 1552 14520 1616
rect 14537 1552 14601 1616
rect 14618 1552 14682 1616
rect 14699 1552 14763 1616
rect 14780 1552 14844 1616
rect 14861 1552 14925 1616
rect 10157 1466 10221 1530
rect 10239 1466 10303 1530
rect 10321 1466 10385 1530
rect 10403 1466 10467 1530
rect 10485 1466 10549 1530
rect 10567 1466 10631 1530
rect 10649 1466 10713 1530
rect 10730 1466 10794 1530
rect 10811 1466 10875 1530
rect 10892 1466 10956 1530
rect 10973 1466 11037 1530
rect 11054 1466 11118 1530
rect 11135 1466 11199 1530
rect 11216 1466 11280 1530
rect 11297 1466 11361 1530
rect 11378 1466 11442 1530
rect 11459 1466 11523 1530
rect 11540 1466 11604 1530
rect 11621 1466 11685 1530
rect 11702 1466 11766 1530
rect 11783 1466 11847 1530
rect 11864 1466 11928 1530
rect 11945 1466 12009 1530
rect 12026 1466 12090 1530
rect 12107 1466 12171 1530
rect 12188 1466 12252 1530
rect 12269 1466 12333 1530
rect 12350 1466 12414 1530
rect 12431 1466 12495 1530
rect 12512 1466 12576 1530
rect 12593 1466 12657 1530
rect 12674 1466 12738 1530
rect 12755 1466 12819 1530
rect 12836 1466 12900 1530
rect 12917 1466 12981 1530
rect 12998 1466 13062 1530
rect 13079 1466 13143 1530
rect 13160 1466 13224 1530
rect 13241 1466 13305 1530
rect 13322 1466 13386 1530
rect 13403 1466 13467 1530
rect 13484 1466 13548 1530
rect 13565 1466 13629 1530
rect 13646 1466 13710 1530
rect 13727 1466 13791 1530
rect 13808 1466 13872 1530
rect 13889 1466 13953 1530
rect 13970 1466 14034 1530
rect 14051 1466 14115 1530
rect 14132 1466 14196 1530
rect 14213 1466 14277 1530
rect 14294 1466 14358 1530
rect 14375 1466 14439 1530
rect 14456 1466 14520 1530
rect 14537 1466 14601 1530
rect 14618 1466 14682 1530
rect 14699 1466 14763 1530
rect 14780 1466 14844 1530
rect 14861 1466 14925 1530
rect 10157 1380 10221 1444
rect 10239 1380 10303 1444
rect 10321 1380 10385 1444
rect 10403 1380 10467 1444
rect 10485 1380 10549 1444
rect 10567 1380 10631 1444
rect 10649 1380 10713 1444
rect 10730 1380 10794 1444
rect 10811 1380 10875 1444
rect 10892 1380 10956 1444
rect 10973 1380 11037 1444
rect 11054 1380 11118 1444
rect 11135 1380 11199 1444
rect 11216 1380 11280 1444
rect 11297 1380 11361 1444
rect 11378 1380 11442 1444
rect 11459 1380 11523 1444
rect 11540 1380 11604 1444
rect 11621 1380 11685 1444
rect 11702 1380 11766 1444
rect 11783 1380 11847 1444
rect 11864 1380 11928 1444
rect 11945 1380 12009 1444
rect 12026 1380 12090 1444
rect 12107 1380 12171 1444
rect 12188 1380 12252 1444
rect 12269 1380 12333 1444
rect 12350 1380 12414 1444
rect 12431 1380 12495 1444
rect 12512 1380 12576 1444
rect 12593 1380 12657 1444
rect 12674 1380 12738 1444
rect 12755 1380 12819 1444
rect 12836 1380 12900 1444
rect 12917 1380 12981 1444
rect 12998 1380 13062 1444
rect 13079 1380 13143 1444
rect 13160 1380 13224 1444
rect 13241 1380 13305 1444
rect 13322 1380 13386 1444
rect 13403 1380 13467 1444
rect 13484 1380 13548 1444
rect 13565 1380 13629 1444
rect 13646 1380 13710 1444
rect 13727 1380 13791 1444
rect 13808 1380 13872 1444
rect 13889 1380 13953 1444
rect 13970 1380 14034 1444
rect 14051 1380 14115 1444
rect 14132 1380 14196 1444
rect 14213 1380 14277 1444
rect 14294 1380 14358 1444
rect 14375 1380 14439 1444
rect 14456 1380 14520 1444
rect 14537 1380 14601 1444
rect 14618 1380 14682 1444
rect 14699 1380 14763 1444
rect 14780 1380 14844 1444
rect 14861 1380 14925 1444
<< metal4 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18600
rect 14746 13607 15000 18600
rect 0 12417 254 13307
rect 14746 12417 15000 13307
rect 0 11247 254 12137
rect 14746 11247 15000 12137
rect 0 10881 254 10947
rect 14746 10881 15000 10947
rect 0 10225 254 10821
rect 14746 10225 15000 10821
rect 0 9929 254 10165
rect 14746 9929 15000 10165
rect 0 9273 254 9869
rect 14746 9273 15000 9869
rect 0 9147 254 9213
rect 14746 9147 15000 9213
rect 0 7917 254 8847
rect 14746 7917 15000 8847
rect 0 6947 254 7637
rect 14746 6947 15000 7637
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 254 5697
rect 14746 4767 15000 5697
rect 0 3557 254 4487
rect 14746 3557 15000 4487
rect 0 2587 193 3277
rect 14807 2587 15000 3277
rect 0 2304 4895 2307
rect 0 2240 126 2304
rect 190 2240 208 2304
rect 272 2240 290 2304
rect 354 2240 372 2304
rect 436 2240 454 2304
rect 518 2240 536 2304
rect 600 2240 618 2304
rect 682 2240 699 2304
rect 763 2240 780 2304
rect 844 2240 861 2304
rect 925 2240 942 2304
rect 1006 2240 1023 2304
rect 1087 2240 1104 2304
rect 1168 2240 1185 2304
rect 1249 2240 1266 2304
rect 1330 2240 1347 2304
rect 1411 2240 1428 2304
rect 1492 2240 1509 2304
rect 1573 2240 1590 2304
rect 1654 2240 1671 2304
rect 1735 2240 1752 2304
rect 1816 2240 1833 2304
rect 1897 2240 1914 2304
rect 1978 2240 1995 2304
rect 2059 2240 2076 2304
rect 2140 2240 2157 2304
rect 2221 2240 2238 2304
rect 2302 2240 2319 2304
rect 2383 2240 2400 2304
rect 2464 2240 2481 2304
rect 2545 2240 2562 2304
rect 2626 2240 2643 2304
rect 2707 2240 2724 2304
rect 2788 2240 2805 2304
rect 2869 2240 2886 2304
rect 2950 2240 2967 2304
rect 3031 2240 3048 2304
rect 3112 2240 3129 2304
rect 3193 2240 3210 2304
rect 3274 2240 3291 2304
rect 3355 2240 3372 2304
rect 3436 2240 3453 2304
rect 3517 2240 3534 2304
rect 3598 2240 3615 2304
rect 3679 2240 3696 2304
rect 3760 2240 3777 2304
rect 3841 2240 3858 2304
rect 3922 2240 3939 2304
rect 4003 2240 4020 2304
rect 4084 2240 4101 2304
rect 4165 2240 4182 2304
rect 4246 2240 4263 2304
rect 4327 2240 4344 2304
rect 4408 2240 4425 2304
rect 4489 2240 4506 2304
rect 4570 2240 4587 2304
rect 4651 2240 4668 2304
rect 4732 2240 4749 2304
rect 4813 2240 4830 2304
rect 4894 2240 4895 2304
rect 0 2218 4895 2240
rect 0 2154 126 2218
rect 190 2154 208 2218
rect 272 2154 290 2218
rect 354 2154 372 2218
rect 436 2154 454 2218
rect 518 2154 536 2218
rect 600 2154 618 2218
rect 682 2154 699 2218
rect 763 2154 780 2218
rect 844 2154 861 2218
rect 925 2154 942 2218
rect 1006 2154 1023 2218
rect 1087 2154 1104 2218
rect 1168 2154 1185 2218
rect 1249 2154 1266 2218
rect 1330 2154 1347 2218
rect 1411 2154 1428 2218
rect 1492 2154 1509 2218
rect 1573 2154 1590 2218
rect 1654 2154 1671 2218
rect 1735 2154 1752 2218
rect 1816 2154 1833 2218
rect 1897 2154 1914 2218
rect 1978 2154 1995 2218
rect 2059 2154 2076 2218
rect 2140 2154 2157 2218
rect 2221 2154 2238 2218
rect 2302 2154 2319 2218
rect 2383 2154 2400 2218
rect 2464 2154 2481 2218
rect 2545 2154 2562 2218
rect 2626 2154 2643 2218
rect 2707 2154 2724 2218
rect 2788 2154 2805 2218
rect 2869 2154 2886 2218
rect 2950 2154 2967 2218
rect 3031 2154 3048 2218
rect 3112 2154 3129 2218
rect 3193 2154 3210 2218
rect 3274 2154 3291 2218
rect 3355 2154 3372 2218
rect 3436 2154 3453 2218
rect 3517 2154 3534 2218
rect 3598 2154 3615 2218
rect 3679 2154 3696 2218
rect 3760 2154 3777 2218
rect 3841 2154 3858 2218
rect 3922 2154 3939 2218
rect 4003 2154 4020 2218
rect 4084 2154 4101 2218
rect 4165 2154 4182 2218
rect 4246 2154 4263 2218
rect 4327 2154 4344 2218
rect 4408 2154 4425 2218
rect 4489 2154 4506 2218
rect 4570 2154 4587 2218
rect 4651 2154 4668 2218
rect 4732 2154 4749 2218
rect 4813 2154 4830 2218
rect 4894 2154 4895 2218
rect 0 2132 4895 2154
rect 0 2068 126 2132
rect 190 2068 208 2132
rect 272 2068 290 2132
rect 354 2068 372 2132
rect 436 2068 454 2132
rect 518 2068 536 2132
rect 600 2068 618 2132
rect 682 2068 699 2132
rect 763 2068 780 2132
rect 844 2068 861 2132
rect 925 2068 942 2132
rect 1006 2068 1023 2132
rect 1087 2068 1104 2132
rect 1168 2068 1185 2132
rect 1249 2068 1266 2132
rect 1330 2068 1347 2132
rect 1411 2068 1428 2132
rect 1492 2068 1509 2132
rect 1573 2068 1590 2132
rect 1654 2068 1671 2132
rect 1735 2068 1752 2132
rect 1816 2068 1833 2132
rect 1897 2068 1914 2132
rect 1978 2068 1995 2132
rect 2059 2068 2076 2132
rect 2140 2068 2157 2132
rect 2221 2068 2238 2132
rect 2302 2068 2319 2132
rect 2383 2068 2400 2132
rect 2464 2068 2481 2132
rect 2545 2068 2562 2132
rect 2626 2068 2643 2132
rect 2707 2068 2724 2132
rect 2788 2068 2805 2132
rect 2869 2068 2886 2132
rect 2950 2068 2967 2132
rect 3031 2068 3048 2132
rect 3112 2068 3129 2132
rect 3193 2068 3210 2132
rect 3274 2068 3291 2132
rect 3355 2068 3372 2132
rect 3436 2068 3453 2132
rect 3517 2068 3534 2132
rect 3598 2068 3615 2132
rect 3679 2068 3696 2132
rect 3760 2068 3777 2132
rect 3841 2068 3858 2132
rect 3922 2068 3939 2132
rect 4003 2068 4020 2132
rect 4084 2068 4101 2132
rect 4165 2068 4182 2132
rect 4246 2068 4263 2132
rect 4327 2068 4344 2132
rect 4408 2068 4425 2132
rect 4489 2068 4506 2132
rect 4570 2068 4587 2132
rect 4651 2068 4668 2132
rect 4732 2068 4749 2132
rect 4813 2068 4830 2132
rect 4894 2068 4895 2132
rect 0 2046 4895 2068
rect 0 1982 126 2046
rect 190 1982 208 2046
rect 272 1982 290 2046
rect 354 1982 372 2046
rect 436 1982 454 2046
rect 518 1982 536 2046
rect 600 1982 618 2046
rect 682 1982 699 2046
rect 763 1982 780 2046
rect 844 1982 861 2046
rect 925 1982 942 2046
rect 1006 1982 1023 2046
rect 1087 1982 1104 2046
rect 1168 1982 1185 2046
rect 1249 1982 1266 2046
rect 1330 1982 1347 2046
rect 1411 1982 1428 2046
rect 1492 1982 1509 2046
rect 1573 1982 1590 2046
rect 1654 1982 1671 2046
rect 1735 1982 1752 2046
rect 1816 1982 1833 2046
rect 1897 1982 1914 2046
rect 1978 1982 1995 2046
rect 2059 1982 2076 2046
rect 2140 1982 2157 2046
rect 2221 1982 2238 2046
rect 2302 1982 2319 2046
rect 2383 1982 2400 2046
rect 2464 1982 2481 2046
rect 2545 1982 2562 2046
rect 2626 1982 2643 2046
rect 2707 1982 2724 2046
rect 2788 1982 2805 2046
rect 2869 1982 2886 2046
rect 2950 1982 2967 2046
rect 3031 1982 3048 2046
rect 3112 1982 3129 2046
rect 3193 1982 3210 2046
rect 3274 1982 3291 2046
rect 3355 1982 3372 2046
rect 3436 1982 3453 2046
rect 3517 1982 3534 2046
rect 3598 1982 3615 2046
rect 3679 1982 3696 2046
rect 3760 1982 3777 2046
rect 3841 1982 3858 2046
rect 3922 1982 3939 2046
rect 4003 1982 4020 2046
rect 4084 1982 4101 2046
rect 4165 1982 4182 2046
rect 4246 1982 4263 2046
rect 4327 1982 4344 2046
rect 4408 1982 4425 2046
rect 4489 1982 4506 2046
rect 4570 1982 4587 2046
rect 4651 1982 4668 2046
rect 4732 1982 4749 2046
rect 4813 1982 4830 2046
rect 4894 1982 4895 2046
rect 0 1960 4895 1982
rect 0 1896 126 1960
rect 190 1896 208 1960
rect 272 1896 290 1960
rect 354 1896 372 1960
rect 436 1896 454 1960
rect 518 1896 536 1960
rect 600 1896 618 1960
rect 682 1896 699 1960
rect 763 1896 780 1960
rect 844 1896 861 1960
rect 925 1896 942 1960
rect 1006 1896 1023 1960
rect 1087 1896 1104 1960
rect 1168 1896 1185 1960
rect 1249 1896 1266 1960
rect 1330 1896 1347 1960
rect 1411 1896 1428 1960
rect 1492 1896 1509 1960
rect 1573 1896 1590 1960
rect 1654 1896 1671 1960
rect 1735 1896 1752 1960
rect 1816 1896 1833 1960
rect 1897 1896 1914 1960
rect 1978 1896 1995 1960
rect 2059 1896 2076 1960
rect 2140 1896 2157 1960
rect 2221 1896 2238 1960
rect 2302 1896 2319 1960
rect 2383 1896 2400 1960
rect 2464 1896 2481 1960
rect 2545 1896 2562 1960
rect 2626 1896 2643 1960
rect 2707 1896 2724 1960
rect 2788 1896 2805 1960
rect 2869 1896 2886 1960
rect 2950 1896 2967 1960
rect 3031 1896 3048 1960
rect 3112 1896 3129 1960
rect 3193 1896 3210 1960
rect 3274 1896 3291 1960
rect 3355 1896 3372 1960
rect 3436 1896 3453 1960
rect 3517 1896 3534 1960
rect 3598 1896 3615 1960
rect 3679 1896 3696 1960
rect 3760 1896 3777 1960
rect 3841 1896 3858 1960
rect 3922 1896 3939 1960
rect 4003 1896 4020 1960
rect 4084 1896 4101 1960
rect 4165 1896 4182 1960
rect 4246 1896 4263 1960
rect 4327 1896 4344 1960
rect 4408 1896 4425 1960
rect 4489 1896 4506 1960
rect 4570 1896 4587 1960
rect 4651 1896 4668 1960
rect 4732 1896 4749 1960
rect 4813 1896 4830 1960
rect 4894 1896 4895 1960
rect 0 1874 4895 1896
rect 0 1810 126 1874
rect 190 1810 208 1874
rect 272 1810 290 1874
rect 354 1810 372 1874
rect 436 1810 454 1874
rect 518 1810 536 1874
rect 600 1810 618 1874
rect 682 1810 699 1874
rect 763 1810 780 1874
rect 844 1810 861 1874
rect 925 1810 942 1874
rect 1006 1810 1023 1874
rect 1087 1810 1104 1874
rect 1168 1810 1185 1874
rect 1249 1810 1266 1874
rect 1330 1810 1347 1874
rect 1411 1810 1428 1874
rect 1492 1810 1509 1874
rect 1573 1810 1590 1874
rect 1654 1810 1671 1874
rect 1735 1810 1752 1874
rect 1816 1810 1833 1874
rect 1897 1810 1914 1874
rect 1978 1810 1995 1874
rect 2059 1810 2076 1874
rect 2140 1810 2157 1874
rect 2221 1810 2238 1874
rect 2302 1810 2319 1874
rect 2383 1810 2400 1874
rect 2464 1810 2481 1874
rect 2545 1810 2562 1874
rect 2626 1810 2643 1874
rect 2707 1810 2724 1874
rect 2788 1810 2805 1874
rect 2869 1810 2886 1874
rect 2950 1810 2967 1874
rect 3031 1810 3048 1874
rect 3112 1810 3129 1874
rect 3193 1810 3210 1874
rect 3274 1810 3291 1874
rect 3355 1810 3372 1874
rect 3436 1810 3453 1874
rect 3517 1810 3534 1874
rect 3598 1810 3615 1874
rect 3679 1810 3696 1874
rect 3760 1810 3777 1874
rect 3841 1810 3858 1874
rect 3922 1810 3939 1874
rect 4003 1810 4020 1874
rect 4084 1810 4101 1874
rect 4165 1810 4182 1874
rect 4246 1810 4263 1874
rect 4327 1810 4344 1874
rect 4408 1810 4425 1874
rect 4489 1810 4506 1874
rect 4570 1810 4587 1874
rect 4651 1810 4668 1874
rect 4732 1810 4749 1874
rect 4813 1810 4830 1874
rect 4894 1810 4895 1874
rect 0 1788 4895 1810
rect 0 1724 126 1788
rect 190 1724 208 1788
rect 272 1724 290 1788
rect 354 1724 372 1788
rect 436 1724 454 1788
rect 518 1724 536 1788
rect 600 1724 618 1788
rect 682 1724 699 1788
rect 763 1724 780 1788
rect 844 1724 861 1788
rect 925 1724 942 1788
rect 1006 1724 1023 1788
rect 1087 1724 1104 1788
rect 1168 1724 1185 1788
rect 1249 1724 1266 1788
rect 1330 1724 1347 1788
rect 1411 1724 1428 1788
rect 1492 1724 1509 1788
rect 1573 1724 1590 1788
rect 1654 1724 1671 1788
rect 1735 1724 1752 1788
rect 1816 1724 1833 1788
rect 1897 1724 1914 1788
rect 1978 1724 1995 1788
rect 2059 1724 2076 1788
rect 2140 1724 2157 1788
rect 2221 1724 2238 1788
rect 2302 1724 2319 1788
rect 2383 1724 2400 1788
rect 2464 1724 2481 1788
rect 2545 1724 2562 1788
rect 2626 1724 2643 1788
rect 2707 1724 2724 1788
rect 2788 1724 2805 1788
rect 2869 1724 2886 1788
rect 2950 1724 2967 1788
rect 3031 1724 3048 1788
rect 3112 1724 3129 1788
rect 3193 1724 3210 1788
rect 3274 1724 3291 1788
rect 3355 1724 3372 1788
rect 3436 1724 3453 1788
rect 3517 1724 3534 1788
rect 3598 1724 3615 1788
rect 3679 1724 3696 1788
rect 3760 1724 3777 1788
rect 3841 1724 3858 1788
rect 3922 1724 3939 1788
rect 4003 1724 4020 1788
rect 4084 1724 4101 1788
rect 4165 1724 4182 1788
rect 4246 1724 4263 1788
rect 4327 1724 4344 1788
rect 4408 1724 4425 1788
rect 4489 1724 4506 1788
rect 4570 1724 4587 1788
rect 4651 1724 4668 1788
rect 4732 1724 4749 1788
rect 4813 1724 4830 1788
rect 4894 1724 4895 1788
rect 0 1702 4895 1724
rect 0 1638 126 1702
rect 190 1638 208 1702
rect 272 1638 290 1702
rect 354 1638 372 1702
rect 436 1638 454 1702
rect 518 1638 536 1702
rect 600 1638 618 1702
rect 682 1638 699 1702
rect 763 1638 780 1702
rect 844 1638 861 1702
rect 925 1638 942 1702
rect 1006 1638 1023 1702
rect 1087 1638 1104 1702
rect 1168 1638 1185 1702
rect 1249 1638 1266 1702
rect 1330 1638 1347 1702
rect 1411 1638 1428 1702
rect 1492 1638 1509 1702
rect 1573 1638 1590 1702
rect 1654 1638 1671 1702
rect 1735 1638 1752 1702
rect 1816 1638 1833 1702
rect 1897 1638 1914 1702
rect 1978 1638 1995 1702
rect 2059 1638 2076 1702
rect 2140 1638 2157 1702
rect 2221 1638 2238 1702
rect 2302 1638 2319 1702
rect 2383 1638 2400 1702
rect 2464 1638 2481 1702
rect 2545 1638 2562 1702
rect 2626 1638 2643 1702
rect 2707 1638 2724 1702
rect 2788 1638 2805 1702
rect 2869 1638 2886 1702
rect 2950 1638 2967 1702
rect 3031 1638 3048 1702
rect 3112 1638 3129 1702
rect 3193 1638 3210 1702
rect 3274 1638 3291 1702
rect 3355 1638 3372 1702
rect 3436 1638 3453 1702
rect 3517 1638 3534 1702
rect 3598 1638 3615 1702
rect 3679 1638 3696 1702
rect 3760 1638 3777 1702
rect 3841 1638 3858 1702
rect 3922 1638 3939 1702
rect 4003 1638 4020 1702
rect 4084 1638 4101 1702
rect 4165 1638 4182 1702
rect 4246 1638 4263 1702
rect 4327 1638 4344 1702
rect 4408 1638 4425 1702
rect 4489 1638 4506 1702
rect 4570 1638 4587 1702
rect 4651 1638 4668 1702
rect 4732 1638 4749 1702
rect 4813 1638 4830 1702
rect 4894 1638 4895 1702
rect 0 1616 4895 1638
rect 0 1552 126 1616
rect 190 1552 208 1616
rect 272 1552 290 1616
rect 354 1552 372 1616
rect 436 1552 454 1616
rect 518 1552 536 1616
rect 600 1552 618 1616
rect 682 1552 699 1616
rect 763 1552 780 1616
rect 844 1552 861 1616
rect 925 1552 942 1616
rect 1006 1552 1023 1616
rect 1087 1552 1104 1616
rect 1168 1552 1185 1616
rect 1249 1552 1266 1616
rect 1330 1552 1347 1616
rect 1411 1552 1428 1616
rect 1492 1552 1509 1616
rect 1573 1552 1590 1616
rect 1654 1552 1671 1616
rect 1735 1552 1752 1616
rect 1816 1552 1833 1616
rect 1897 1552 1914 1616
rect 1978 1552 1995 1616
rect 2059 1552 2076 1616
rect 2140 1552 2157 1616
rect 2221 1552 2238 1616
rect 2302 1552 2319 1616
rect 2383 1552 2400 1616
rect 2464 1552 2481 1616
rect 2545 1552 2562 1616
rect 2626 1552 2643 1616
rect 2707 1552 2724 1616
rect 2788 1552 2805 1616
rect 2869 1552 2886 1616
rect 2950 1552 2967 1616
rect 3031 1552 3048 1616
rect 3112 1552 3129 1616
rect 3193 1552 3210 1616
rect 3274 1552 3291 1616
rect 3355 1552 3372 1616
rect 3436 1552 3453 1616
rect 3517 1552 3534 1616
rect 3598 1552 3615 1616
rect 3679 1552 3696 1616
rect 3760 1552 3777 1616
rect 3841 1552 3858 1616
rect 3922 1552 3939 1616
rect 4003 1552 4020 1616
rect 4084 1552 4101 1616
rect 4165 1552 4182 1616
rect 4246 1552 4263 1616
rect 4327 1552 4344 1616
rect 4408 1552 4425 1616
rect 4489 1552 4506 1616
rect 4570 1552 4587 1616
rect 4651 1552 4668 1616
rect 4732 1552 4749 1616
rect 4813 1552 4830 1616
rect 4894 1552 4895 1616
rect 0 1530 4895 1552
rect 0 1466 126 1530
rect 190 1466 208 1530
rect 272 1466 290 1530
rect 354 1466 372 1530
rect 436 1466 454 1530
rect 518 1466 536 1530
rect 600 1466 618 1530
rect 682 1466 699 1530
rect 763 1466 780 1530
rect 844 1466 861 1530
rect 925 1466 942 1530
rect 1006 1466 1023 1530
rect 1087 1466 1104 1530
rect 1168 1466 1185 1530
rect 1249 1466 1266 1530
rect 1330 1466 1347 1530
rect 1411 1466 1428 1530
rect 1492 1466 1509 1530
rect 1573 1466 1590 1530
rect 1654 1466 1671 1530
rect 1735 1466 1752 1530
rect 1816 1466 1833 1530
rect 1897 1466 1914 1530
rect 1978 1466 1995 1530
rect 2059 1466 2076 1530
rect 2140 1466 2157 1530
rect 2221 1466 2238 1530
rect 2302 1466 2319 1530
rect 2383 1466 2400 1530
rect 2464 1466 2481 1530
rect 2545 1466 2562 1530
rect 2626 1466 2643 1530
rect 2707 1466 2724 1530
rect 2788 1466 2805 1530
rect 2869 1466 2886 1530
rect 2950 1466 2967 1530
rect 3031 1466 3048 1530
rect 3112 1466 3129 1530
rect 3193 1466 3210 1530
rect 3274 1466 3291 1530
rect 3355 1466 3372 1530
rect 3436 1466 3453 1530
rect 3517 1466 3534 1530
rect 3598 1466 3615 1530
rect 3679 1466 3696 1530
rect 3760 1466 3777 1530
rect 3841 1466 3858 1530
rect 3922 1466 3939 1530
rect 4003 1466 4020 1530
rect 4084 1466 4101 1530
rect 4165 1466 4182 1530
rect 4246 1466 4263 1530
rect 4327 1466 4344 1530
rect 4408 1466 4425 1530
rect 4489 1466 4506 1530
rect 4570 1466 4587 1530
rect 4651 1466 4668 1530
rect 4732 1466 4749 1530
rect 4813 1466 4830 1530
rect 4894 1466 4895 1530
rect 0 1444 4895 1466
rect 0 1380 126 1444
rect 190 1380 208 1444
rect 272 1380 290 1444
rect 354 1380 372 1444
rect 436 1380 454 1444
rect 518 1380 536 1444
rect 600 1380 618 1444
rect 682 1380 699 1444
rect 763 1380 780 1444
rect 844 1380 861 1444
rect 925 1380 942 1444
rect 1006 1380 1023 1444
rect 1087 1380 1104 1444
rect 1168 1380 1185 1444
rect 1249 1380 1266 1444
rect 1330 1380 1347 1444
rect 1411 1380 1428 1444
rect 1492 1380 1509 1444
rect 1573 1380 1590 1444
rect 1654 1380 1671 1444
rect 1735 1380 1752 1444
rect 1816 1380 1833 1444
rect 1897 1380 1914 1444
rect 1978 1380 1995 1444
rect 2059 1380 2076 1444
rect 2140 1380 2157 1444
rect 2221 1380 2238 1444
rect 2302 1380 2319 1444
rect 2383 1380 2400 1444
rect 2464 1380 2481 1444
rect 2545 1380 2562 1444
rect 2626 1380 2643 1444
rect 2707 1380 2724 1444
rect 2788 1380 2805 1444
rect 2869 1380 2886 1444
rect 2950 1380 2967 1444
rect 3031 1380 3048 1444
rect 3112 1380 3129 1444
rect 3193 1380 3210 1444
rect 3274 1380 3291 1444
rect 3355 1380 3372 1444
rect 3436 1380 3453 1444
rect 3517 1380 3534 1444
rect 3598 1380 3615 1444
rect 3679 1380 3696 1444
rect 3760 1380 3777 1444
rect 3841 1380 3858 1444
rect 3922 1380 3939 1444
rect 4003 1380 4020 1444
rect 4084 1380 4101 1444
rect 4165 1380 4182 1444
rect 4246 1380 4263 1444
rect 4327 1380 4344 1444
rect 4408 1380 4425 1444
rect 4489 1380 4506 1444
rect 4570 1380 4587 1444
rect 4651 1380 4668 1444
rect 4732 1380 4749 1444
rect 4813 1380 4830 1444
rect 4894 1380 4895 1444
rect 0 1377 4895 1380
rect 10156 2304 15000 2307
rect 10156 2240 10157 2304
rect 10221 2240 10239 2304
rect 10303 2240 10321 2304
rect 10385 2240 10403 2304
rect 10467 2240 10485 2304
rect 10549 2240 10567 2304
rect 10631 2240 10649 2304
rect 10713 2240 10730 2304
rect 10794 2240 10811 2304
rect 10875 2240 10892 2304
rect 10956 2240 10973 2304
rect 11037 2240 11054 2304
rect 11118 2240 11135 2304
rect 11199 2240 11216 2304
rect 11280 2240 11297 2304
rect 11361 2240 11378 2304
rect 11442 2240 11459 2304
rect 11523 2240 11540 2304
rect 11604 2240 11621 2304
rect 11685 2240 11702 2304
rect 11766 2240 11783 2304
rect 11847 2240 11864 2304
rect 11928 2240 11945 2304
rect 12009 2240 12026 2304
rect 12090 2240 12107 2304
rect 12171 2240 12188 2304
rect 12252 2240 12269 2304
rect 12333 2240 12350 2304
rect 12414 2240 12431 2304
rect 12495 2240 12512 2304
rect 12576 2240 12593 2304
rect 12657 2240 12674 2304
rect 12738 2240 12755 2304
rect 12819 2240 12836 2304
rect 12900 2240 12917 2304
rect 12981 2240 12998 2304
rect 13062 2240 13079 2304
rect 13143 2240 13160 2304
rect 13224 2240 13241 2304
rect 13305 2240 13322 2304
rect 13386 2240 13403 2304
rect 13467 2240 13484 2304
rect 13548 2240 13565 2304
rect 13629 2240 13646 2304
rect 13710 2240 13727 2304
rect 13791 2240 13808 2304
rect 13872 2240 13889 2304
rect 13953 2240 13970 2304
rect 14034 2240 14051 2304
rect 14115 2240 14132 2304
rect 14196 2240 14213 2304
rect 14277 2240 14294 2304
rect 14358 2240 14375 2304
rect 14439 2240 14456 2304
rect 14520 2240 14537 2304
rect 14601 2240 14618 2304
rect 14682 2240 14699 2304
rect 14763 2240 14780 2304
rect 14844 2240 14861 2304
rect 14925 2240 15000 2304
rect 10156 2218 15000 2240
rect 10156 2154 10157 2218
rect 10221 2154 10239 2218
rect 10303 2154 10321 2218
rect 10385 2154 10403 2218
rect 10467 2154 10485 2218
rect 10549 2154 10567 2218
rect 10631 2154 10649 2218
rect 10713 2154 10730 2218
rect 10794 2154 10811 2218
rect 10875 2154 10892 2218
rect 10956 2154 10973 2218
rect 11037 2154 11054 2218
rect 11118 2154 11135 2218
rect 11199 2154 11216 2218
rect 11280 2154 11297 2218
rect 11361 2154 11378 2218
rect 11442 2154 11459 2218
rect 11523 2154 11540 2218
rect 11604 2154 11621 2218
rect 11685 2154 11702 2218
rect 11766 2154 11783 2218
rect 11847 2154 11864 2218
rect 11928 2154 11945 2218
rect 12009 2154 12026 2218
rect 12090 2154 12107 2218
rect 12171 2154 12188 2218
rect 12252 2154 12269 2218
rect 12333 2154 12350 2218
rect 12414 2154 12431 2218
rect 12495 2154 12512 2218
rect 12576 2154 12593 2218
rect 12657 2154 12674 2218
rect 12738 2154 12755 2218
rect 12819 2154 12836 2218
rect 12900 2154 12917 2218
rect 12981 2154 12998 2218
rect 13062 2154 13079 2218
rect 13143 2154 13160 2218
rect 13224 2154 13241 2218
rect 13305 2154 13322 2218
rect 13386 2154 13403 2218
rect 13467 2154 13484 2218
rect 13548 2154 13565 2218
rect 13629 2154 13646 2218
rect 13710 2154 13727 2218
rect 13791 2154 13808 2218
rect 13872 2154 13889 2218
rect 13953 2154 13970 2218
rect 14034 2154 14051 2218
rect 14115 2154 14132 2218
rect 14196 2154 14213 2218
rect 14277 2154 14294 2218
rect 14358 2154 14375 2218
rect 14439 2154 14456 2218
rect 14520 2154 14537 2218
rect 14601 2154 14618 2218
rect 14682 2154 14699 2218
rect 14763 2154 14780 2218
rect 14844 2154 14861 2218
rect 14925 2154 15000 2218
rect 10156 2132 15000 2154
rect 10156 2068 10157 2132
rect 10221 2068 10239 2132
rect 10303 2068 10321 2132
rect 10385 2068 10403 2132
rect 10467 2068 10485 2132
rect 10549 2068 10567 2132
rect 10631 2068 10649 2132
rect 10713 2068 10730 2132
rect 10794 2068 10811 2132
rect 10875 2068 10892 2132
rect 10956 2068 10973 2132
rect 11037 2068 11054 2132
rect 11118 2068 11135 2132
rect 11199 2068 11216 2132
rect 11280 2068 11297 2132
rect 11361 2068 11378 2132
rect 11442 2068 11459 2132
rect 11523 2068 11540 2132
rect 11604 2068 11621 2132
rect 11685 2068 11702 2132
rect 11766 2068 11783 2132
rect 11847 2068 11864 2132
rect 11928 2068 11945 2132
rect 12009 2068 12026 2132
rect 12090 2068 12107 2132
rect 12171 2068 12188 2132
rect 12252 2068 12269 2132
rect 12333 2068 12350 2132
rect 12414 2068 12431 2132
rect 12495 2068 12512 2132
rect 12576 2068 12593 2132
rect 12657 2068 12674 2132
rect 12738 2068 12755 2132
rect 12819 2068 12836 2132
rect 12900 2068 12917 2132
rect 12981 2068 12998 2132
rect 13062 2068 13079 2132
rect 13143 2068 13160 2132
rect 13224 2068 13241 2132
rect 13305 2068 13322 2132
rect 13386 2068 13403 2132
rect 13467 2068 13484 2132
rect 13548 2068 13565 2132
rect 13629 2068 13646 2132
rect 13710 2068 13727 2132
rect 13791 2068 13808 2132
rect 13872 2068 13889 2132
rect 13953 2068 13970 2132
rect 14034 2068 14051 2132
rect 14115 2068 14132 2132
rect 14196 2068 14213 2132
rect 14277 2068 14294 2132
rect 14358 2068 14375 2132
rect 14439 2068 14456 2132
rect 14520 2068 14537 2132
rect 14601 2068 14618 2132
rect 14682 2068 14699 2132
rect 14763 2068 14780 2132
rect 14844 2068 14861 2132
rect 14925 2068 15000 2132
rect 10156 2046 15000 2068
rect 10156 1982 10157 2046
rect 10221 1982 10239 2046
rect 10303 1982 10321 2046
rect 10385 1982 10403 2046
rect 10467 1982 10485 2046
rect 10549 1982 10567 2046
rect 10631 1982 10649 2046
rect 10713 1982 10730 2046
rect 10794 1982 10811 2046
rect 10875 1982 10892 2046
rect 10956 1982 10973 2046
rect 11037 1982 11054 2046
rect 11118 1982 11135 2046
rect 11199 1982 11216 2046
rect 11280 1982 11297 2046
rect 11361 1982 11378 2046
rect 11442 1982 11459 2046
rect 11523 1982 11540 2046
rect 11604 1982 11621 2046
rect 11685 1982 11702 2046
rect 11766 1982 11783 2046
rect 11847 1982 11864 2046
rect 11928 1982 11945 2046
rect 12009 1982 12026 2046
rect 12090 1982 12107 2046
rect 12171 1982 12188 2046
rect 12252 1982 12269 2046
rect 12333 1982 12350 2046
rect 12414 1982 12431 2046
rect 12495 1982 12512 2046
rect 12576 1982 12593 2046
rect 12657 1982 12674 2046
rect 12738 1982 12755 2046
rect 12819 1982 12836 2046
rect 12900 1982 12917 2046
rect 12981 1982 12998 2046
rect 13062 1982 13079 2046
rect 13143 1982 13160 2046
rect 13224 1982 13241 2046
rect 13305 1982 13322 2046
rect 13386 1982 13403 2046
rect 13467 1982 13484 2046
rect 13548 1982 13565 2046
rect 13629 1982 13646 2046
rect 13710 1982 13727 2046
rect 13791 1982 13808 2046
rect 13872 1982 13889 2046
rect 13953 1982 13970 2046
rect 14034 1982 14051 2046
rect 14115 1982 14132 2046
rect 14196 1982 14213 2046
rect 14277 1982 14294 2046
rect 14358 1982 14375 2046
rect 14439 1982 14456 2046
rect 14520 1982 14537 2046
rect 14601 1982 14618 2046
rect 14682 1982 14699 2046
rect 14763 1982 14780 2046
rect 14844 1982 14861 2046
rect 14925 1982 15000 2046
rect 10156 1960 15000 1982
rect 10156 1896 10157 1960
rect 10221 1896 10239 1960
rect 10303 1896 10321 1960
rect 10385 1896 10403 1960
rect 10467 1896 10485 1960
rect 10549 1896 10567 1960
rect 10631 1896 10649 1960
rect 10713 1896 10730 1960
rect 10794 1896 10811 1960
rect 10875 1896 10892 1960
rect 10956 1896 10973 1960
rect 11037 1896 11054 1960
rect 11118 1896 11135 1960
rect 11199 1896 11216 1960
rect 11280 1896 11297 1960
rect 11361 1896 11378 1960
rect 11442 1896 11459 1960
rect 11523 1896 11540 1960
rect 11604 1896 11621 1960
rect 11685 1896 11702 1960
rect 11766 1896 11783 1960
rect 11847 1896 11864 1960
rect 11928 1896 11945 1960
rect 12009 1896 12026 1960
rect 12090 1896 12107 1960
rect 12171 1896 12188 1960
rect 12252 1896 12269 1960
rect 12333 1896 12350 1960
rect 12414 1896 12431 1960
rect 12495 1896 12512 1960
rect 12576 1896 12593 1960
rect 12657 1896 12674 1960
rect 12738 1896 12755 1960
rect 12819 1896 12836 1960
rect 12900 1896 12917 1960
rect 12981 1896 12998 1960
rect 13062 1896 13079 1960
rect 13143 1896 13160 1960
rect 13224 1896 13241 1960
rect 13305 1896 13322 1960
rect 13386 1896 13403 1960
rect 13467 1896 13484 1960
rect 13548 1896 13565 1960
rect 13629 1896 13646 1960
rect 13710 1896 13727 1960
rect 13791 1896 13808 1960
rect 13872 1896 13889 1960
rect 13953 1896 13970 1960
rect 14034 1896 14051 1960
rect 14115 1896 14132 1960
rect 14196 1896 14213 1960
rect 14277 1896 14294 1960
rect 14358 1896 14375 1960
rect 14439 1896 14456 1960
rect 14520 1896 14537 1960
rect 14601 1896 14618 1960
rect 14682 1896 14699 1960
rect 14763 1896 14780 1960
rect 14844 1896 14861 1960
rect 14925 1896 15000 1960
rect 10156 1874 15000 1896
rect 10156 1810 10157 1874
rect 10221 1810 10239 1874
rect 10303 1810 10321 1874
rect 10385 1810 10403 1874
rect 10467 1810 10485 1874
rect 10549 1810 10567 1874
rect 10631 1810 10649 1874
rect 10713 1810 10730 1874
rect 10794 1810 10811 1874
rect 10875 1810 10892 1874
rect 10956 1810 10973 1874
rect 11037 1810 11054 1874
rect 11118 1810 11135 1874
rect 11199 1810 11216 1874
rect 11280 1810 11297 1874
rect 11361 1810 11378 1874
rect 11442 1810 11459 1874
rect 11523 1810 11540 1874
rect 11604 1810 11621 1874
rect 11685 1810 11702 1874
rect 11766 1810 11783 1874
rect 11847 1810 11864 1874
rect 11928 1810 11945 1874
rect 12009 1810 12026 1874
rect 12090 1810 12107 1874
rect 12171 1810 12188 1874
rect 12252 1810 12269 1874
rect 12333 1810 12350 1874
rect 12414 1810 12431 1874
rect 12495 1810 12512 1874
rect 12576 1810 12593 1874
rect 12657 1810 12674 1874
rect 12738 1810 12755 1874
rect 12819 1810 12836 1874
rect 12900 1810 12917 1874
rect 12981 1810 12998 1874
rect 13062 1810 13079 1874
rect 13143 1810 13160 1874
rect 13224 1810 13241 1874
rect 13305 1810 13322 1874
rect 13386 1810 13403 1874
rect 13467 1810 13484 1874
rect 13548 1810 13565 1874
rect 13629 1810 13646 1874
rect 13710 1810 13727 1874
rect 13791 1810 13808 1874
rect 13872 1810 13889 1874
rect 13953 1810 13970 1874
rect 14034 1810 14051 1874
rect 14115 1810 14132 1874
rect 14196 1810 14213 1874
rect 14277 1810 14294 1874
rect 14358 1810 14375 1874
rect 14439 1810 14456 1874
rect 14520 1810 14537 1874
rect 14601 1810 14618 1874
rect 14682 1810 14699 1874
rect 14763 1810 14780 1874
rect 14844 1810 14861 1874
rect 14925 1810 15000 1874
rect 10156 1788 15000 1810
rect 10156 1724 10157 1788
rect 10221 1724 10239 1788
rect 10303 1724 10321 1788
rect 10385 1724 10403 1788
rect 10467 1724 10485 1788
rect 10549 1724 10567 1788
rect 10631 1724 10649 1788
rect 10713 1724 10730 1788
rect 10794 1724 10811 1788
rect 10875 1724 10892 1788
rect 10956 1724 10973 1788
rect 11037 1724 11054 1788
rect 11118 1724 11135 1788
rect 11199 1724 11216 1788
rect 11280 1724 11297 1788
rect 11361 1724 11378 1788
rect 11442 1724 11459 1788
rect 11523 1724 11540 1788
rect 11604 1724 11621 1788
rect 11685 1724 11702 1788
rect 11766 1724 11783 1788
rect 11847 1724 11864 1788
rect 11928 1724 11945 1788
rect 12009 1724 12026 1788
rect 12090 1724 12107 1788
rect 12171 1724 12188 1788
rect 12252 1724 12269 1788
rect 12333 1724 12350 1788
rect 12414 1724 12431 1788
rect 12495 1724 12512 1788
rect 12576 1724 12593 1788
rect 12657 1724 12674 1788
rect 12738 1724 12755 1788
rect 12819 1724 12836 1788
rect 12900 1724 12917 1788
rect 12981 1724 12998 1788
rect 13062 1724 13079 1788
rect 13143 1724 13160 1788
rect 13224 1724 13241 1788
rect 13305 1724 13322 1788
rect 13386 1724 13403 1788
rect 13467 1724 13484 1788
rect 13548 1724 13565 1788
rect 13629 1724 13646 1788
rect 13710 1724 13727 1788
rect 13791 1724 13808 1788
rect 13872 1724 13889 1788
rect 13953 1724 13970 1788
rect 14034 1724 14051 1788
rect 14115 1724 14132 1788
rect 14196 1724 14213 1788
rect 14277 1724 14294 1788
rect 14358 1724 14375 1788
rect 14439 1724 14456 1788
rect 14520 1724 14537 1788
rect 14601 1724 14618 1788
rect 14682 1724 14699 1788
rect 14763 1724 14780 1788
rect 14844 1724 14861 1788
rect 14925 1724 15000 1788
rect 10156 1702 15000 1724
rect 10156 1638 10157 1702
rect 10221 1638 10239 1702
rect 10303 1638 10321 1702
rect 10385 1638 10403 1702
rect 10467 1638 10485 1702
rect 10549 1638 10567 1702
rect 10631 1638 10649 1702
rect 10713 1638 10730 1702
rect 10794 1638 10811 1702
rect 10875 1638 10892 1702
rect 10956 1638 10973 1702
rect 11037 1638 11054 1702
rect 11118 1638 11135 1702
rect 11199 1638 11216 1702
rect 11280 1638 11297 1702
rect 11361 1638 11378 1702
rect 11442 1638 11459 1702
rect 11523 1638 11540 1702
rect 11604 1638 11621 1702
rect 11685 1638 11702 1702
rect 11766 1638 11783 1702
rect 11847 1638 11864 1702
rect 11928 1638 11945 1702
rect 12009 1638 12026 1702
rect 12090 1638 12107 1702
rect 12171 1638 12188 1702
rect 12252 1638 12269 1702
rect 12333 1638 12350 1702
rect 12414 1638 12431 1702
rect 12495 1638 12512 1702
rect 12576 1638 12593 1702
rect 12657 1638 12674 1702
rect 12738 1638 12755 1702
rect 12819 1638 12836 1702
rect 12900 1638 12917 1702
rect 12981 1638 12998 1702
rect 13062 1638 13079 1702
rect 13143 1638 13160 1702
rect 13224 1638 13241 1702
rect 13305 1638 13322 1702
rect 13386 1638 13403 1702
rect 13467 1638 13484 1702
rect 13548 1638 13565 1702
rect 13629 1638 13646 1702
rect 13710 1638 13727 1702
rect 13791 1638 13808 1702
rect 13872 1638 13889 1702
rect 13953 1638 13970 1702
rect 14034 1638 14051 1702
rect 14115 1638 14132 1702
rect 14196 1638 14213 1702
rect 14277 1638 14294 1702
rect 14358 1638 14375 1702
rect 14439 1638 14456 1702
rect 14520 1638 14537 1702
rect 14601 1638 14618 1702
rect 14682 1638 14699 1702
rect 14763 1638 14780 1702
rect 14844 1638 14861 1702
rect 14925 1638 15000 1702
rect 10156 1616 15000 1638
rect 10156 1552 10157 1616
rect 10221 1552 10239 1616
rect 10303 1552 10321 1616
rect 10385 1552 10403 1616
rect 10467 1552 10485 1616
rect 10549 1552 10567 1616
rect 10631 1552 10649 1616
rect 10713 1552 10730 1616
rect 10794 1552 10811 1616
rect 10875 1552 10892 1616
rect 10956 1552 10973 1616
rect 11037 1552 11054 1616
rect 11118 1552 11135 1616
rect 11199 1552 11216 1616
rect 11280 1552 11297 1616
rect 11361 1552 11378 1616
rect 11442 1552 11459 1616
rect 11523 1552 11540 1616
rect 11604 1552 11621 1616
rect 11685 1552 11702 1616
rect 11766 1552 11783 1616
rect 11847 1552 11864 1616
rect 11928 1552 11945 1616
rect 12009 1552 12026 1616
rect 12090 1552 12107 1616
rect 12171 1552 12188 1616
rect 12252 1552 12269 1616
rect 12333 1552 12350 1616
rect 12414 1552 12431 1616
rect 12495 1552 12512 1616
rect 12576 1552 12593 1616
rect 12657 1552 12674 1616
rect 12738 1552 12755 1616
rect 12819 1552 12836 1616
rect 12900 1552 12917 1616
rect 12981 1552 12998 1616
rect 13062 1552 13079 1616
rect 13143 1552 13160 1616
rect 13224 1552 13241 1616
rect 13305 1552 13322 1616
rect 13386 1552 13403 1616
rect 13467 1552 13484 1616
rect 13548 1552 13565 1616
rect 13629 1552 13646 1616
rect 13710 1552 13727 1616
rect 13791 1552 13808 1616
rect 13872 1552 13889 1616
rect 13953 1552 13970 1616
rect 14034 1552 14051 1616
rect 14115 1552 14132 1616
rect 14196 1552 14213 1616
rect 14277 1552 14294 1616
rect 14358 1552 14375 1616
rect 14439 1552 14456 1616
rect 14520 1552 14537 1616
rect 14601 1552 14618 1616
rect 14682 1552 14699 1616
rect 14763 1552 14780 1616
rect 14844 1552 14861 1616
rect 14925 1552 15000 1616
rect 10156 1530 15000 1552
rect 10156 1466 10157 1530
rect 10221 1466 10239 1530
rect 10303 1466 10321 1530
rect 10385 1466 10403 1530
rect 10467 1466 10485 1530
rect 10549 1466 10567 1530
rect 10631 1466 10649 1530
rect 10713 1466 10730 1530
rect 10794 1466 10811 1530
rect 10875 1466 10892 1530
rect 10956 1466 10973 1530
rect 11037 1466 11054 1530
rect 11118 1466 11135 1530
rect 11199 1466 11216 1530
rect 11280 1466 11297 1530
rect 11361 1466 11378 1530
rect 11442 1466 11459 1530
rect 11523 1466 11540 1530
rect 11604 1466 11621 1530
rect 11685 1466 11702 1530
rect 11766 1466 11783 1530
rect 11847 1466 11864 1530
rect 11928 1466 11945 1530
rect 12009 1466 12026 1530
rect 12090 1466 12107 1530
rect 12171 1466 12188 1530
rect 12252 1466 12269 1530
rect 12333 1466 12350 1530
rect 12414 1466 12431 1530
rect 12495 1466 12512 1530
rect 12576 1466 12593 1530
rect 12657 1466 12674 1530
rect 12738 1466 12755 1530
rect 12819 1466 12836 1530
rect 12900 1466 12917 1530
rect 12981 1466 12998 1530
rect 13062 1466 13079 1530
rect 13143 1466 13160 1530
rect 13224 1466 13241 1530
rect 13305 1466 13322 1530
rect 13386 1466 13403 1530
rect 13467 1466 13484 1530
rect 13548 1466 13565 1530
rect 13629 1466 13646 1530
rect 13710 1466 13727 1530
rect 13791 1466 13808 1530
rect 13872 1466 13889 1530
rect 13953 1466 13970 1530
rect 14034 1466 14051 1530
rect 14115 1466 14132 1530
rect 14196 1466 14213 1530
rect 14277 1466 14294 1530
rect 14358 1466 14375 1530
rect 14439 1466 14456 1530
rect 14520 1466 14537 1530
rect 14601 1466 14618 1530
rect 14682 1466 14699 1530
rect 14763 1466 14780 1530
rect 14844 1466 14861 1530
rect 14925 1466 15000 1530
rect 10156 1444 15000 1466
rect 10156 1380 10157 1444
rect 10221 1380 10239 1444
rect 10303 1380 10321 1444
rect 10385 1380 10403 1444
rect 10467 1380 10485 1444
rect 10549 1380 10567 1444
rect 10631 1380 10649 1444
rect 10713 1380 10730 1444
rect 10794 1380 10811 1444
rect 10875 1380 10892 1444
rect 10956 1380 10973 1444
rect 11037 1380 11054 1444
rect 11118 1380 11135 1444
rect 11199 1380 11216 1444
rect 11280 1380 11297 1444
rect 11361 1380 11378 1444
rect 11442 1380 11459 1444
rect 11523 1380 11540 1444
rect 11604 1380 11621 1444
rect 11685 1380 11702 1444
rect 11766 1380 11783 1444
rect 11847 1380 11864 1444
rect 11928 1380 11945 1444
rect 12009 1380 12026 1444
rect 12090 1380 12107 1444
rect 12171 1380 12188 1444
rect 12252 1380 12269 1444
rect 12333 1380 12350 1444
rect 12414 1380 12431 1444
rect 12495 1380 12512 1444
rect 12576 1380 12593 1444
rect 12657 1380 12674 1444
rect 12738 1380 12755 1444
rect 12819 1380 12836 1444
rect 12900 1380 12917 1444
rect 12981 1380 12998 1444
rect 13062 1380 13079 1444
rect 13143 1380 13160 1444
rect 13224 1380 13241 1444
rect 13305 1380 13322 1444
rect 13386 1380 13403 1444
rect 13467 1380 13484 1444
rect 13548 1380 13565 1444
rect 13629 1380 13646 1444
rect 13710 1380 13727 1444
rect 13791 1380 13808 1444
rect 13872 1380 13889 1444
rect 13953 1380 13970 1444
rect 14034 1380 14051 1444
rect 14115 1380 14132 1444
rect 14196 1380 14213 1444
rect 14277 1380 14294 1444
rect 14358 1380 14375 1444
rect 14439 1380 14456 1444
rect 14520 1380 14537 1444
rect 14601 1380 14618 1444
rect 14682 1380 14699 1444
rect 14763 1380 14780 1444
rect 14844 1380 14861 1444
rect 14925 1380 15000 1444
rect 10156 1377 15000 1380
rect 0 7 254 1097
rect 14746 7 15000 1097
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18597
rect 14746 13607 15000 18597
rect 0 12437 254 13287
rect 14746 12437 15000 13287
rect 0 11267 254 12117
rect 14746 11267 15000 12117
rect 0 9147 254 10947
rect 14746 9147 15000 10947
rect 0 7937 254 8827
rect 14746 7937 15000 8827
rect 0 6968 254 7617
rect 14746 6968 15000 7617
rect 0 5997 254 6647
rect 14746 5997 15000 6647
rect 0 4787 254 5677
rect 14746 4787 15000 5677
rect 0 3577 254 4467
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 14746 1397 15000 2287
rect 0 27 254 1077
rect 14746 27 15000 1077
use sky130_fd_io__com_bus_hookup  sky130_fd_io__com_bus_hookup_0
timestamp 1640697850
transform 1 0 0 0 1 149
box 0 -142 15000 39451
<< labels >>
flabel metal5 s 0 12437 254 13287 3 FreeSans 520 0 0 0 VDDIO_Q
port 1 nsew power bidirectional
flabel metal5 s 0 13607 254 18597 3 FreeSans 520 0 0 0 VDDIO
port 2 nsew power bidirectional
flabel metal5 s 0 9147 254 10947 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 14746 27 15000 1077 3 FreeSans 520 180 0 0 VCCHIB
port 4 nsew power bidirectional
flabel metal5 s 14746 1397 15000 2287 3 FreeSans 520 180 0 0 VCCD
port 5 nsew power bidirectional
flabel metal5 s 14807 2607 15000 3257 3 FreeSans 520 180 0 0 VDDA
port 6 nsew power bidirectional
flabel metal5 s 14746 3577 15000 4467 3 FreeSans 520 180 0 0 VDDIO
port 2 nsew power bidirectional
flabel metal5 s 14746 11267 15000 12117 3 FreeSans 520 180 0 0 VSSIO_Q
port 7 nsew ground bidirectional
flabel metal5 s 14746 5997 15000 6647 3 FreeSans 520 180 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal5 s 14746 4787 15000 5677 3 FreeSans 520 180 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal5 s 14746 7937 15000 8827 3 FreeSans 520 180 0 0 VSSD
port 10 nsew ground bidirectional
flabel metal5 s 14746 6968 15000 7617 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 14746 12437 15000 13287 3 FreeSans 520 180 0 0 VDDIO_Q
port 1 nsew power bidirectional
flabel metal5 s 14746 13607 15000 18597 3 FreeSans 520 180 0 0 VDDIO
port 2 nsew power bidirectional
flabel metal5 s 14746 9147 15000 10947 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal5 s 14746 34757 15000 39600 3 FreeSans 520 180 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal5 s 0 34757 254 39600 3 FreeSans 520 0 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal5 s 0 27 254 1077 3 FreeSans 520 0 0 0 VCCHIB
port 4 nsew power bidirectional
flabel metal5 s 0 1397 254 2287 3 FreeSans 520 0 0 0 VCCD
port 5 nsew power bidirectional
flabel metal5 s 0 2607 193 3257 3 FreeSans 520 0 0 0 VDDA
port 6 nsew power bidirectional
flabel metal5 s 0 3577 254 4467 3 FreeSans 520 0 0 0 VDDIO
port 2 nsew power bidirectional
flabel metal5 s 0 11267 254 12117 3 FreeSans 520 0 0 0 VSSIO_Q
port 7 nsew ground bidirectional
flabel metal5 s 0 5997 254 6647 3 FreeSans 520 0 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal5 s 0 4787 254 5677 3 FreeSans 520 0 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal5 s 0 7937 254 8827 3 FreeSans 520 0 0 0 VSSD
port 10 nsew ground bidirectional
flabel metal5 s 0 6968 254 7617 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 14746 7 15000 1097 3 FreeSans 520 180 0 0 VCCHIB
port 4 nsew power bidirectional
flabel metal4 s 14746 1377 15000 2307 3 FreeSans 520 180 0 0 VCCD
port 5 nsew power bidirectional
flabel metal4 s 14807 2587 15000 3277 3 FreeSans 520 180 0 0 VDDA
port 6 nsew power bidirectional
flabel metal4 s 14746 9929 15000 10165 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 14746 9147 15000 9213 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 14746 11247 15000 12137 3 FreeSans 520 180 0 0 VSSIO_Q
port 7 nsew ground bidirectional
flabel metal4 s 14746 10881 15000 10947 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 14746 4767 15000 5697 3 FreeSans 520 180 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal4 s 14746 5977 15000 6667 3 FreeSans 520 180 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal4 s 14746 13607 15000 18600 3 FreeSans 520 180 0 0 VDDIO
port 2 nsew power bidirectional
flabel metal4 s 14746 12417 15000 13307 3 FreeSans 520 180 0 0 VDDIO_Q
port 1 nsew power bidirectional
flabel metal4 s 14746 10225 15000 10821 3 FreeSans 520 180 0 0 AMUXBUS_A
port 11 nsew signal bidirectional
flabel metal4 s 14746 9273 15000 9869 3 FreeSans 520 180 0 0 AMUXBUS_B
port 12 nsew signal bidirectional
flabel metal4 s 14746 7917 15000 8847 3 FreeSans 520 180 0 0 VSSD
port 10 nsew ground bidirectional
flabel metal4 s 14746 6947 15000 7637 3 FreeSans 520 180 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 14746 3557 15000 4487 3 FreeSans 520 180 0 0 VDDIO
port 2 nsew power bidirectional
flabel metal4 s 0 7 254 1097 3 FreeSans 520 0 0 0 VCCHIB
port 4 nsew power bidirectional
flabel metal4 s 0 1377 254 2307 3 FreeSans 520 0 0 0 VCCD
port 5 nsew power bidirectional
flabel metal4 s 0 2587 193 3277 3 FreeSans 520 0 0 0 VDDA
port 6 nsew power bidirectional
flabel metal4 s 0 9929 254 10165 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 0 9147 254 9213 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 0 11247 254 12137 3 FreeSans 520 0 0 0 VSSIO_Q
port 7 nsew ground bidirectional
flabel metal4 s 0 10881 254 10947 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 0 4767 254 5697 3 FreeSans 520 0 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal4 s 0 5977 254 6667 3 FreeSans 520 0 0 0 VSWITCH
port 8 nsew power bidirectional
flabel metal4 s 0 13607 254 18600 3 FreeSans 520 0 0 0 VDDIO
port 2 nsew power bidirectional
flabel metal4 s 0 12417 254 13307 3 FreeSans 520 0 0 0 VDDIO_Q
port 1 nsew power bidirectional
flabel metal4 s 0 10225 254 10821 3 FreeSans 520 0 0 0 AMUXBUS_A
port 11 nsew signal bidirectional
flabel metal4 s 0 9273 254 9869 3 FreeSans 520 0 0 0 AMUXBUS_B
port 12 nsew signal bidirectional
flabel metal4 s 0 7917 254 8847 3 FreeSans 520 0 0 0 VSSD
port 10 nsew ground bidirectional
flabel metal4 s 0 6947 254 7637 3 FreeSans 520 0 0 0 VSSA
port 3 nsew ground bidirectional
flabel metal4 s 14746 34757 15000 39600 3 FreeSans 520 180 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal4 s 14873 37932 14873 37932 3 FreeSans 520 180 0 0 VSSIO
port 9 nsew
flabel metal4 s 0 34757 254 39600 3 FreeSans 520 0 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal4 s 127 37932 127 37932 3 FreeSans 520 0 0 0 VSSIO
port 9 nsew
flabel metal4 s 0 3557 254 4487 3 FreeSans 520 0 0 0 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 10225 15000 10821 1 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 14746 9273 15000 9869 1 AMUXBUS_B
port 12 nsew signal bidirectional
rlabel metal3 s 10151 1378 14931 2306 1 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 0 1377 4895 2307 1 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 10156 1377 15000 2307 1 VCCD
port 5 nsew power bidirectional
rlabel metal5 s 0 1397 254 2287 1 VCCD
port 5 nsew power bidirectional
rlabel metal5 s 14746 1397 15000 2287 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14873 2252 14913 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14873 2166 14913 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14873 2080 14913 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14873 1994 14913 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14873 1908 14913 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14873 1822 14913 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14873 1736 14913 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14873 1650 14913 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14873 1564 14913 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14873 1478 14913 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14873 1392 14913 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14792 2252 14832 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14792 2166 14832 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14792 2080 14832 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14792 1994 14832 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14792 1908 14832 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14792 1822 14832 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14792 1736 14832 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14792 1650 14832 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14792 1564 14832 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14792 1478 14832 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14792 1392 14832 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14711 2252 14751 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14711 2166 14751 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14711 2080 14751 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14711 1994 14751 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14711 1908 14751 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14711 1822 14751 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14711 1736 14751 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14711 1650 14751 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14711 1564 14751 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14711 1478 14751 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14711 1392 14751 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14630 2252 14670 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14630 2166 14670 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14630 2080 14670 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14630 1994 14670 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14630 1908 14670 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14630 1822 14670 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14630 1736 14670 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14630 1650 14670 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14630 1564 14670 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14630 1478 14670 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14630 1392 14670 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14549 2252 14589 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14549 2166 14589 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14549 2080 14589 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14549 1994 14589 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14549 1908 14589 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14549 1822 14589 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14549 1736 14589 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14549 1650 14589 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14549 1564 14589 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14549 1478 14589 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14549 1392 14589 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14468 2252 14508 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14468 2166 14508 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14468 2080 14508 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14468 1994 14508 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14468 1908 14508 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14468 1822 14508 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14468 1736 14508 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14468 1650 14508 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14468 1564 14508 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14468 1478 14508 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14468 1392 14508 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14387 2252 14427 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14387 2166 14427 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14387 2080 14427 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14387 1994 14427 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14387 1908 14427 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14387 1822 14427 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14387 1736 14427 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14387 1650 14427 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14387 1564 14427 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14387 1478 14427 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14387 1392 14427 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14306 2252 14346 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14306 2166 14346 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14306 2080 14346 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14306 1994 14346 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14306 1908 14346 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14306 1822 14346 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14306 1736 14346 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14306 1650 14346 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14306 1564 14346 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14306 1478 14346 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14306 1392 14346 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14225 2252 14265 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14225 2166 14265 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14225 2080 14265 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14225 1994 14265 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14225 1908 14265 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14225 1822 14265 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14225 1736 14265 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14225 1650 14265 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14225 1564 14265 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14225 1478 14265 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14225 1392 14265 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14144 2252 14184 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14144 2166 14184 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14144 2080 14184 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14144 1994 14184 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14144 1908 14184 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14144 1822 14184 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14144 1736 14184 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14144 1650 14184 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14144 1564 14184 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14144 1478 14184 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14144 1392 14184 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14063 2252 14103 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14063 2166 14103 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14063 2080 14103 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14063 1994 14103 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14063 1908 14103 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14063 1822 14103 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14063 1736 14103 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14063 1650 14103 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14063 1564 14103 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14063 1478 14103 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 14063 1392 14103 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13982 2252 14022 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13982 2166 14022 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13982 2080 14022 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13982 1994 14022 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13982 1908 14022 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13982 1822 14022 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13982 1736 14022 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13982 1650 14022 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13982 1564 14022 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13982 1478 14022 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13982 1392 14022 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13901 2252 13941 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13901 2166 13941 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13901 2080 13941 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13901 1994 13941 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13901 1908 13941 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13901 1822 13941 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13901 1736 13941 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13901 1650 13941 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13901 1564 13941 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13901 1478 13941 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13901 1392 13941 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13820 2252 13860 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13820 2166 13860 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13820 2080 13860 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13820 1994 13860 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13820 1908 13860 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13820 1822 13860 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13820 1736 13860 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13820 1650 13860 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13820 1564 13860 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13820 1478 13860 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13820 1392 13860 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13739 2252 13779 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13739 2166 13779 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13739 2080 13779 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13739 1994 13779 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13739 1908 13779 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13739 1822 13779 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13739 1736 13779 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13739 1650 13779 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13739 1564 13779 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13739 1478 13779 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13739 1392 13779 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13658 2252 13698 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13658 2166 13698 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13658 2080 13698 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13658 1994 13698 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13658 1908 13698 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13658 1822 13698 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13658 1736 13698 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13658 1650 13698 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13658 1564 13698 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13658 1478 13698 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13658 1392 13698 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13577 2252 13617 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13577 2166 13617 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13577 2080 13617 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13577 1994 13617 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13577 1908 13617 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13577 1822 13617 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13577 1736 13617 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13577 1650 13617 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13577 1564 13617 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13577 1478 13617 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13577 1392 13617 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13496 2252 13536 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13496 2166 13536 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13496 2080 13536 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13496 1994 13536 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13496 1908 13536 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13496 1822 13536 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13496 1736 13536 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13496 1650 13536 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13496 1564 13536 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13496 1478 13536 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13496 1392 13536 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13415 2252 13455 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13415 2166 13455 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13415 2080 13455 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13415 1994 13455 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13415 1908 13455 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13415 1822 13455 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13415 1736 13455 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13415 1650 13455 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13415 1564 13455 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13415 1478 13455 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13415 1392 13455 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13334 2252 13374 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13334 2166 13374 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13334 2080 13374 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13334 1994 13374 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13334 1908 13374 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13334 1822 13374 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13334 1736 13374 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13334 1650 13374 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13334 1564 13374 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13334 1478 13374 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13334 1392 13374 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13253 2252 13293 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13253 2166 13293 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13253 2080 13293 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13253 1994 13293 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13253 1908 13293 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13253 1822 13293 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13253 1736 13293 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13253 1650 13293 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13253 1564 13293 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13253 1478 13293 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13253 1392 13293 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13172 2252 13212 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13172 2166 13212 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13172 2080 13212 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13172 1994 13212 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13172 1908 13212 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13172 1822 13212 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13172 1736 13212 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13172 1650 13212 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13172 1564 13212 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13172 1478 13212 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13172 1392 13212 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13091 2252 13131 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13091 2166 13131 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13091 2080 13131 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13091 1994 13131 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13091 1908 13131 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13091 1822 13131 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13091 1736 13131 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13091 1650 13131 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13091 1564 13131 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13091 1478 13131 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13091 1392 13131 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13010 2252 13050 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13010 2166 13050 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13010 2080 13050 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13010 1994 13050 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13010 1908 13050 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13010 1822 13050 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13010 1736 13050 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13010 1650 13050 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13010 1564 13050 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13010 1478 13050 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 13010 1392 13050 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12929 2252 12969 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12929 2166 12969 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12929 2080 12969 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12929 1994 12969 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12929 1908 12969 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12929 1822 12969 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12929 1736 12969 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12929 1650 12969 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12929 1564 12969 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12929 1478 12969 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12929 1392 12969 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12848 2252 12888 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12848 2166 12888 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12848 2080 12888 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12848 1994 12888 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12848 1908 12888 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12848 1822 12888 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12848 1736 12888 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12848 1650 12888 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12848 1564 12888 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12848 1478 12888 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12848 1392 12888 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12767 2252 12807 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12767 2166 12807 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12767 2080 12807 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12767 1994 12807 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12767 1908 12807 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12767 1822 12807 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12767 1736 12807 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12767 1650 12807 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12767 1564 12807 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12767 1478 12807 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12767 1392 12807 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12686 2252 12726 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12686 2166 12726 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12686 2080 12726 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12686 1994 12726 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12686 1908 12726 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12686 1822 12726 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12686 1736 12726 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12686 1650 12726 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12686 1564 12726 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12686 1478 12726 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12686 1392 12726 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12605 2252 12645 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12605 2166 12645 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12605 2080 12645 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12605 1994 12645 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12605 1908 12645 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12605 1822 12645 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12605 1736 12645 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12605 1650 12645 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12605 1564 12645 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12605 1478 12645 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12605 1392 12645 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12524 2252 12564 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12524 2166 12564 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12524 2080 12564 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12524 1994 12564 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12524 1908 12564 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12524 1822 12564 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12524 1736 12564 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12524 1650 12564 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12524 1564 12564 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12524 1478 12564 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12524 1392 12564 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12443 2252 12483 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12443 2166 12483 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12443 2080 12483 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12443 1994 12483 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12443 1908 12483 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12443 1822 12483 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12443 1736 12483 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12443 1650 12483 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12443 1564 12483 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12443 1478 12483 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12443 1392 12483 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12362 2252 12402 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12362 2166 12402 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12362 2080 12402 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12362 1994 12402 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12362 1908 12402 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12362 1822 12402 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12362 1736 12402 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12362 1650 12402 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12362 1564 12402 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12362 1478 12402 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12362 1392 12402 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12281 2252 12321 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12281 2166 12321 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12281 2080 12321 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12281 1994 12321 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12281 1908 12321 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12281 1822 12321 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12281 1736 12321 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12281 1650 12321 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12281 1564 12321 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12281 1478 12321 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12281 1392 12321 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12200 2252 12240 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12200 2166 12240 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12200 2080 12240 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12200 1994 12240 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12200 1908 12240 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12200 1822 12240 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12200 1736 12240 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12200 1650 12240 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12200 1564 12240 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12200 1478 12240 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12200 1392 12240 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12119 2252 12159 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12119 2166 12159 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12119 2080 12159 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12119 1994 12159 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12119 1908 12159 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12119 1822 12159 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12119 1736 12159 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12119 1650 12159 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12119 1564 12159 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12119 1478 12159 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12119 1392 12159 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12038 2252 12078 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12038 2166 12078 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12038 2080 12078 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12038 1994 12078 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12038 1908 12078 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12038 1822 12078 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12038 1736 12078 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12038 1650 12078 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12038 1564 12078 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12038 1478 12078 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 12038 1392 12078 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11957 2252 11997 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11957 2166 11997 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11957 2080 11997 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11957 1994 11997 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11957 1908 11997 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11957 1822 11997 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11957 1736 11997 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11957 1650 11997 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11957 1564 11997 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11957 1478 11997 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11957 1392 11997 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11876 2252 11916 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11876 2166 11916 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11876 2080 11916 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11876 1994 11916 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11876 1908 11916 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11876 1822 11916 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11876 1736 11916 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11876 1650 11916 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11876 1564 11916 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11876 1478 11916 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11876 1392 11916 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11795 2252 11835 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11795 2166 11835 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11795 2080 11835 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11795 1994 11835 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11795 1908 11835 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11795 1822 11835 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11795 1736 11835 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11795 1650 11835 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11795 1564 11835 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11795 1478 11835 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11795 1392 11835 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11714 2252 11754 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11714 2166 11754 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11714 2080 11754 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11714 1994 11754 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11714 1908 11754 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11714 1822 11754 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11714 1736 11754 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11714 1650 11754 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11714 1564 11754 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11714 1478 11754 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11714 1392 11754 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11633 2252 11673 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11633 2166 11673 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11633 2080 11673 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11633 1994 11673 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11633 1908 11673 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11633 1822 11673 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11633 1736 11673 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11633 1650 11673 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11633 1564 11673 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11633 1478 11673 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11633 1392 11673 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11552 2252 11592 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11552 2166 11592 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11552 2080 11592 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11552 1994 11592 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11552 1908 11592 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11552 1822 11592 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11552 1736 11592 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11552 1650 11592 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11552 1564 11592 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11552 1478 11592 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11552 1392 11592 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11471 2252 11511 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11471 2166 11511 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11471 2080 11511 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11471 1994 11511 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11471 1908 11511 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11471 1822 11511 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11471 1736 11511 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11471 1650 11511 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11471 1564 11511 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11471 1478 11511 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11471 1392 11511 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11390 2252 11430 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11390 2166 11430 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11390 2080 11430 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11390 1994 11430 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11390 1908 11430 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11390 1822 11430 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11390 1736 11430 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11390 1650 11430 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11390 1564 11430 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11390 1478 11430 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11390 1392 11430 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11309 2252 11349 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11309 2166 11349 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11309 2080 11349 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11309 1994 11349 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11309 1908 11349 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11309 1822 11349 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11309 1736 11349 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11309 1650 11349 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11309 1564 11349 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11309 1478 11349 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11309 1392 11349 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11228 2252 11268 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11228 2166 11268 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11228 2080 11268 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11228 1994 11268 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11228 1908 11268 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11228 1822 11268 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11228 1736 11268 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11228 1650 11268 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11228 1564 11268 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11228 1478 11268 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11228 1392 11268 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11147 2252 11187 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11147 2166 11187 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11147 2080 11187 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11147 1994 11187 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11147 1908 11187 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11147 1822 11187 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11147 1736 11187 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11147 1650 11187 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11147 1564 11187 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11147 1478 11187 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11147 1392 11187 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11066 2252 11106 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11066 2166 11106 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11066 2080 11106 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11066 1994 11106 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11066 1908 11106 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11066 1822 11106 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11066 1736 11106 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11066 1650 11106 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11066 1564 11106 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11066 1478 11106 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 11066 1392 11106 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10985 2252 11025 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10985 2166 11025 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10985 2080 11025 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10985 1994 11025 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10985 1908 11025 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10985 1822 11025 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10985 1736 11025 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10985 1650 11025 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10985 1564 11025 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10985 1478 11025 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10985 1392 11025 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10904 2252 10944 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10904 2166 10944 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10904 2080 10944 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10904 1994 10944 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10904 1908 10944 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10904 1822 10944 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10904 1736 10944 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10904 1650 10944 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10904 1564 10944 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10904 1478 10944 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10904 1392 10944 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10823 2252 10863 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10823 2166 10863 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10823 2080 10863 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10823 1994 10863 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10823 1908 10863 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10823 1822 10863 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10823 1736 10863 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10823 1650 10863 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10823 1564 10863 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10823 1478 10863 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10823 1392 10863 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10742 2252 10782 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10742 2166 10782 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10742 2080 10782 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10742 1994 10782 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10742 1908 10782 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10742 1822 10782 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10742 1736 10782 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10742 1650 10782 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10742 1564 10782 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10742 1478 10782 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10742 1392 10782 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10661 2252 10701 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10661 2166 10701 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10661 2080 10701 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10661 1994 10701 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10661 1908 10701 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10661 1822 10701 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10661 1736 10701 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10661 1650 10701 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10661 1564 10701 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10661 1478 10701 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10661 1392 10701 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10579 2252 10619 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10579 2166 10619 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10579 2080 10619 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10579 1994 10619 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10579 1908 10619 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10579 1822 10619 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10579 1736 10619 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10579 1650 10619 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10579 1564 10619 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10579 1478 10619 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10579 1392 10619 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10497 2252 10537 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10497 2166 10537 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10497 2080 10537 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10497 1994 10537 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10497 1908 10537 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10497 1822 10537 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10497 1736 10537 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10497 1650 10537 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10497 1564 10537 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10497 1478 10537 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10497 1392 10537 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10415 2252 10455 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10415 2166 10455 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10415 2080 10455 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10415 1994 10455 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10415 1908 10455 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10415 1822 10455 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10415 1736 10455 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10415 1650 10455 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10415 1564 10455 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10415 1478 10455 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10415 1392 10455 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10333 2252 10373 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10333 2166 10373 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10333 2080 10373 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10333 1994 10373 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10333 1908 10373 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10333 1822 10373 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10333 1736 10373 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10333 1650 10373 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10333 1564 10373 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10333 1478 10373 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10333 1392 10373 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10251 2252 10291 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10251 2166 10291 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10251 2080 10291 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10251 1994 10291 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10251 1908 10291 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10251 1822 10291 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10251 1736 10291 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10251 1650 10291 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10251 1564 10291 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10251 1478 10291 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10251 1392 10291 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10169 2252 10209 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10169 2166 10209 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10169 2080 10209 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10169 1994 10209 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10169 1908 10209 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10169 1822 10209 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10169 1736 10209 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10169 1650 10209 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10169 1564 10209 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10169 1478 10209 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 10169 1392 10209 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4842 2252 4882 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4842 2166 4882 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4842 2080 4882 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4842 1994 4882 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4842 1908 4882 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4842 1822 4882 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4842 1736 4882 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4842 1650 4882 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4842 1564 4882 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4842 1478 4882 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4842 1392 4882 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4761 2252 4801 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4761 2166 4801 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4761 2080 4801 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4761 1994 4801 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4761 1908 4801 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4761 1822 4801 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4761 1736 4801 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4761 1650 4801 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4761 1564 4801 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4761 1478 4801 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4761 1392 4801 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4680 2252 4720 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4680 2166 4720 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4680 2080 4720 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4680 1994 4720 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4680 1908 4720 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4680 1822 4720 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4680 1736 4720 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4680 1650 4720 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4680 1564 4720 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4680 1478 4720 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4680 1392 4720 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4599 2252 4639 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4599 2166 4639 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4599 2080 4639 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4599 1994 4639 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4599 1908 4639 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4599 1822 4639 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4599 1736 4639 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4599 1650 4639 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4599 1564 4639 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4599 1478 4639 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4599 1392 4639 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4518 2252 4558 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4518 2166 4558 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4518 2080 4558 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4518 1994 4558 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4518 1908 4558 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4518 1822 4558 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4518 1736 4558 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4518 1650 4558 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4518 1564 4558 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4518 1478 4558 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4518 1392 4558 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4437 2252 4477 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4437 2166 4477 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4437 2080 4477 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4437 1994 4477 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4437 1908 4477 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4437 1822 4477 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4437 1736 4477 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4437 1650 4477 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4437 1564 4477 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4437 1478 4477 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4437 1392 4477 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4356 2252 4396 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4356 2166 4396 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4356 2080 4396 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4356 1994 4396 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4356 1908 4396 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4356 1822 4396 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4356 1736 4396 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4356 1650 4396 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4356 1564 4396 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4356 1478 4396 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4356 1392 4396 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4275 2252 4315 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4275 2166 4315 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4275 2080 4315 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4275 1994 4315 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4275 1908 4315 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4275 1822 4315 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4275 1736 4315 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4275 1650 4315 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4275 1564 4315 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4275 1478 4315 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4275 1392 4315 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4194 2252 4234 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4194 2166 4234 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4194 2080 4234 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4194 1994 4234 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4194 1908 4234 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4194 1822 4234 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4194 1736 4234 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4194 1650 4234 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4194 1564 4234 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4194 1478 4234 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4194 1392 4234 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4113 2252 4153 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4113 2166 4153 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4113 2080 4153 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4113 1994 4153 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4113 1908 4153 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4113 1822 4153 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4113 1736 4153 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4113 1650 4153 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4113 1564 4153 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4113 1478 4153 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4113 1392 4153 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4032 2252 4072 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4032 2166 4072 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4032 2080 4072 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4032 1994 4072 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4032 1908 4072 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4032 1822 4072 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4032 1736 4072 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4032 1650 4072 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4032 1564 4072 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4032 1478 4072 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 4032 1392 4072 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3951 2252 3991 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3951 2166 3991 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3951 2080 3991 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3951 1994 3991 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3951 1908 3991 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3951 1822 3991 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3951 1736 3991 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3951 1650 3991 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3951 1564 3991 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3951 1478 3991 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3951 1392 3991 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3870 2252 3910 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3870 2166 3910 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3870 2080 3910 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3870 1994 3910 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3870 1908 3910 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3870 1822 3910 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3870 1736 3910 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3870 1650 3910 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3870 1564 3910 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3870 1478 3910 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3870 1392 3910 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3789 2252 3829 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3789 2166 3829 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3789 2080 3829 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3789 1994 3829 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3789 1908 3829 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3789 1822 3829 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3789 1736 3829 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3789 1650 3829 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3789 1564 3829 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3789 1478 3829 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3789 1392 3829 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3708 2252 3748 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3708 2166 3748 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3708 2080 3748 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3708 1994 3748 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3708 1908 3748 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3708 1822 3748 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3708 1736 3748 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3708 1650 3748 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3708 1564 3748 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3708 1478 3748 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3708 1392 3748 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3627 2252 3667 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3627 2166 3667 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3627 2080 3667 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3627 1994 3667 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3627 1908 3667 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3627 1822 3667 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3627 1736 3667 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3627 1650 3667 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3627 1564 3667 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3627 1478 3667 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3627 1392 3667 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3546 2252 3586 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3546 2166 3586 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3546 2080 3586 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3546 1994 3586 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3546 1908 3586 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3546 1822 3586 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3546 1736 3586 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3546 1650 3586 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3546 1564 3586 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3546 1478 3586 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3546 1392 3586 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3465 2252 3505 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3465 2166 3505 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3465 2080 3505 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3465 1994 3505 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3465 1908 3505 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3465 1822 3505 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3465 1736 3505 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3465 1650 3505 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3465 1564 3505 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3465 1478 3505 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3465 1392 3505 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3384 2252 3424 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3384 2166 3424 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3384 2080 3424 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3384 1994 3424 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3384 1908 3424 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3384 1822 3424 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3384 1736 3424 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3384 1650 3424 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3384 1564 3424 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3384 1478 3424 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3384 1392 3424 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3303 2252 3343 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3303 2166 3343 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3303 2080 3343 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3303 1994 3343 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3303 1908 3343 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3303 1822 3343 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3303 1736 3343 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3303 1650 3343 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3303 1564 3343 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3303 1478 3343 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3303 1392 3343 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3222 2252 3262 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3222 2166 3262 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3222 2080 3262 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3222 1994 3262 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3222 1908 3262 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3222 1822 3262 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3222 1736 3262 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3222 1650 3262 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3222 1564 3262 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3222 1478 3262 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3222 1392 3262 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3141 2252 3181 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3141 2166 3181 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3141 2080 3181 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3141 1994 3181 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3141 1908 3181 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3141 1822 3181 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3141 1736 3181 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3141 1650 3181 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3141 1564 3181 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3141 1478 3181 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3141 1392 3181 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3060 2252 3100 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3060 2166 3100 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3060 2080 3100 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3060 1994 3100 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3060 1908 3100 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3060 1822 3100 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3060 1736 3100 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3060 1650 3100 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3060 1564 3100 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3060 1478 3100 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 3060 1392 3100 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2979 2252 3019 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2979 2166 3019 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2979 2080 3019 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2979 1994 3019 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2979 1908 3019 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2979 1822 3019 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2979 1736 3019 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2979 1650 3019 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2979 1564 3019 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2979 1478 3019 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2979 1392 3019 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2898 2252 2938 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2898 2166 2938 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2898 2080 2938 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2898 1994 2938 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2898 1908 2938 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2898 1822 2938 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2898 1736 2938 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2898 1650 2938 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2898 1564 2938 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2898 1478 2938 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2898 1392 2938 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2817 2252 2857 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2817 2166 2857 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2817 2080 2857 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2817 1994 2857 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2817 1908 2857 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2817 1822 2857 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2817 1736 2857 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2817 1650 2857 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2817 1564 2857 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2817 1478 2857 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2817 1392 2857 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2736 2252 2776 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2736 2166 2776 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2736 2080 2776 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2736 1994 2776 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2736 1908 2776 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2736 1822 2776 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2736 1736 2776 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2736 1650 2776 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2736 1564 2776 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2736 1478 2776 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2736 1392 2776 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2655 2252 2695 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2655 2166 2695 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2655 2080 2695 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2655 1994 2695 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2655 1908 2695 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2655 1822 2695 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2655 1736 2695 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2655 1650 2695 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2655 1564 2695 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2655 1478 2695 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2655 1392 2695 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2574 2252 2614 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2574 2166 2614 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2574 2080 2614 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2574 1994 2614 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2574 1908 2614 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2574 1822 2614 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2574 1736 2614 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2574 1650 2614 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2574 1564 2614 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2574 1478 2614 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2574 1392 2614 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2493 2252 2533 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2493 2166 2533 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2493 2080 2533 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2493 1994 2533 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2493 1908 2533 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2493 1822 2533 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2493 1736 2533 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2493 1650 2533 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2493 1564 2533 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2493 1478 2533 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2493 1392 2533 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2412 2252 2452 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2412 2166 2452 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2412 2080 2452 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2412 1994 2452 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2412 1908 2452 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2412 1822 2452 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2412 1736 2452 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2412 1650 2452 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2412 1564 2452 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2412 1478 2452 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2412 1392 2452 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2331 2252 2371 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2331 2166 2371 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2331 2080 2371 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2331 1994 2371 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2331 1908 2371 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2331 1822 2371 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2331 1736 2371 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2331 1650 2371 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2331 1564 2371 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2331 1478 2371 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2331 1392 2371 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2250 2252 2290 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2250 2166 2290 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2250 2080 2290 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2250 1994 2290 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2250 1908 2290 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2250 1822 2290 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2250 1736 2290 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2250 1650 2290 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2250 1564 2290 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2250 1478 2290 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2250 1392 2290 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2169 2252 2209 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2169 2166 2209 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2169 2080 2209 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2169 1994 2209 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2169 1908 2209 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2169 1822 2209 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2169 1736 2209 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2169 1650 2209 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2169 1564 2209 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2169 1478 2209 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2169 1392 2209 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2088 2252 2128 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2088 2166 2128 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2088 2080 2128 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2088 1994 2128 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2088 1908 2128 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2088 1822 2128 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2088 1736 2128 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2088 1650 2128 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2088 1564 2128 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2088 1478 2128 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2088 1392 2128 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2007 2252 2047 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2007 2166 2047 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2007 2080 2047 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2007 1994 2047 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2007 1908 2047 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2007 1822 2047 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2007 1736 2047 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2007 1650 2047 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2007 1564 2047 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2007 1478 2047 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 2007 1392 2047 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1926 2252 1966 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1926 2166 1966 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1926 2080 1966 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1926 1994 1966 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1926 1908 1966 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1926 1822 1966 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1926 1736 1966 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1926 1650 1966 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1926 1564 1966 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1926 1478 1966 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1926 1392 1966 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1845 2252 1885 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1845 2166 1885 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1845 2080 1885 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1845 1994 1885 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1845 1908 1885 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1845 1822 1885 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1845 1736 1885 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1845 1650 1885 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1845 1564 1885 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1845 1478 1885 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1845 1392 1885 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1764 2252 1804 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1764 2166 1804 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1764 2080 1804 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1764 1994 1804 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1764 1908 1804 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1764 1822 1804 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1764 1736 1804 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1764 1650 1804 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1764 1564 1804 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1764 1478 1804 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1764 1392 1804 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1683 2252 1723 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1683 2166 1723 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1683 2080 1723 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1683 1994 1723 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1683 1908 1723 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1683 1822 1723 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1683 1736 1723 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1683 1650 1723 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1683 1564 1723 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1683 1478 1723 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1683 1392 1723 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1602 2252 1642 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1602 2166 1642 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1602 2080 1642 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1602 1994 1642 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1602 1908 1642 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1602 1822 1642 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1602 1736 1642 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1602 1650 1642 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1602 1564 1642 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1602 1478 1642 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1602 1392 1642 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1521 2252 1561 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1521 2166 1561 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1521 2080 1561 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1521 1994 1561 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1521 1908 1561 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1521 1822 1561 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1521 1736 1561 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1521 1650 1561 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1521 1564 1561 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1521 1478 1561 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1521 1392 1561 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1440 2252 1480 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1440 2166 1480 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1440 2080 1480 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1440 1994 1480 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1440 1908 1480 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1440 1822 1480 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1440 1736 1480 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1440 1650 1480 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1440 1564 1480 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1440 1478 1480 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1440 1392 1480 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1359 2252 1399 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1359 2166 1399 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1359 2080 1399 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1359 1994 1399 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1359 1908 1399 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1359 1822 1399 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1359 1736 1399 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1359 1650 1399 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1359 1564 1399 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1359 1478 1399 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1359 1392 1399 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1278 2252 1318 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1278 2166 1318 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1278 2080 1318 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1278 1994 1318 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1278 1908 1318 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1278 1822 1318 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1278 1736 1318 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1278 1650 1318 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1278 1564 1318 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1278 1478 1318 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1278 1392 1318 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1197 2252 1237 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1197 2166 1237 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1197 2080 1237 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1197 1994 1237 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1197 1908 1237 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1197 1822 1237 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1197 1736 1237 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1197 1650 1237 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1197 1564 1237 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1197 1478 1237 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1197 1392 1237 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1116 2252 1156 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1116 2166 1156 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1116 2080 1156 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1116 1994 1156 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1116 1908 1156 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1116 1822 1156 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1116 1736 1156 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1116 1650 1156 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1116 1564 1156 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1116 1478 1156 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1116 1392 1156 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1035 2252 1075 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1035 2166 1075 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1035 2080 1075 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1035 1994 1075 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1035 1908 1075 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1035 1822 1075 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1035 1736 1075 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1035 1650 1075 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1035 1564 1075 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1035 1478 1075 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 1035 1392 1075 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 954 2252 994 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 954 2166 994 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 954 2080 994 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 954 1994 994 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 954 1908 994 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 954 1822 994 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 954 1736 994 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 954 1650 994 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 954 1564 994 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 954 1478 994 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 954 1392 994 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 873 2252 913 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 873 2166 913 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 873 2080 913 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 873 1994 913 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 873 1908 913 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 873 1822 913 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 873 1736 913 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 873 1650 913 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 873 1564 913 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 873 1478 913 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 873 1392 913 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 792 2252 832 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 792 2166 832 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 792 2080 832 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 792 1994 832 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 792 1908 832 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 792 1822 832 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 792 1736 832 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 792 1650 832 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 792 1564 832 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 792 1478 832 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 792 1392 832 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 711 2252 751 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 711 2166 751 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 711 2080 751 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 711 1994 751 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 711 1908 751 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 711 1822 751 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 711 1736 751 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 711 1650 751 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 711 1564 751 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 711 1478 751 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 711 1392 751 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 630 2252 670 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 630 2166 670 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 630 2080 670 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 630 1994 670 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 630 1908 670 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 630 1822 670 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 630 1736 670 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 630 1650 670 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 630 1564 670 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 630 1478 670 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 630 1392 670 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 548 2252 588 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 548 2166 588 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 548 2080 588 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 548 1994 588 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 548 1908 588 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 548 1822 588 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 548 1736 588 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 548 1650 588 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 548 1564 588 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 548 1478 588 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 548 1392 588 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 466 2252 506 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 466 2166 506 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 466 2080 506 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 466 1994 506 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 466 1908 506 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 466 1822 506 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 466 1736 506 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 466 1650 506 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 466 1564 506 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 466 1478 506 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 466 1392 506 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 384 2252 424 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 384 2166 424 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 384 2080 424 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 384 1994 424 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 384 1908 424 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 384 1822 424 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 384 1736 424 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 384 1650 424 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 384 1564 424 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 384 1478 424 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 384 1392 424 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 302 2252 342 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 302 2166 342 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 302 2080 342 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 302 1994 342 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 302 1908 342 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 302 1822 342 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 302 1736 342 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 302 1650 342 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 302 1564 342 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 302 1478 342 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 302 1392 342 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 220 2252 260 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 220 2166 260 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 220 2080 260 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 220 1994 260 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 220 1908 260 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 220 1822 260 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 220 1736 260 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 220 1650 260 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 220 1564 260 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 220 1478 260 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 220 1392 260 1432 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 138 2252 178 2292 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 138 2166 178 2206 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 138 2080 178 2120 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 138 1994 178 2034 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 138 1908 178 1948 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 138 1822 178 1862 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 138 1736 178 1776 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 138 1650 178 1690 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 138 1564 178 1604 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 138 1478 178 1518 1 VCCD
port 5 nsew power bidirectional
rlabel via3 s 138 1392 178 1432 1 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 1 VCCHIB
port 4 nsew power bidirectional
rlabel metal5 s 0 27 254 1077 1 VCCHIB
port 4 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 1 VCCHIB
port 4 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 1 VDDA
port 6 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 1 VDDA
port 6 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 1 VDDA
port 6 nsew power bidirectional
rlabel metal4 s 0 13607 254 18600 1 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 3557 15000 4487 1 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 18600 1 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 1 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 1 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 1 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 13607 15000 18597 1 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 12417 15000 13307 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 0 12437 254 13287 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 0 9147 254 9213 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10881 254 10947 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 9147 15000 9213 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 10881 15000 10947 1 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 1 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 9147 254 10947 1 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 1 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 9147 15000 10947 1 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 1 VSSD
port 10 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 1 VSSD
port 10 nsew ground bidirectional
rlabel metal5 s 14746 7937 15000 8827 1 VSSD
port 10 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 1 VSSIO
port 9 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 1 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 1 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 1 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 1 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 1 VSSIO
port 9 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 1 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 0 11267 254 12117 1 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 1 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14746 5977 15000 6667 1 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 0 5997 254 6647 1 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 14746 5997 15000 6647 1 VSWITCH
port 8 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 15000 39600
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string LEFsymmetry X Y R90
string GDS_END 538092
string GDS_START 446284
<< end >>
