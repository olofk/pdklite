magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1245 -1243 3285 1278
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_0
timestamp 1619729480
transform -1 0 16 0 1 17
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_1
timestamp 1619729480
transform 1 0 2024 0 1 17
box 0 0 1 1
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 1339954
string GDS_START 1339472
<< end >>
