magic
tech sky130A
magscale 1 2
timestamp 1640697996
<< nwell >>
rect -66 377 1986 897
<< pwell >>
rect 23 43 1901 317
rect -26 -43 1946 43
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1920 831
rect 123 729 1901 759
rect 157 695 195 729
rect 229 695 267 729
rect 301 695 339 729
rect 373 725 554 729
rect 123 489 373 695
rect 553 695 554 725
rect 588 695 626 729
rect 660 725 821 729
rect 660 695 687 725
rect 553 477 687 695
rect 855 695 893 729
rect 927 695 965 729
rect 999 725 1133 729
rect 821 477 999 695
rect 1167 695 1205 729
rect 1239 695 1277 729
rect 1311 725 1446 729
rect 1133 477 1311 695
rect 1445 695 1446 725
rect 1480 695 1589 729
rect 1623 725 1853 729
rect 1781 695 1853 725
rect 1887 695 1901 729
rect 1445 477 1623 695
rect 1827 477 1901 695
rect 127 316 449 363
rect 135 110 385 277
rect 553 152 699 289
rect 521 110 699 152
rect 809 110 1011 289
rect 1121 110 1323 289
rect 1433 110 1635 289
rect 1827 120 1901 289
rect 1795 110 1901 120
rect 135 76 207 110
rect 241 76 279 110
rect 313 76 351 110
rect 385 76 521 110
rect 555 76 593 110
rect 627 76 665 110
rect 699 76 814 110
rect 848 76 886 110
rect 920 76 958 110
rect 992 76 1134 110
rect 1168 76 1206 110
rect 1240 76 1278 110
rect 1312 76 1447 110
rect 1481 76 1519 110
rect 1553 76 1591 110
rect 1625 76 1795 110
rect 1829 76 1867 110
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 123 695 157 729
rect 195 695 229 729
rect 267 695 301 729
rect 339 695 373 729
rect 554 695 588 729
rect 626 695 660 729
rect 821 695 855 729
rect 893 695 927 729
rect 965 695 999 729
rect 1133 695 1167 729
rect 1205 695 1239 729
rect 1277 695 1311 729
rect 1446 695 1480 729
rect 1589 695 1623 729
rect 1853 695 1887 729
rect 207 76 241 110
rect 279 76 313 110
rect 351 76 385 110
rect 521 76 555 110
rect 593 76 627 110
rect 665 76 699 110
rect 814 76 848 110
rect 886 76 920 110
rect 958 76 992 110
rect 1134 76 1168 110
rect 1206 76 1240 110
rect 1278 76 1312 110
rect 1447 76 1481 110
rect 1519 76 1553 110
rect 1591 76 1625 110
rect 1795 76 1829 110
rect 1867 76 1901 110
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< obsli1 >>
rect 49 453 87 709
rect 409 453 519 689
rect 49 419 519 453
rect 49 295 87 419
rect 485 391 519 419
rect 721 441 787 689
rect 1033 441 1099 689
rect 1345 441 1411 689
rect 1657 646 1747 689
rect 1657 441 1793 646
rect 721 424 1793 441
rect 721 391 1124 424
rect 485 325 676 391
rect 733 390 1124 391
rect 1158 390 1196 424
rect 1230 390 1793 424
rect 733 325 1793 390
rect 49 161 91 295
rect 485 280 519 325
rect 421 246 519 280
rect 421 146 463 246
rect 733 161 775 325
rect 1045 161 1087 325
rect 1357 161 1399 325
rect 1669 161 1793 325
<< obsli1c >>
rect 1124 390 1158 424
rect 1196 390 1230 424
<< metal1 >>
rect 0 831 1920 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1920 831
rect 0 791 1920 797
rect 0 753 1920 763
rect 0 729 1862 753
rect 0 695 123 729
rect 157 695 195 729
rect 229 695 267 729
rect 301 695 339 729
rect 373 695 554 729
rect 588 695 626 729
rect 660 695 821 729
rect 855 695 893 729
rect 927 695 965 729
rect 999 695 1133 729
rect 1167 695 1205 729
rect 1239 695 1277 729
rect 1311 695 1446 729
rect 1480 695 1589 729
rect 1623 695 1853 729
rect 1914 701 1926 753
rect 1978 701 1984 753
rect 1887 695 1920 701
rect 0 689 1920 695
rect 1112 381 1120 433
rect 1172 381 1184 433
rect 1236 381 1242 433
rect 0 113 1920 125
rect 0 110 1862 113
rect 0 76 207 110
rect 241 76 279 110
rect 313 76 351 110
rect 385 76 521 110
rect 555 76 593 110
rect 627 76 665 110
rect 699 76 814 110
rect 848 76 886 110
rect 920 76 958 110
rect 992 76 1134 110
rect 1168 76 1206 110
rect 1240 76 1278 110
rect 1312 76 1447 110
rect 1481 76 1519 110
rect 1553 76 1591 110
rect 1625 76 1795 110
rect 1829 76 1862 110
rect 0 61 1862 76
rect 1914 61 1926 113
rect 1978 61 1984 113
rect 0 51 1920 61
rect 0 17 1920 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -23 1920 -17
<< via1 >>
rect 1862 729 1914 753
rect 1862 701 1887 729
rect 1887 701 1914 729
rect 1926 701 1978 753
rect 1120 424 1172 433
rect 1120 390 1124 424
rect 1124 390 1158 424
rect 1158 390 1172 424
rect 1120 381 1172 390
rect 1184 424 1236 433
rect 1184 390 1196 424
rect 1196 390 1230 424
rect 1230 390 1236 424
rect 1184 381 1236 390
rect 1862 110 1914 113
rect 1862 76 1867 110
rect 1867 76 1901 110
rect 1901 76 1914 110
rect 1862 61 1914 76
rect 1926 61 1978 113
<< metal2 >>
rect 1843 701 1852 757
rect 1908 753 1932 757
rect 1914 701 1926 753
rect 1988 701 1997 757
rect 1088 379 1097 435
rect 1153 433 1177 435
rect 1233 433 1242 435
rect 1172 381 1177 433
rect 1236 381 1242 433
rect 1153 379 1177 381
rect 1233 379 1242 381
rect 1843 57 1852 113
rect 1914 61 1926 113
rect 1908 57 1932 61
rect 1988 57 1997 113
<< via2 >>
rect 1852 753 1908 757
rect 1932 753 1988 757
rect 1852 701 1862 753
rect 1862 701 1908 753
rect 1932 701 1978 753
rect 1978 701 1988 753
rect 1097 433 1153 435
rect 1177 433 1233 435
rect 1097 381 1120 433
rect 1120 381 1153 433
rect 1177 381 1184 433
rect 1184 381 1233 433
rect 1097 379 1153 381
rect 1177 379 1233 381
rect 1852 61 1862 113
rect 1862 61 1908 113
rect 1932 61 1978 113
rect 1978 61 1988 113
rect 1852 57 1908 61
rect 1932 57 1988 61
<< metal3 >>
rect 1842 761 1998 762
rect 1842 697 1848 761
rect 1912 697 1928 761
rect 1992 697 1998 761
rect 1842 696 1998 697
rect 1087 439 1243 440
rect 567 375 573 439
rect 637 375 653 439
rect 717 375 723 439
rect 1087 375 1093 439
rect 1157 375 1173 439
rect 1237 375 1243 439
rect 1087 374 1243 375
rect 1842 117 1998 118
rect 1842 53 1848 117
rect 1912 53 1928 117
rect 1992 53 1998 117
rect 1842 52 1998 53
<< via3 >>
rect 1848 757 1912 761
rect 1848 701 1852 757
rect 1852 701 1908 757
rect 1908 701 1912 757
rect 1848 697 1912 701
rect 1928 757 1992 761
rect 1928 701 1932 757
rect 1932 701 1988 757
rect 1988 701 1992 757
rect 1928 697 1992 701
rect 573 375 637 439
rect 653 375 717 439
rect 1093 435 1157 439
rect 1093 379 1097 435
rect 1097 379 1153 435
rect 1153 379 1157 435
rect 1093 375 1157 379
rect 1173 435 1237 439
rect 1173 379 1177 435
rect 1177 379 1233 435
rect 1233 379 1237 435
rect 1173 375 1237 379
rect 1848 113 1912 117
rect 1848 57 1852 113
rect 1852 57 1908 113
rect 1908 57 1912 113
rect 1848 53 1912 57
rect 1928 113 1992 117
rect 1928 57 1932 113
rect 1932 57 1988 113
rect 1988 57 1992 113
rect 1928 53 1992 57
<< metal4 >>
rect 1802 761 2038 845
rect 1802 697 1848 761
rect 1912 697 1928 761
rect 1992 697 2038 761
rect 1802 609 2038 697
rect 482 439 718 525
rect 482 375 573 439
rect 637 375 653 439
rect 717 375 718 439
rect 482 289 718 375
rect 1002 439 1238 525
rect 1002 375 1093 439
rect 1157 375 1173 439
rect 1237 375 1238 439
rect 1002 289 1238 375
rect 1802 117 2038 205
rect 1802 53 1848 117
rect 1912 53 1928 117
rect 1992 53 2038 117
rect 1802 -31 2038 53
<< metal5 >>
rect 942 567 1262 887
rect 1582 567 2082 887
rect 458 247 1262 567
rect 942 -73 1262 247
rect 1582 -73 2082 247
<< labels >>
rlabel locali s 127 316 449 363 6 A
port 1 nsew signal input
rlabel metal5 s 1582 -73 2082 247 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 1802 -31 2038 205 6 VGND
port 2 nsew ground bidirectional
rlabel via3 s 1928 53 1992 117 6 VGND
port 2 nsew ground bidirectional
rlabel via3 s 1848 53 1912 117 6 VGND
port 2 nsew ground bidirectional
rlabel metal3 s 1842 52 1998 118 6 VGND
port 2 nsew ground bidirectional
rlabel via2 s 1932 57 1988 113 6 VGND
port 2 nsew ground bidirectional
rlabel via2 s 1852 57 1908 113 6 VGND
port 2 nsew ground bidirectional
rlabel metal2 s 1843 57 1997 113 6 VGND
port 2 nsew ground bidirectional
rlabel via1 s 1926 61 1978 113 6 VGND
port 2 nsew ground bidirectional
rlabel via1 s 1862 61 1914 113 6 VGND
port 2 nsew ground bidirectional
rlabel metal1 s 0 51 1920 61 6 VGND
port 2 nsew ground bidirectional
rlabel metal1 s 0 61 1984 113 6 VGND
port 2 nsew ground bidirectional
rlabel metal1 s 0 113 1920 125 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 1867 76 1901 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 1795 76 1829 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 1591 76 1625 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 1519 76 1553 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 1447 76 1481 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 1278 76 1312 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 1206 76 1240 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 1134 76 1168 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 958 76 992 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 886 76 920 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 814 76 848 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 665 76 699 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 593 76 627 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 521 76 555 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 351 76 385 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 279 76 313 110 6 VGND
port 2 nsew ground bidirectional
rlabel viali s 207 76 241 110 6 VGND
port 2 nsew ground bidirectional
rlabel locali s 135 76 1901 110 6 VGND
port 2 nsew ground bidirectional
rlabel locali s 1795 110 1901 120 6 VGND
port 2 nsew ground bidirectional
rlabel locali s 1827 120 1901 289 6 VGND
port 2 nsew ground bidirectional
rlabel locali s 1433 110 1635 289 6 VGND
port 2 nsew ground bidirectional
rlabel locali s 1121 110 1323 289 6 VGND
port 2 nsew ground bidirectional
rlabel locali s 809 110 1011 289 6 VGND
port 2 nsew ground bidirectional
rlabel locali s 521 110 699 152 6 VGND
port 2 nsew ground bidirectional
rlabel locali s 553 152 699 289 6 VGND
port 2 nsew ground bidirectional
rlabel locali s 135 110 385 277 6 VGND
port 2 nsew ground bidirectional
rlabel metal1 s 0 -23 1920 23 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s -26 -43 1946 43 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 23 43 1901 317 6 VNB
port 3 nsew ground bidirectional
rlabel viali s 1855 -17 1889 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1759 -17 1793 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1663 -17 1697 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1567 -17 1601 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1471 -17 1505 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1375 -17 1409 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1279 -17 1313 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1183 -17 1217 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 1087 -17 1121 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 991 -17 1025 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 895 -17 929 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 799 -17 833 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 703 -17 737 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 607 -17 641 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 511 -17 545 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 415 -17 449 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 319 -17 353 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 223 -17 257 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 127 -17 161 17 8 VNB
port 3 nsew ground bidirectional
rlabel viali s 31 -17 65 17 8 VNB
port 3 nsew ground bidirectional
rlabel locali s 0 -17 1920 17 8 VNB
port 3 nsew ground bidirectional
rlabel metal1 s 0 791 1920 837 6 VPB
port 4 nsew power bidirectional
rlabel nwell s -66 377 1986 897 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1855 797 1889 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1759 797 1793 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1663 797 1697 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1567 797 1601 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1471 797 1505 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1375 797 1409 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1279 797 1313 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1183 797 1217 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 1087 797 1121 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 991 797 1025 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 895 797 929 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 799 797 833 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 703 797 737 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 607 797 641 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 511 797 545 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 415 797 449 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 319 797 353 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 223 797 257 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 127 797 161 831 6 VPB
port 4 nsew power bidirectional
rlabel viali s 31 797 65 831 6 VPB
port 4 nsew power bidirectional
rlabel locali s 0 797 1920 831 6 VPB
port 4 nsew power bidirectional
rlabel metal5 s 1582 567 2082 887 6 VPWR
port 5 nsew power bidirectional
rlabel metal4 s 1802 609 2038 845 6 VPWR
port 5 nsew power bidirectional
rlabel via3 s 1928 697 1992 761 6 VPWR
port 5 nsew power bidirectional
rlabel via3 s 1848 697 1912 761 6 VPWR
port 5 nsew power bidirectional
rlabel metal3 s 1842 696 1998 762 6 VPWR
port 5 nsew power bidirectional
rlabel via2 s 1932 701 1988 757 6 VPWR
port 5 nsew power bidirectional
rlabel via2 s 1852 701 1908 757 6 VPWR
port 5 nsew power bidirectional
rlabel metal2 s 1843 701 1997 757 6 VPWR
port 5 nsew power bidirectional
rlabel via1 s 1926 701 1978 753 6 VPWR
port 5 nsew power bidirectional
rlabel via1 s 1862 701 1914 753 6 VPWR
port 5 nsew power bidirectional
rlabel metal1 s 0 689 1920 701 6 VPWR
port 5 nsew power bidirectional
rlabel metal1 s 0 701 1984 753 6 VPWR
port 5 nsew power bidirectional
rlabel metal1 s 0 753 1920 763 6 VPWR
port 5 nsew power bidirectional
rlabel viali s 1853 695 1887 729 6 VPWR
port 5 nsew power bidirectional
rlabel viali s 1589 695 1623 729 6 VPWR
port 5 nsew power bidirectional
rlabel viali s 1446 695 1480 729 6 VPWR
port 5 nsew power bidirectional
rlabel viali s 1277 695 1311 729 6 VPWR
port 5 nsew power bidirectional
rlabel viali s 1205 695 1239 729 6 VPWR
port 5 nsew power bidirectional
rlabel viali s 1133 695 1167 729 6 VPWR
port 5 nsew power bidirectional
rlabel viali s 965 695 999 729 6 VPWR
port 5 nsew power bidirectional
rlabel viali s 893 695 927 729 6 VPWR
port 5 nsew power bidirectional
rlabel viali s 821 695 855 729 6 VPWR
port 5 nsew power bidirectional
rlabel viali s 626 695 660 729 6 VPWR
port 5 nsew power bidirectional
rlabel viali s 554 695 588 729 6 VPWR
port 5 nsew power bidirectional
rlabel viali s 339 695 373 729 6 VPWR
port 5 nsew power bidirectional
rlabel viali s 267 695 301 729 6 VPWR
port 5 nsew power bidirectional
rlabel viali s 195 695 229 729 6 VPWR
port 5 nsew power bidirectional
rlabel viali s 123 695 157 729 6 VPWR
port 5 nsew power bidirectional
rlabel locali s 1827 477 1901 695 6 VPWR
port 5 nsew power bidirectional
rlabel locali s 1781 695 1901 725 6 VPWR
port 5 nsew power bidirectional
rlabel locali s 1445 477 1623 725 6 VPWR
port 5 nsew power bidirectional
rlabel locali s 1133 477 1311 725 6 VPWR
port 5 nsew power bidirectional
rlabel locali s 821 477 999 725 6 VPWR
port 5 nsew power bidirectional
rlabel locali s 553 477 687 725 6 VPWR
port 5 nsew power bidirectional
rlabel locali s 123 489 373 725 6 VPWR
port 5 nsew power bidirectional
rlabel locali s 123 725 1901 759 6 VPWR
port 5 nsew power bidirectional
rlabel metal5 s 942 -73 1262 247 6 X
port 6 nsew signal output
rlabel metal5 s 458 247 1262 567 6 X
port 6 nsew signal output
rlabel metal5 s 942 567 1262 887 6 X
port 6 nsew signal output
rlabel metal4 s 1002 289 1238 525 6 X
port 6 nsew signal output
rlabel via3 s 1173 375 1237 439 6 X
port 6 nsew signal output
rlabel via3 s 1093 375 1157 439 6 X
port 6 nsew signal output
rlabel metal3 s 1087 374 1243 440 6 X
port 6 nsew signal output
rlabel metal4 s 482 289 718 525 6 X
port 6 nsew signal output
rlabel via2 s 1177 379 1233 435 6 X
port 6 nsew signal output
rlabel via2 s 1097 379 1153 435 6 X
port 6 nsew signal output
rlabel metal2 s 1088 379 1242 435 6 X
port 6 nsew signal output
rlabel via3 s 653 375 717 439 6 X
port 6 nsew signal output
rlabel via3 s 573 375 637 439 6 X
port 6 nsew signal output
rlabel metal3 s 567 375 723 439 6 X
port 6 nsew signal output
rlabel via1 s 1184 381 1236 433 6 X
port 6 nsew signal output
rlabel via1 s 1120 381 1172 433 6 X
port 6 nsew signal output
rlabel metal1 s 1112 381 1242 433 6 X
port 6 nsew signal output
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 1920 814
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_END 336350
string GDS_START 313384
<< end >>
