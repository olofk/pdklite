magic
tech sky130A
magscale 1 2
timestamp 1640697980
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 275 157 459 203
rect 1 21 459 157
rect 29 -17 63 21
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 17 416 138 527
rect 173 425 269 493
rect 303 418 354 527
rect 17 396 140 416
rect 103 391 140 396
rect 103 342 169 391
rect 388 353 443 493
rect 17 127 127 204
rect 229 158 295 243
rect 229 61 273 158
rect 409 147 443 353
rect 307 17 357 125
rect 391 51 443 147
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< obsli1 >>
rect 17 272 69 362
rect 203 327 354 377
rect 200 320 354 327
rect 197 318 354 320
rect 196 315 375 318
rect 192 312 375 315
rect 188 310 375 312
rect 183 308 375 310
rect 169 302 375 308
rect 165 296 375 302
rect 161 290 375 296
rect 155 285 375 290
rect 148 278 375 285
rect 142 277 375 278
rect 142 276 220 277
rect 142 274 215 276
rect 142 273 212 274
rect 142 272 209 273
rect 17 271 209 272
rect 17 269 207 271
rect 17 268 205 269
rect 17 266 203 268
rect 17 264 202 266
rect 17 263 201 264
rect 17 260 199 263
rect 17 257 198 260
rect 17 252 196 257
rect 17 238 195 252
rect 161 93 195 238
rect 17 59 195 93
rect 329 198 375 277
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 17 127 127 204 6 A
port 1 nsew signal input
rlabel locali s 173 425 269 493 6 B
port 2 nsew signal input
rlabel locali s 229 61 273 158 6 C
port 3 nsew signal input
rlabel locali s 229 158 295 243 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 460 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 397 -17 431 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 305 -17 339 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 213 -17 247 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 121 -17 155 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 29 -17 63 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 460 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 307 17 357 125 6 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 459 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 275 157 459 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 397 527 431 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 305 527 339 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 213 527 247 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 121 527 155 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 29 527 63 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 342 169 391 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 391 140 396 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 17 396 140 416 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 303 418 354 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 17 416 138 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 460 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 391 51 443 147 6 X
port 8 nsew signal output
rlabel locali s 409 147 443 353 6 X
port 8 nsew signal output
rlabel locali s 388 353 443 493 6 X
port 8 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3858454
string GDS_START 3851348
<< end >>
