magic
tech sky130A
magscale 1 2
timestamp 1640697995
<< nwell >>
rect -66 377 3426 897
<< pwell >>
rect 2641 283 2907 317
rect 545 217 1976 283
rect 2641 217 3356 283
rect 11 43 3356 217
rect -26 -43 3386 43
<< mvnmos >>
rect 94 107 194 191
rect 250 107 350 191
rect 628 173 728 257
rect 770 173 870 257
rect 926 173 1026 257
rect 1115 173 1215 257
rect 1257 173 1357 257
rect 1403 173 1503 257
rect 1644 107 1744 257
rect 1800 107 1900 257
rect 2014 107 2114 191
rect 2156 107 2256 191
rect 2312 107 2412 191
rect 2454 107 2554 191
rect 2724 141 2824 291
rect 2998 173 3098 257
rect 3177 107 3277 257
<< mvpmos >>
rect 94 533 194 683
rect 292 533 392 683
rect 566 608 666 692
rect 722 608 822 692
rect 878 608 978 692
rect 1034 608 1134 692
rect 1176 608 1276 692
rect 1332 608 1432 692
rect 1644 462 1744 662
rect 1800 462 1900 662
rect 1979 462 2079 546
rect 2122 462 2222 546
rect 2298 462 2398 546
rect 2454 462 2554 546
rect 2715 443 2815 743
rect 2994 443 3094 593
rect 3173 443 3273 743
<< mvndiff >>
rect 571 232 628 257
rect 571 198 583 232
rect 617 198 628 232
rect 37 166 94 191
rect 37 132 49 166
rect 83 132 94 166
rect 37 107 94 132
rect 194 166 250 191
rect 194 132 205 166
rect 239 132 250 166
rect 194 107 250 132
rect 350 166 407 191
rect 571 173 628 198
rect 728 173 770 257
rect 870 232 926 257
rect 870 198 881 232
rect 915 198 926 232
rect 870 173 926 198
rect 1026 232 1115 257
rect 1026 198 1070 232
rect 1104 198 1115 232
rect 1026 173 1115 198
rect 1215 173 1257 257
rect 1357 173 1403 257
rect 1503 173 1644 257
rect 350 132 361 166
rect 395 132 407 166
rect 1571 169 1644 173
rect 350 107 407 132
rect 1571 135 1583 169
rect 1617 135 1644 169
rect 1571 107 1644 135
rect 1744 249 1800 257
rect 1744 215 1755 249
rect 1789 215 1800 249
rect 1744 157 1800 215
rect 1744 123 1755 157
rect 1789 123 1800 157
rect 1744 107 1800 123
rect 1900 191 1950 257
rect 2667 283 2724 291
rect 2667 249 2679 283
rect 2713 249 2724 283
rect 1900 170 2014 191
rect 1900 136 1932 170
rect 1966 136 2014 170
rect 1900 107 2014 136
rect 2114 107 2156 191
rect 2256 152 2312 191
rect 2256 118 2267 152
rect 2301 118 2312 152
rect 2256 107 2312 118
rect 2412 107 2454 191
rect 2554 166 2607 191
rect 2554 132 2565 166
rect 2599 132 2607 166
rect 2667 183 2724 249
rect 2667 149 2679 183
rect 2713 149 2724 183
rect 2667 141 2724 149
rect 2824 283 2881 291
rect 2824 249 2835 283
rect 2869 249 2881 283
rect 2824 183 2881 249
rect 2824 149 2835 183
rect 2869 149 2881 183
rect 2941 232 2998 257
rect 2941 198 2953 232
rect 2987 198 2998 232
rect 2941 173 2998 198
rect 3098 249 3177 257
rect 3098 215 3132 249
rect 3166 215 3177 249
rect 3098 173 3177 215
rect 2824 141 2881 149
rect 3120 149 3177 173
rect 2554 107 2607 132
rect 3120 115 3132 149
rect 3166 115 3177 149
rect 3120 107 3177 115
rect 3277 245 3330 257
rect 3277 211 3288 245
rect 3322 211 3330 245
rect 3277 153 3330 211
rect 3277 119 3288 153
rect 3322 119 3330 153
rect 3277 107 3330 119
<< mvpdiff >>
rect 2658 735 2715 743
rect 2658 701 2670 735
rect 2704 701 2715 735
rect 37 675 94 683
rect 37 641 49 675
rect 83 641 94 675
rect 37 575 94 641
rect 37 541 49 575
rect 83 541 94 575
rect 37 533 94 541
rect 194 675 292 683
rect 194 641 205 675
rect 239 641 292 675
rect 194 575 292 641
rect 194 541 205 575
rect 239 541 292 575
rect 194 533 292 541
rect 392 675 449 683
rect 392 641 403 675
rect 437 641 449 675
rect 392 575 449 641
rect 509 667 566 692
rect 509 633 521 667
rect 555 633 566 667
rect 509 608 566 633
rect 666 667 722 692
rect 666 633 677 667
rect 711 633 722 667
rect 666 608 722 633
rect 822 667 878 692
rect 822 633 833 667
rect 867 633 878 667
rect 822 608 878 633
rect 978 667 1034 692
rect 978 633 989 667
rect 1023 633 1034 667
rect 978 608 1034 633
rect 1134 608 1176 692
rect 1276 681 1332 692
rect 1276 647 1287 681
rect 1321 647 1332 681
rect 1276 608 1332 647
rect 1432 662 1489 692
rect 1432 628 1443 662
rect 1477 628 1489 662
rect 1432 608 1489 628
rect 1587 649 1644 662
rect 1587 615 1599 649
rect 1633 615 1644 649
rect 392 541 403 575
rect 437 541 449 575
rect 392 533 449 541
rect 1587 462 1644 615
rect 1744 504 1800 662
rect 1744 470 1755 504
rect 1789 470 1800 504
rect 1744 462 1800 470
rect 1900 654 1957 662
rect 1900 620 1911 654
rect 1945 620 1957 654
rect 1900 579 1957 620
rect 1900 545 1911 579
rect 1945 546 1957 579
rect 2658 652 2715 701
rect 2658 618 2670 652
rect 2704 618 2715 652
rect 2658 568 2715 618
rect 2658 546 2670 568
rect 1945 545 1979 546
rect 1900 504 1979 545
rect 1900 470 1911 504
rect 1945 470 1979 504
rect 1900 462 1979 470
rect 2079 462 2122 546
rect 2222 521 2298 546
rect 2222 487 2233 521
rect 2267 487 2298 521
rect 2222 462 2298 487
rect 2398 521 2454 546
rect 2398 487 2409 521
rect 2443 487 2454 521
rect 2398 462 2454 487
rect 2554 534 2670 546
rect 2704 534 2715 568
rect 2554 485 2715 534
rect 2554 462 2670 485
rect 2658 451 2670 462
rect 2704 451 2715 485
rect 2658 443 2715 451
rect 2815 735 2872 743
rect 2815 701 2826 735
rect 2860 701 2872 735
rect 2815 652 2872 701
rect 2815 618 2826 652
rect 2860 618 2872 652
rect 3116 735 3173 743
rect 3116 701 3128 735
rect 3162 701 3173 735
rect 3116 652 3173 701
rect 2815 568 2872 618
rect 3116 618 3128 652
rect 3162 618 3173 652
rect 3116 593 3173 618
rect 2815 534 2826 568
rect 2860 534 2872 568
rect 2815 485 2872 534
rect 2815 451 2826 485
rect 2860 451 2872 485
rect 2815 443 2872 451
rect 2937 585 2994 593
rect 2937 551 2949 585
rect 2983 551 2994 585
rect 2937 485 2994 551
rect 2937 451 2949 485
rect 2983 451 2994 485
rect 2937 443 2994 451
rect 3094 568 3173 593
rect 3094 534 3128 568
rect 3162 534 3173 568
rect 3094 485 3173 534
rect 3094 451 3128 485
rect 3162 451 3173 485
rect 3094 443 3173 451
rect 3273 735 3330 743
rect 3273 701 3284 735
rect 3318 701 3330 735
rect 3273 652 3330 701
rect 3273 618 3284 652
rect 3318 618 3330 652
rect 3273 568 3330 618
rect 3273 534 3284 568
rect 3318 534 3330 568
rect 3273 485 3330 534
rect 3273 451 3284 485
rect 3318 451 3330 485
rect 3273 443 3330 451
<< mvndiffc >>
rect 583 198 617 232
rect 49 132 83 166
rect 205 132 239 166
rect 881 198 915 232
rect 1070 198 1104 232
rect 361 132 395 166
rect 1583 135 1617 169
rect 1755 215 1789 249
rect 1755 123 1789 157
rect 2679 249 2713 283
rect 1932 136 1966 170
rect 2267 118 2301 152
rect 2565 132 2599 166
rect 2679 149 2713 183
rect 2835 249 2869 283
rect 2835 149 2869 183
rect 2953 198 2987 232
rect 3132 215 3166 249
rect 3132 115 3166 149
rect 3288 211 3322 245
rect 3288 119 3322 153
<< mvpdiffc >>
rect 2670 701 2704 735
rect 49 641 83 675
rect 49 541 83 575
rect 205 641 239 675
rect 205 541 239 575
rect 403 641 437 675
rect 521 633 555 667
rect 677 633 711 667
rect 833 633 867 667
rect 989 633 1023 667
rect 1287 647 1321 681
rect 1443 628 1477 662
rect 1599 615 1633 649
rect 403 541 437 575
rect 1755 470 1789 504
rect 1911 620 1945 654
rect 1911 545 1945 579
rect 2670 618 2704 652
rect 1911 470 1945 504
rect 2233 487 2267 521
rect 2409 487 2443 521
rect 2670 534 2704 568
rect 2670 451 2704 485
rect 2826 701 2860 735
rect 2826 618 2860 652
rect 3128 701 3162 735
rect 3128 618 3162 652
rect 2826 534 2860 568
rect 2826 451 2860 485
rect 2949 551 2983 585
rect 2949 451 2983 485
rect 3128 534 3162 568
rect 3128 451 3162 485
rect 3284 701 3318 735
rect 3284 618 3318 652
rect 3284 534 3318 568
rect 3284 451 3318 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3360 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
<< poly >>
rect 2715 743 2815 769
rect 3173 743 3273 769
rect 94 683 194 709
rect 292 683 392 709
rect 566 692 666 718
rect 722 692 822 718
rect 878 692 978 718
rect 1034 692 1134 718
rect 1176 692 1276 718
rect 1332 692 1432 718
rect 1644 662 1744 688
rect 1800 662 1900 688
rect 94 341 194 533
rect 292 507 392 533
rect 94 307 135 341
rect 169 307 194 341
rect 94 273 194 307
rect 94 239 135 273
rect 169 239 194 273
rect 94 191 194 239
rect 250 485 392 507
rect 250 451 317 485
rect 351 451 392 485
rect 250 417 392 451
rect 250 383 317 417
rect 351 383 392 417
rect 250 363 392 383
rect 566 413 666 608
rect 722 527 822 608
rect 878 582 978 608
rect 878 548 992 582
rect 722 427 836 527
rect 566 379 612 413
rect 646 379 666 413
rect 770 405 836 427
rect 878 514 939 548
rect 973 514 992 548
rect 878 480 992 514
rect 878 446 939 480
rect 973 446 992 480
rect 878 426 992 446
rect 1034 560 1134 608
rect 1034 526 1080 560
rect 1114 526 1134 560
rect 1034 482 1134 526
rect 1176 582 1276 608
rect 1332 586 1432 608
rect 1176 487 1290 582
rect 1332 529 1503 586
rect 250 191 350 363
rect 566 345 728 379
rect 566 311 612 345
rect 646 311 728 345
rect 566 279 728 311
rect 628 257 728 279
rect 770 371 786 405
rect 820 383 836 405
rect 1034 383 1073 482
rect 1176 467 1361 487
rect 1176 466 1307 467
rect 1257 433 1307 466
rect 1341 433 1361 467
rect 820 371 870 383
rect 770 337 870 371
rect 770 303 786 337
rect 820 303 870 337
rect 770 257 870 303
rect 926 283 1073 383
rect 1115 404 1215 424
rect 1115 370 1135 404
rect 1169 370 1215 404
rect 1115 336 1215 370
rect 1115 302 1135 336
rect 1169 302 1215 336
rect 926 257 1026 283
rect 1115 257 1215 302
rect 1257 399 1361 433
rect 1257 365 1307 399
rect 1341 365 1361 399
rect 1257 283 1361 365
rect 1403 399 1503 529
rect 1979 546 2079 572
rect 2122 546 2222 572
rect 2298 546 2398 572
rect 2454 546 2554 572
rect 1403 365 1449 399
rect 1483 365 1503 399
rect 1644 379 1744 462
rect 1257 257 1357 283
rect 1403 257 1503 365
rect 1563 329 1744 379
rect 1800 414 1900 462
rect 1979 440 2079 462
rect 1800 380 1841 414
rect 1875 380 1900 414
rect 1800 360 1900 380
rect 1942 402 2079 440
rect 1942 368 1962 402
rect 1996 368 2079 402
rect 1563 295 1583 329
rect 1617 295 1744 329
rect 1942 348 2079 368
rect 2122 440 2222 462
rect 2122 364 2256 440
rect 2122 348 2202 364
rect 1942 318 1972 348
rect 1563 279 1744 295
rect 1644 257 1744 279
rect 1800 279 1972 318
rect 2156 330 2202 348
rect 2236 330 2256 364
rect 1800 257 1900 279
rect 2014 264 2114 306
rect 628 147 728 173
rect 770 147 870 173
rect 926 147 1026 173
rect 1115 147 1215 173
rect 1257 147 1357 173
rect 1403 147 1503 173
rect 2014 230 2034 264
rect 2068 230 2114 264
rect 2014 191 2114 230
rect 2156 296 2256 330
rect 2156 262 2202 296
rect 2236 262 2256 296
rect 2156 191 2256 262
rect 2298 305 2398 462
rect 2454 440 2554 462
rect 2994 593 3094 619
rect 2440 417 2554 440
rect 2715 417 2815 443
rect 2994 417 3094 443
rect 2440 414 3098 417
rect 2440 380 2456 414
rect 2490 380 3098 414
rect 3173 383 3273 443
rect 2440 347 3098 380
rect 2454 317 3098 347
rect 2298 267 2412 305
rect 2298 233 2318 267
rect 2352 233 2412 267
rect 2298 213 2412 233
rect 2312 191 2412 213
rect 2454 191 2554 317
rect 2724 291 2824 317
rect 2994 283 3098 317
rect 3162 351 3277 383
rect 3162 317 3182 351
rect 3216 317 3277 351
rect 3162 283 3277 317
rect 2998 257 3098 283
rect 3177 257 3277 283
rect 2998 147 3098 173
rect 2724 115 2824 141
rect 94 81 194 107
rect 250 81 350 107
rect 1644 81 1744 107
rect 1800 81 1900 107
rect 2014 81 2114 107
rect 2156 81 2256 107
rect 2312 81 2412 107
rect 2454 81 2554 107
rect 3177 81 3277 107
<< polycont >>
rect 135 307 169 341
rect 135 239 169 273
rect 317 451 351 485
rect 317 383 351 417
rect 612 379 646 413
rect 939 514 973 548
rect 939 446 973 480
rect 1080 526 1114 560
rect 612 311 646 345
rect 786 371 820 405
rect 1307 433 1341 467
rect 786 303 820 337
rect 1135 370 1169 404
rect 1135 302 1169 336
rect 1307 365 1341 399
rect 1449 365 1483 399
rect 1841 380 1875 414
rect 1962 368 1996 402
rect 1583 295 1617 329
rect 2202 330 2236 364
rect 2034 230 2068 264
rect 2202 262 2236 296
rect 2456 380 2490 414
rect 2318 233 2352 267
rect 3182 317 3216 351
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3360 831
rect 119 735 297 741
rect 153 701 191 735
rect 225 701 263 735
rect 33 675 83 691
rect 33 641 49 675
rect 33 575 83 641
rect 33 541 49 575
rect 33 489 83 541
rect 119 675 297 701
rect 119 641 205 675
rect 239 641 297 675
rect 119 575 297 641
rect 119 541 205 575
rect 239 541 297 575
rect 119 525 297 541
rect 333 727 641 761
rect 333 489 367 727
rect 33 485 367 489
rect 33 455 317 485
rect 33 199 83 455
rect 301 451 317 455
rect 351 451 367 485
rect 301 417 367 451
rect 301 383 317 417
rect 351 383 367 417
rect 301 380 367 383
rect 403 675 455 691
rect 437 641 455 675
rect 403 575 455 641
rect 437 541 455 575
rect 403 350 455 541
rect 505 667 571 684
rect 505 633 521 667
rect 555 633 571 667
rect 505 494 571 633
rect 607 564 641 727
rect 677 735 711 741
rect 677 667 711 701
rect 677 600 711 633
rect 747 720 1113 754
rect 747 564 781 720
rect 817 667 903 684
rect 817 633 833 667
rect 867 633 903 667
rect 817 600 903 633
rect 973 667 1043 684
rect 973 633 989 667
rect 1023 633 1043 667
rect 973 600 1043 633
rect 607 530 781 564
rect 869 494 903 600
rect 505 460 903 494
rect 119 341 185 344
rect 119 307 135 341
rect 169 307 185 341
rect 119 273 185 307
rect 119 239 135 273
rect 169 239 185 273
rect 119 235 185 239
rect 403 316 415 350
rect 449 316 455 350
rect 403 310 455 316
rect 596 413 733 424
rect 596 379 612 413
rect 646 379 733 413
rect 596 345 733 379
rect 596 311 612 345
rect 646 311 733 345
rect 403 199 437 310
rect 596 301 733 311
rect 33 166 99 199
rect 33 132 49 166
rect 83 132 99 166
rect 33 99 99 132
rect 135 166 325 199
rect 135 132 205 166
rect 239 132 325 166
rect 135 113 325 132
rect 135 79 141 113
rect 175 79 213 113
rect 247 79 285 113
rect 319 79 325 113
rect 361 166 437 199
rect 395 132 437 166
rect 361 99 437 132
rect 473 232 663 265
rect 473 198 583 232
rect 617 198 663 232
rect 473 113 663 198
rect 135 73 325 79
rect 473 79 479 113
rect 513 79 551 113
rect 585 79 623 113
rect 657 79 663 113
rect 699 126 733 301
rect 770 405 833 421
rect 770 371 786 405
rect 820 371 833 405
rect 770 337 833 371
rect 770 303 786 337
rect 820 303 833 337
rect 770 162 833 303
rect 869 265 903 460
rect 939 548 973 564
rect 939 480 973 514
rect 939 356 973 446
rect 1009 474 1043 600
rect 1079 609 1113 720
rect 1149 735 1337 741
rect 1149 701 1154 735
rect 1188 701 1226 735
rect 1260 701 1298 735
rect 1332 701 1337 735
rect 1149 681 1337 701
rect 1149 647 1287 681
rect 1321 647 1337 681
rect 1149 645 1337 647
rect 1373 727 1547 761
rect 1373 609 1407 727
rect 1079 575 1407 609
rect 1443 662 1477 691
rect 1079 560 1130 575
rect 1079 526 1080 560
rect 1114 526 1130 560
rect 1443 539 1477 628
rect 1513 574 1547 727
rect 1583 735 1773 741
rect 1583 701 1589 735
rect 1623 701 1661 735
rect 1695 701 1733 735
rect 1767 701 1773 735
rect 1583 649 1773 701
rect 2118 735 2308 741
rect 2118 701 2124 735
rect 2158 701 2196 735
rect 2230 701 2268 735
rect 2302 701 2308 735
rect 1583 615 1599 649
rect 1633 615 1773 649
rect 1583 610 1773 615
rect 1911 654 1961 670
rect 1945 620 1961 654
rect 1911 579 1961 620
rect 1513 540 1875 574
rect 1079 510 1130 526
rect 1221 505 1477 539
rect 1221 474 1255 505
rect 1009 440 1255 474
rect 1739 470 1755 504
rect 1789 470 1805 504
rect 1739 469 1805 470
rect 1119 370 1135 404
rect 1169 370 1185 404
rect 1119 356 1185 370
rect 939 350 1185 356
rect 939 316 991 350
rect 1025 336 1185 350
rect 1025 316 1135 336
rect 939 302 1135 316
rect 1169 302 1185 336
rect 939 301 1185 302
rect 1221 329 1255 440
rect 1291 467 1805 469
rect 1291 433 1307 467
rect 1341 435 1805 467
rect 1341 433 1357 435
rect 1291 399 1357 433
rect 1291 365 1307 399
rect 1341 365 1357 399
rect 1433 365 1449 399
rect 1483 365 1703 399
rect 1221 295 1583 329
rect 1617 295 1633 329
rect 1221 265 1255 295
rect 869 232 931 265
rect 869 198 881 232
rect 915 198 931 232
rect 869 165 931 198
rect 1054 232 1255 265
rect 1669 259 1703 365
rect 1054 198 1070 232
rect 1104 231 1255 232
rect 1104 198 1120 231
rect 1054 165 1120 198
rect 1291 225 1703 259
rect 1291 126 1325 225
rect 699 92 1325 126
rect 1443 169 1633 189
rect 1443 135 1583 169
rect 1617 135 1633 169
rect 1443 113 1633 135
rect 473 73 663 79
rect 1443 79 1449 113
rect 1483 79 1521 113
rect 1555 79 1593 113
rect 1627 79 1633 113
rect 1443 73 1633 79
rect 1669 87 1703 225
rect 1739 249 1805 435
rect 1739 215 1755 249
rect 1789 215 1805 249
rect 1841 414 1875 540
rect 1945 545 1961 579
rect 1911 504 1961 545
rect 1945 488 1961 504
rect 2118 521 2308 701
rect 2612 735 2790 751
rect 2646 701 2670 735
rect 2718 701 2756 735
rect 2612 652 2790 701
rect 2612 618 2670 652
rect 2704 618 2790 652
rect 2612 568 2790 618
rect 1945 470 2082 488
rect 2118 487 2233 521
rect 2267 487 2308 521
rect 2118 470 2308 487
rect 2393 521 2459 554
rect 2393 487 2409 521
rect 2443 504 2459 521
rect 2612 534 2670 568
rect 2704 534 2790 568
rect 2443 487 2576 504
rect 2393 470 2576 487
rect 1911 454 2082 470
rect 2048 434 2082 454
rect 1841 280 1875 380
rect 1945 402 2012 418
rect 1945 368 1962 402
rect 1996 368 2012 402
rect 2048 414 2506 434
rect 2048 400 2456 414
rect 1945 350 2012 368
rect 1945 316 1951 350
rect 1985 316 2012 350
rect 1841 264 2075 280
rect 1841 246 2034 264
rect 1739 157 1805 215
rect 2018 230 2034 246
rect 2068 230 2075 264
rect 2018 214 2075 230
rect 1739 123 1755 157
rect 1789 123 1805 157
rect 1916 170 1982 199
rect 1916 136 1932 170
rect 1966 157 1982 170
rect 2111 157 2145 400
rect 2440 380 2456 400
rect 2490 380 2506 414
rect 2440 376 2506 380
rect 2186 330 2202 364
rect 2236 340 2252 364
rect 2542 340 2576 470
rect 2612 485 2790 534
rect 2612 451 2670 485
rect 2704 451 2790 485
rect 2612 435 2790 451
rect 2826 735 2876 751
rect 2860 701 2876 735
rect 2826 652 2876 701
rect 2860 618 2876 652
rect 2826 568 2876 618
rect 3035 735 3225 751
rect 3035 701 3041 735
rect 3075 701 3113 735
rect 3162 701 3185 735
rect 3219 701 3225 735
rect 3035 652 3225 701
rect 3035 618 3128 652
rect 3162 618 3225 652
rect 2860 534 2876 568
rect 2826 485 2876 534
rect 2860 451 2876 485
rect 2826 356 2876 451
rect 2236 330 2576 340
rect 2186 306 2576 330
rect 2186 296 2252 306
rect 2186 262 2202 296
rect 2236 262 2252 296
rect 2302 267 2368 270
rect 2302 233 2318 267
rect 2352 233 2368 267
rect 2302 226 2368 233
rect 1966 136 2145 157
rect 1916 123 2145 136
rect 2181 192 2368 226
rect 2542 195 2576 306
rect 2809 299 2876 356
rect 2933 585 2999 601
rect 2933 551 2949 585
rect 2983 551 2999 585
rect 2933 485 2999 551
rect 2933 451 2949 485
rect 2983 451 2999 485
rect 2933 367 2999 451
rect 3035 568 3225 618
rect 3035 534 3128 568
rect 3162 534 3225 568
rect 3035 485 3225 534
rect 3035 451 3128 485
rect 3162 451 3225 485
rect 3035 435 3225 451
rect 3268 735 3338 751
rect 3268 701 3284 735
rect 3318 701 3338 735
rect 3268 652 3338 701
rect 3268 618 3284 652
rect 3318 618 3338 652
rect 3268 568 3338 618
rect 3268 534 3284 568
rect 3318 534 3338 568
rect 3268 485 3338 534
rect 3268 451 3284 485
rect 3318 451 3338 485
rect 2933 351 3232 367
rect 2933 317 3182 351
rect 3216 317 3232 351
rect 2933 301 3232 317
rect 2651 283 2769 299
rect 2651 249 2679 283
rect 2713 249 2769 283
rect 2181 87 2215 192
rect 2542 166 2615 195
rect 1669 53 2215 87
rect 2251 152 2441 156
rect 2251 118 2267 152
rect 2301 118 2441 152
rect 2251 113 2441 118
rect 2251 79 2257 113
rect 2291 79 2329 113
rect 2363 79 2401 113
rect 2435 79 2441 113
rect 2542 132 2565 166
rect 2599 132 2615 166
rect 2542 103 2615 132
rect 2651 183 2769 249
rect 2651 149 2679 183
rect 2713 149 2769 183
rect 2651 113 2769 149
rect 2809 283 2885 299
rect 2809 249 2835 283
rect 2869 249 2885 283
rect 2809 183 2885 249
rect 2809 149 2835 183
rect 2869 149 2885 183
rect 2933 232 3003 301
rect 2933 198 2953 232
rect 2987 198 3003 232
rect 2933 165 3003 198
rect 3039 249 3229 265
rect 3039 215 3132 249
rect 3166 215 3229 249
rect 2809 133 2885 149
rect 3039 149 3229 215
rect 2251 73 2441 79
rect 2651 79 2657 113
rect 2691 79 2729 113
rect 2763 79 2769 113
rect 2651 73 2769 79
rect 3039 115 3132 149
rect 3166 115 3229 149
rect 3039 113 3229 115
rect 3039 79 3045 113
rect 3079 79 3117 113
rect 3151 79 3189 113
rect 3223 79 3229 113
rect 3268 245 3338 451
rect 3268 211 3288 245
rect 3322 211 3338 245
rect 3268 153 3338 211
rect 3268 119 3288 153
rect 3322 119 3338 153
rect 3268 103 3338 119
rect 3039 73 3229 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 119 701 153 735
rect 191 701 225 735
rect 263 701 297 735
rect 677 701 711 735
rect 415 316 449 350
rect 141 79 175 113
rect 213 79 247 113
rect 285 79 319 113
rect 479 79 513 113
rect 551 79 585 113
rect 623 79 657 113
rect 1154 701 1188 735
rect 1226 701 1260 735
rect 1298 701 1332 735
rect 1589 701 1623 735
rect 1661 701 1695 735
rect 1733 701 1767 735
rect 2124 701 2158 735
rect 2196 701 2230 735
rect 2268 701 2302 735
rect 991 316 1025 350
rect 1449 79 1483 113
rect 1521 79 1555 113
rect 1593 79 1627 113
rect 2612 701 2646 735
rect 2684 701 2704 735
rect 2704 701 2718 735
rect 2756 701 2790 735
rect 1951 316 1985 350
rect 3041 701 3075 735
rect 3113 701 3128 735
rect 3128 701 3147 735
rect 3185 701 3219 735
rect 2257 79 2291 113
rect 2329 79 2363 113
rect 2401 79 2435 113
rect 2657 79 2691 113
rect 2729 79 2763 113
rect 3045 79 3079 113
rect 3117 79 3151 113
rect 3189 79 3223 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
<< metal1 >>
rect 0 831 3360 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3360 831
rect 0 791 3360 797
rect 0 735 3360 763
rect 0 701 119 735
rect 153 701 191 735
rect 225 701 263 735
rect 297 701 677 735
rect 711 701 1154 735
rect 1188 701 1226 735
rect 1260 701 1298 735
rect 1332 701 1589 735
rect 1623 701 1661 735
rect 1695 701 1733 735
rect 1767 701 2124 735
rect 2158 701 2196 735
rect 2230 701 2268 735
rect 2302 701 2612 735
rect 2646 701 2684 735
rect 2718 701 2756 735
rect 2790 701 3041 735
rect 3075 701 3113 735
rect 3147 701 3185 735
rect 3219 701 3360 735
rect 0 689 3360 701
rect 403 350 461 356
rect 403 316 415 350
rect 449 347 461 350
rect 979 350 1037 356
rect 979 347 991 350
rect 449 319 991 347
rect 449 316 461 319
rect 403 310 461 316
rect 979 316 991 319
rect 1025 347 1037 350
rect 1939 350 1997 356
rect 1939 347 1951 350
rect 1025 319 1951 347
rect 1025 316 1037 319
rect 979 310 1037 316
rect 1939 316 1951 319
rect 1985 316 1997 350
rect 1939 310 1997 316
rect 0 113 3360 125
rect 0 79 141 113
rect 175 79 213 113
rect 247 79 285 113
rect 319 79 479 113
rect 513 79 551 113
rect 585 79 623 113
rect 657 79 1449 113
rect 1483 79 1521 113
rect 1555 79 1593 113
rect 1627 79 2257 113
rect 2291 79 2329 113
rect 2363 79 2401 113
rect 2435 79 2657 113
rect 2691 79 2729 113
rect 2763 79 3045 113
rect 3079 79 3117 113
rect 3151 79 3189 113
rect 3223 79 3360 113
rect 0 51 3360 79
rect 0 17 3360 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
rect 0 -23 3360 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfrbp_1
flabel metal1 s 0 51 3360 125 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 0 3360 23 0 FreeSans 340 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 0 689 3360 763 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 791 3360 814 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 3295 168 3329 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3295 242 3329 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3295 316 3329 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3295 390 3329 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3295 464 3329 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3295 538 3329 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3295 612 3329 646 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2815 168 2849 202 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2815 242 2849 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2815 316 2849 350 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 3360 814
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string LEFsymmetry X Y
string GDS_END 1031540
string GDS_START 1000276
<< end >>
