magic
tech sky130A
magscale 1 2
timestamp 1619729571
<< checkpaint >>
rect -1298 -1308 3690 1852
<< nwell >>
rect -38 261 2430 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 423 47 453 131
rect 611 47 641 131
rect 699 47 729 131
rect 801 47 831 131
rect 983 47 1013 119
rect 1071 47 1101 119
rect 1177 47 1207 131
rect 1296 47 1326 175
rect 1484 47 1514 131
rect 1581 47 1611 119
rect 1687 47 1717 119
rect 1782 47 1812 131
rect 1879 47 1909 177
rect 2122 47 2152 131
rect 2219 47 2249 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 423 369 453 497
rect 611 369 641 497
rect 699 369 729 497
rect 801 369 831 497
rect 956 413 986 497
rect 1047 413 1077 497
rect 1150 413 1180 497
rect 1282 347 1312 497
rect 1470 413 1500 497
rect 1561 413 1591 497
rect 1645 413 1675 497
rect 1759 413 1789 497
rect 1856 297 1886 497
rect 2122 369 2152 497
rect 2219 297 2249 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 100 351 131
rect 299 66 307 100
rect 341 66 351 100
rect 299 47 351 66
rect 381 47 423 131
rect 453 93 505 131
rect 453 59 463 93
rect 497 59 505 93
rect 453 47 505 59
rect 559 119 611 131
rect 559 85 567 119
rect 601 85 611 119
rect 559 47 611 85
rect 641 106 699 131
rect 641 72 653 106
rect 687 72 699 106
rect 641 47 699 72
rect 729 47 801 131
rect 831 119 883 131
rect 1246 131 1296 175
rect 1127 119 1177 131
rect 831 106 983 119
rect 831 72 841 106
rect 875 72 983 106
rect 831 47 983 72
rect 1013 99 1071 119
rect 1013 65 1023 99
rect 1057 65 1071 99
rect 1013 47 1071 65
rect 1101 47 1177 119
rect 1207 101 1296 131
rect 1207 67 1218 101
rect 1252 67 1296 101
rect 1207 47 1296 67
rect 1326 163 1378 175
rect 1326 129 1336 163
rect 1370 129 1378 163
rect 1326 95 1378 129
rect 1326 61 1336 95
rect 1370 61 1378 95
rect 1326 47 1378 61
rect 1432 107 1484 131
rect 1432 73 1440 107
rect 1474 73 1484 107
rect 1432 47 1484 73
rect 1514 119 1564 131
rect 1827 164 1879 177
rect 1827 131 1835 164
rect 1732 119 1782 131
rect 1514 47 1581 119
rect 1611 104 1687 119
rect 1611 70 1624 104
rect 1658 70 1687 104
rect 1611 47 1687 70
rect 1717 47 1782 119
rect 1812 130 1835 131
rect 1869 130 1879 164
rect 1812 96 1879 130
rect 1812 62 1835 96
rect 1869 62 1879 96
rect 1812 47 1879 62
rect 1909 164 1961 177
rect 1909 130 1919 164
rect 1953 130 1961 164
rect 2167 164 2219 177
rect 2167 131 2175 164
rect 1909 96 1961 130
rect 1909 62 1919 96
rect 1953 62 1961 96
rect 1909 47 1961 62
rect 2070 94 2122 131
rect 2070 60 2078 94
rect 2112 60 2122 94
rect 2070 47 2122 60
rect 2152 130 2175 131
rect 2209 130 2219 164
rect 2152 96 2219 130
rect 2152 62 2175 96
rect 2209 62 2219 96
rect 2152 47 2219 62
rect 2249 164 2305 177
rect 2249 130 2261 164
rect 2295 130 2305 164
rect 2249 96 2305 130
rect 2249 62 2261 96
rect 2295 62 2305 96
rect 2249 47 2305 62
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 485 351 497
rect 299 451 307 485
rect 341 451 351 485
rect 299 415 351 451
rect 299 381 307 415
rect 341 381 351 415
rect 299 369 351 381
rect 381 369 423 497
rect 453 485 505 497
rect 453 451 463 485
rect 497 451 505 485
rect 453 417 505 451
rect 453 383 463 417
rect 497 383 505 417
rect 453 369 505 383
rect 559 485 611 497
rect 559 451 567 485
rect 601 451 611 485
rect 559 415 611 451
rect 559 381 567 415
rect 601 381 611 415
rect 559 369 611 381
rect 641 485 699 497
rect 641 451 653 485
rect 687 451 699 485
rect 641 415 699 451
rect 641 381 653 415
rect 687 381 699 415
rect 641 369 699 381
rect 729 369 801 497
rect 831 485 956 497
rect 831 451 841 485
rect 875 451 956 485
rect 831 417 956 451
rect 831 383 841 417
rect 875 413 956 417
rect 986 472 1047 497
rect 986 438 999 472
rect 1033 438 1047 472
rect 986 413 1047 438
rect 1077 413 1150 497
rect 1180 485 1282 497
rect 1180 451 1232 485
rect 1266 451 1282 485
rect 1180 417 1282 451
rect 1180 413 1232 417
rect 875 383 883 413
rect 831 369 883 383
rect 1195 383 1232 413
rect 1266 383 1282 417
rect 1195 347 1282 383
rect 1312 485 1364 497
rect 1312 451 1322 485
rect 1356 451 1364 485
rect 1312 393 1364 451
rect 1418 472 1470 497
rect 1418 438 1426 472
rect 1460 438 1470 472
rect 1418 413 1470 438
rect 1500 413 1561 497
rect 1591 469 1645 497
rect 1591 435 1601 469
rect 1635 435 1645 469
rect 1591 413 1645 435
rect 1675 413 1759 497
rect 1789 485 1856 497
rect 1789 451 1812 485
rect 1846 451 1856 485
rect 1789 417 1856 451
rect 1789 413 1812 417
rect 1312 359 1322 393
rect 1356 359 1364 393
rect 1312 347 1364 359
rect 1804 383 1812 413
rect 1846 383 1856 417
rect 1804 349 1856 383
rect 1804 315 1812 349
rect 1846 315 1856 349
rect 1804 297 1856 315
rect 1886 479 1938 497
rect 1886 445 1896 479
rect 1930 445 1938 479
rect 1886 411 1938 445
rect 1886 377 1896 411
rect 1930 377 1938 411
rect 2068 485 2122 497
rect 2068 451 2076 485
rect 2110 451 2122 485
rect 2068 415 2122 451
rect 2068 381 2076 415
rect 2110 381 2122 415
rect 1886 343 1938 377
rect 1886 309 1896 343
rect 1930 309 1938 343
rect 1886 297 1938 309
rect 2068 369 2122 381
rect 2152 479 2219 497
rect 2152 445 2175 479
rect 2209 445 2219 479
rect 2152 411 2219 445
rect 2152 377 2175 411
rect 2209 377 2219 411
rect 2152 369 2219 377
rect 2167 343 2219 369
rect 2167 309 2175 343
rect 2209 309 2219 343
rect 2167 297 2219 309
rect 2249 479 2305 497
rect 2249 445 2261 479
rect 2295 445 2305 479
rect 2249 411 2305 445
rect 2249 377 2261 411
rect 2295 377 2305 411
rect 2249 343 2305 377
rect 2249 309 2261 343
rect 2295 309 2305 343
rect 2249 297 2305 309
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 66 341 100
rect 463 59 497 93
rect 567 85 601 119
rect 653 72 687 106
rect 841 72 875 106
rect 1023 65 1057 99
rect 1218 67 1252 101
rect 1336 129 1370 163
rect 1336 61 1370 95
rect 1440 73 1474 107
rect 1624 70 1658 104
rect 1835 130 1869 164
rect 1835 62 1869 96
rect 1919 130 1953 164
rect 1919 62 1953 96
rect 2078 60 2112 94
rect 2175 130 2209 164
rect 2175 62 2209 96
rect 2261 130 2295 164
rect 2261 62 2295 96
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 451 341 485
rect 307 381 341 415
rect 463 451 497 485
rect 463 383 497 417
rect 567 451 601 485
rect 567 381 601 415
rect 653 451 687 485
rect 653 381 687 415
rect 841 451 875 485
rect 841 383 875 417
rect 999 438 1033 472
rect 1232 451 1266 485
rect 1232 383 1266 417
rect 1322 451 1356 485
rect 1426 438 1460 472
rect 1601 435 1635 469
rect 1812 451 1846 485
rect 1322 359 1356 393
rect 1812 383 1846 417
rect 1812 315 1846 349
rect 1896 445 1930 479
rect 1896 377 1930 411
rect 2076 451 2110 485
rect 2076 381 2110 415
rect 1896 309 1930 343
rect 2175 445 2209 479
rect 2175 377 2209 411
rect 2175 309 2209 343
rect 2261 445 2295 479
rect 2261 377 2295 411
rect 2261 309 2295 343
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 423 497 453 523
rect 611 497 641 523
rect 699 497 729 523
rect 801 497 831 523
rect 956 497 986 523
rect 1047 497 1077 523
rect 1150 497 1180 523
rect 1282 497 1312 523
rect 1470 497 1500 523
rect 1561 497 1591 523
rect 1645 497 1675 523
rect 1759 497 1789 523
rect 1856 497 1886 523
rect 2122 497 2152 523
rect 2219 497 2249 523
rect 79 348 109 363
rect 47 318 109 348
rect 47 265 77 318
rect 163 274 193 363
rect 351 330 381 369
rect 423 354 453 369
rect 423 343 549 354
rect 23 249 77 265
rect 23 215 33 249
rect 67 215 77 249
rect 119 264 193 274
rect 119 230 135 264
rect 169 230 193 264
rect 119 220 193 230
rect 23 199 77 215
rect 47 176 77 199
rect 47 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 323 314 383 330
rect 425 324 549 343
rect 323 280 339 314
rect 373 280 383 314
rect 323 246 383 280
rect 483 321 549 324
rect 483 287 499 321
rect 533 287 549 321
rect 483 277 549 287
rect 611 322 641 369
rect 699 322 729 369
rect 801 330 831 369
rect 611 292 729 322
rect 791 314 845 330
rect 323 212 339 246
rect 373 212 383 246
rect 323 196 383 212
rect 425 219 491 235
rect 351 131 381 196
rect 425 185 441 219
rect 475 200 491 219
rect 611 200 641 292
rect 791 280 801 314
rect 835 280 845 314
rect 956 297 986 413
rect 1047 381 1077 413
rect 1047 365 1108 381
rect 1047 331 1064 365
rect 1098 331 1108 365
rect 1047 315 1108 331
rect 791 264 845 280
rect 943 287 1009 297
rect 475 185 641 200
rect 425 176 641 185
rect 423 170 641 176
rect 423 162 491 170
rect 423 131 453 162
rect 611 131 641 170
rect 683 219 737 235
rect 683 185 693 219
rect 727 185 737 219
rect 683 169 737 185
rect 699 131 729 169
rect 801 131 831 264
rect 943 253 959 287
rect 993 273 1009 287
rect 993 253 1101 273
rect 943 243 1101 253
rect 963 191 1029 201
rect 963 157 979 191
rect 1013 157 1029 191
rect 963 147 1029 157
rect 983 119 1013 147
rect 1071 119 1101 243
rect 1150 213 1180 413
rect 1282 309 1312 347
rect 1222 299 1312 309
rect 1222 265 1238 299
rect 1272 265 1312 299
rect 1470 275 1500 413
rect 1561 315 1591 413
rect 1645 375 1675 413
rect 1644 365 1710 375
rect 1644 331 1660 365
rect 1694 331 1710 365
rect 1644 321 1710 331
rect 1222 255 1312 265
rect 1282 220 1312 255
rect 1445 259 1500 275
rect 1445 225 1455 259
rect 1489 225 1500 259
rect 1548 299 1602 315
rect 1548 265 1558 299
rect 1592 279 1602 299
rect 1592 265 1717 279
rect 1548 249 1717 265
rect 1150 203 1224 213
rect 1150 169 1174 203
rect 1208 169 1224 203
rect 1282 190 1326 220
rect 1296 175 1326 190
rect 1445 209 1500 225
rect 1445 179 1514 209
rect 1150 159 1224 169
rect 1177 131 1207 159
rect 1484 131 1514 179
rect 1581 191 1645 207
rect 1581 157 1601 191
rect 1635 157 1645 191
rect 1581 141 1645 157
rect 1581 119 1611 141
rect 1687 119 1717 249
rect 1759 244 1789 413
rect 1976 365 2030 381
rect 1976 331 1986 365
rect 2020 331 2030 365
rect 2122 331 2152 369
rect 1856 244 1886 297
rect 1976 286 2152 331
rect 2122 265 2152 286
rect 2219 265 2249 297
rect 1759 228 2047 244
rect 1759 207 2003 228
rect 1782 131 1812 207
rect 1879 177 1909 207
rect 1993 194 2003 207
rect 2037 194 2047 228
rect 1993 178 2047 194
rect 2122 199 2249 265
rect 2122 131 2152 199
rect 2219 177 2249 199
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 423 21 453 47
rect 611 21 641 47
rect 699 21 729 47
rect 801 21 831 47
rect 983 21 1013 47
rect 1071 21 1101 47
rect 1177 21 1207 47
rect 1296 21 1326 47
rect 1484 21 1514 47
rect 1581 21 1611 47
rect 1687 21 1717 47
rect 1782 21 1812 47
rect 1879 21 1909 47
rect 2122 21 2152 47
rect 2219 21 2249 47
<< polycont >>
rect 33 215 67 249
rect 135 230 169 264
rect 339 280 373 314
rect 499 287 533 321
rect 339 212 373 246
rect 441 185 475 219
rect 801 280 835 314
rect 1064 331 1098 365
rect 693 185 727 219
rect 959 253 993 287
rect 979 157 1013 191
rect 1238 265 1272 299
rect 1660 331 1694 365
rect 1455 225 1489 259
rect 1558 265 1592 299
rect 1174 169 1208 203
rect 1601 157 1635 191
rect 1986 331 2020 365
rect 2003 194 2037 228
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 237 493
rect 203 409 237 443
rect 69 391 169 393
rect 69 375 127 391
rect 35 359 127 375
rect 123 357 127 359
rect 161 357 169 391
rect 19 249 89 325
rect 19 215 33 249
rect 67 215 89 249
rect 19 195 89 215
rect 123 264 169 357
rect 123 230 135 264
rect 123 161 169 230
rect 35 127 169 161
rect 203 323 237 375
rect 35 119 69 127
rect 203 119 237 289
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 271 485 357 493
rect 271 451 307 485
rect 341 451 357 485
rect 271 415 357 451
rect 271 381 307 415
rect 341 381 357 415
rect 271 378 357 381
rect 447 485 513 527
rect 653 485 692 527
rect 447 451 463 485
rect 497 451 513 485
rect 447 417 513 451
rect 447 383 463 417
rect 497 383 513 417
rect 447 378 513 383
rect 551 451 567 485
rect 601 451 617 485
rect 551 415 617 451
rect 551 381 567 415
rect 601 381 617 415
rect 271 119 305 378
rect 551 344 617 381
rect 687 451 692 485
rect 653 415 692 451
rect 687 381 692 415
rect 653 365 692 381
rect 825 485 891 493
rect 825 451 841 485
rect 875 451 891 485
rect 1225 485 1272 527
rect 825 417 891 451
rect 983 472 1191 475
rect 983 438 999 472
rect 1033 438 1191 472
rect 983 435 1191 438
rect 825 383 841 417
rect 875 404 891 417
rect 875 383 903 404
rect 825 364 903 383
rect 339 314 383 344
rect 373 280 383 314
rect 339 246 383 280
rect 499 321 617 344
rect 533 287 617 321
rect 373 212 383 246
rect 339 153 383 212
rect 422 237 465 274
rect 499 271 617 287
rect 422 219 513 237
rect 422 185 441 219
rect 475 185 513 219
rect 422 153 513 185
rect 556 235 617 271
rect 761 314 835 330
rect 761 280 801 314
rect 761 264 835 280
rect 556 219 727 235
rect 556 185 693 219
rect 556 169 727 185
rect 761 187 795 264
rect 869 230 903 364
rect 1030 391 1123 401
rect 1030 357 1042 391
rect 1076 365 1123 391
rect 556 119 601 169
rect 761 137 795 153
rect 829 196 903 230
rect 959 323 996 344
rect 959 289 960 323
rect 994 289 996 323
rect 959 287 996 289
rect 993 253 996 287
rect 959 225 996 253
rect 305 100 357 103
rect 305 85 307 100
rect 103 17 169 59
rect 271 66 307 85
rect 341 66 357 100
rect 271 51 357 66
rect 447 93 513 103
rect 447 59 463 93
rect 497 59 513 93
rect 447 17 513 59
rect 556 85 567 119
rect 556 51 601 85
rect 637 106 703 122
rect 637 72 653 106
rect 687 72 703 106
rect 637 17 703 72
rect 829 119 883 196
rect 1030 191 1064 357
rect 1098 331 1123 365
rect 1157 315 1191 435
rect 1225 451 1232 485
rect 1266 451 1272 485
rect 1225 417 1272 451
rect 1225 383 1232 417
rect 1266 383 1272 417
rect 1225 367 1272 383
rect 1306 485 1372 493
rect 1306 451 1322 485
rect 1356 451 1372 485
rect 1306 393 1372 451
rect 1414 472 1472 527
rect 1414 438 1426 472
rect 1460 438 1472 472
rect 1812 485 1846 527
rect 1414 421 1472 438
rect 1585 469 1778 471
rect 1585 435 1601 469
rect 1635 435 1778 469
rect 1585 433 1778 435
rect 1306 359 1322 393
rect 1356 359 1372 393
rect 1157 299 1272 315
rect 1157 297 1238 299
rect 963 157 979 191
rect 1013 157 1064 191
rect 963 147 1064 157
rect 1102 265 1238 297
rect 1102 263 1272 265
rect 829 85 837 119
rect 871 106 883 119
rect 1102 113 1136 263
rect 1238 249 1272 263
rect 1306 275 1372 359
rect 1558 391 1596 393
rect 1558 357 1560 391
rect 1594 357 1596 391
rect 1558 299 1596 357
rect 1306 259 1489 275
rect 1306 225 1455 259
rect 1592 265 1596 299
rect 1558 249 1596 265
rect 1630 365 1694 399
rect 1630 331 1660 365
rect 1630 323 1694 331
rect 1630 289 1644 323
rect 1678 289 1694 323
rect 1174 213 1214 219
rect 1306 213 1489 225
rect 1174 209 1489 213
rect 1174 203 1387 209
rect 1630 207 1694 289
rect 1208 169 1387 203
rect 1174 163 1387 169
rect 1174 153 1336 163
rect 829 72 841 85
rect 875 72 883 106
rect 829 51 883 72
rect 1001 99 1136 113
rect 1306 129 1336 153
rect 1370 129 1387 163
rect 1601 191 1694 207
rect 1635 157 1694 191
rect 1601 141 1694 157
rect 1728 391 1778 433
rect 1728 357 1736 391
rect 1770 357 1778 391
rect 1001 65 1023 99
rect 1057 65 1136 99
rect 1001 51 1136 65
rect 1189 101 1268 112
rect 1189 67 1218 101
rect 1252 67 1268 101
rect 1189 17 1268 67
rect 1306 95 1387 129
rect 1306 61 1336 95
rect 1370 61 1387 95
rect 1306 51 1387 61
rect 1433 107 1488 123
rect 1728 107 1778 357
rect 1812 417 1846 451
rect 1812 349 1846 383
rect 1812 299 1846 315
rect 1880 479 1946 493
rect 1880 445 1896 479
rect 1930 445 1946 479
rect 1880 411 1946 445
rect 1880 377 1896 411
rect 1930 377 1946 411
rect 2060 485 2128 493
rect 2060 451 2076 485
rect 2110 451 2128 485
rect 2060 415 2128 451
rect 1880 343 1946 377
rect 1880 309 1896 343
rect 1930 309 1946 343
rect 1980 391 2026 402
rect 1980 331 1986 391
rect 2020 331 2026 391
rect 1980 315 2026 331
rect 2060 381 2076 415
rect 2110 381 2128 415
rect 1880 282 1946 309
rect 1880 213 1969 282
rect 2060 244 2128 381
rect 2162 479 2211 527
rect 2162 445 2175 479
rect 2209 445 2211 479
rect 2162 411 2211 445
rect 2162 377 2175 411
rect 2209 377 2211 411
rect 2162 343 2211 377
rect 2162 309 2175 343
rect 2209 309 2211 343
rect 2162 293 2211 309
rect 2245 479 2311 484
rect 2245 445 2261 479
rect 2295 445 2311 479
rect 2245 411 2311 445
rect 2245 377 2261 411
rect 2295 377 2311 411
rect 2245 343 2311 377
rect 2245 309 2261 343
rect 2295 309 2311 343
rect 1433 73 1440 107
rect 1474 73 1488 107
rect 1433 17 1488 73
rect 1605 104 1778 107
rect 1605 70 1624 104
rect 1658 70 1778 104
rect 1605 66 1778 70
rect 1819 164 1869 180
rect 1819 130 1835 164
rect 1819 96 1869 130
rect 1819 62 1835 96
rect 1819 17 1869 62
rect 1903 164 1969 213
rect 2003 228 2128 244
rect 2037 194 2128 228
rect 2003 187 2128 194
rect 2003 178 2078 187
rect 1903 130 1919 164
rect 1953 130 1969 164
rect 1903 96 1969 130
rect 1903 62 1919 96
rect 1953 62 1969 96
rect 1903 51 1969 62
rect 2060 153 2078 178
rect 2112 153 2128 187
rect 2060 94 2128 153
rect 2060 60 2078 94
rect 2112 60 2128 94
rect 2060 51 2128 60
rect 2162 164 2211 180
rect 2162 130 2175 164
rect 2209 130 2211 164
rect 2162 96 2211 130
rect 2162 62 2175 96
rect 2209 62 2211 96
rect 2162 17 2211 62
rect 2245 164 2311 309
rect 2245 130 2261 164
rect 2295 130 2311 164
rect 2245 96 2311 130
rect 2245 62 2261 96
rect 2295 62 2311 96
rect 2245 51 2311 62
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 127 357 161 391
rect 203 289 237 323
rect 1042 365 1076 391
rect 1042 357 1064 365
rect 1064 357 1076 365
rect 271 85 305 119
rect 761 153 795 187
rect 960 289 994 323
rect 837 106 871 119
rect 1560 357 1594 391
rect 1644 289 1678 323
rect 837 85 841 106
rect 841 85 871 106
rect 1736 357 1770 391
rect 1986 365 2020 391
rect 1986 357 2020 365
rect 2078 153 2112 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 496 2392 527
rect 115 391 173 397
rect 115 357 127 391
rect 161 388 173 391
rect 1030 391 1088 397
rect 1030 388 1042 391
rect 161 360 1042 388
rect 161 357 173 360
rect 115 351 173 357
rect 1030 357 1042 360
rect 1076 388 1088 391
rect 1548 391 1606 397
rect 1548 388 1560 391
rect 1076 360 1560 388
rect 1076 357 1088 360
rect 1030 351 1088 357
rect 1548 357 1560 360
rect 1594 357 1606 391
rect 1548 351 1606 357
rect 1724 391 1782 397
rect 1724 357 1736 391
rect 1770 388 1782 391
rect 1974 391 2032 397
rect 1974 388 1986 391
rect 1770 360 1986 388
rect 1770 357 1782 360
rect 1724 351 1782 357
rect 1974 357 1986 360
rect 2020 357 2032 391
rect 1974 351 2032 357
rect 191 323 249 329
rect 191 289 203 323
rect 237 320 249 323
rect 948 323 1006 329
rect 948 320 960 323
rect 237 292 960 320
rect 237 289 249 292
rect 191 283 249 289
rect 948 289 960 292
rect 994 320 1006 323
rect 1632 323 1690 329
rect 1632 320 1644 323
rect 994 292 1644 320
rect 994 289 1006 292
rect 948 283 1006 289
rect 1632 289 1644 292
rect 1678 289 1690 323
rect 1632 283 1690 289
rect 749 187 807 193
rect 749 153 761 187
rect 795 184 807 187
rect 2066 187 2124 193
rect 2066 184 2078 187
rect 795 156 2078 184
rect 795 153 807 156
rect 749 147 807 153
rect 2066 153 2078 156
rect 2112 153 2124 187
rect 2066 147 2124 153
rect 259 119 317 125
rect 259 85 271 119
rect 305 116 317 119
rect 825 119 883 125
rect 825 116 837 119
rect 305 85 837 116
rect 871 85 883 119
rect 259 79 883 85
rect 0 17 2392 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< labels >>
rlabel comment s 0 0 0 0 4 edfxbp_1
flabel comment s 973 304 973 304 0 FreeSans 200 0 0 0 clkpos
flabel comment s 1060 374 1060 374 0 FreeSans 200 0 0 0 clkneg
flabel comment s 2005 374 2005 374 0 FreeSans 200 0 0 0 S0
flabel comment s 219 304 219 304 0 FreeSans 200 0 0 0 clkpos
flabel comment s 147 374 147 374 0 FreeSans 200 0 0 0 clkneg
flabel comment s 623 209 623 209 0 FreeSans 200 0 0 0 deneg
flabel comment s 855 104 855 104 0 FreeSans 200 0 0 0 db
flabel comment s 749 446 749 446 0 FreeSans 200 0 0 0 q1
flabel comment s 2096 446 2096 446 0 FreeSans 200 0 0 0 q1
flabel comment s 1660 304 1660 304 0 FreeSans 200 0 0 0 clkpos
flabel comment s 1577 374 1577 374 0 FreeSans 200 0 0 0 clkneg
flabel comment s 1752 374 1752 374 0 FreeSans 200 0 0 0 S0
flabel comment s 1256 269 1256 269 0 FreeSans 200 0 0 0 M0
flabel comment s 1342 269 1342 269 0 FreeSans 200 0 0 0 M1
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1905 221 1939 255 0 FreeSans 400 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 426 153 460 187 0 FreeSans 400 0 0 0 DE
port 3 nsew signal input
flabel locali s 344 221 378 255 0 FreeSans 400 0 0 0 D
port 2 nsew signal input
flabel locali s 2259 221 2293 255 0 FreeSans 400 0 0 0 Q
port 8 nsew signal output
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel pwell s 29 -17 63 17 0 FreeSans 400 0 0 0 VNB
port 5 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2392 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 386760
string GDS_START 367776
<< end >>
