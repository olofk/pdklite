magic
tech sky130A
magscale 1 2
timestamp 1640697850
<< nwell >>
rect 1 37 1415 346
rect 1 14 1490 37
rect 1 -101 483 14
rect 1280 -294 1490 14
<< pwell >>
rect 41 613 1375 749
<< mvnmos >>
rect 120 639 240 723
rect 296 639 416 723
rect 472 639 592 723
rect 648 639 768 723
rect 824 639 944 723
rect 1000 639 1120 723
rect 1176 639 1296 723
<< mvpmos >>
rect 120 80 240 280
rect 296 80 416 280
rect 472 80 592 280
rect 648 80 768 280
rect 824 80 944 280
rect 1000 80 1120 280
rect 1176 80 1296 280
<< mvndiff >>
rect 67 685 120 723
rect 67 651 75 685
rect 109 651 120 685
rect 67 639 120 651
rect 240 685 296 723
rect 240 651 251 685
rect 285 651 296 685
rect 240 639 296 651
rect 416 685 472 723
rect 416 651 427 685
rect 461 651 472 685
rect 416 639 472 651
rect 592 685 648 723
rect 592 651 603 685
rect 637 651 648 685
rect 592 639 648 651
rect 768 685 824 723
rect 768 651 779 685
rect 813 651 824 685
rect 768 639 824 651
rect 944 685 1000 723
rect 944 651 955 685
rect 989 651 1000 685
rect 944 639 1000 651
rect 1120 685 1176 723
rect 1120 651 1131 685
rect 1165 651 1176 685
rect 1120 639 1176 651
rect 1296 685 1349 723
rect 1296 651 1307 685
rect 1341 651 1349 685
rect 1296 639 1349 651
<< mvpdiff >>
rect 67 262 120 280
rect 67 228 75 262
rect 109 228 120 262
rect 67 194 120 228
rect 67 160 75 194
rect 109 160 120 194
rect 67 126 120 160
rect 67 92 75 126
rect 109 92 120 126
rect 67 80 120 92
rect 240 262 296 280
rect 240 228 251 262
rect 285 228 296 262
rect 240 194 296 228
rect 240 160 251 194
rect 285 160 296 194
rect 240 126 296 160
rect 240 92 251 126
rect 285 92 296 126
rect 240 80 296 92
rect 416 262 472 280
rect 416 228 427 262
rect 461 228 472 262
rect 416 194 472 228
rect 416 160 427 194
rect 461 160 472 194
rect 416 126 472 160
rect 416 92 427 126
rect 461 92 472 126
rect 416 80 472 92
rect 592 262 648 280
rect 592 228 603 262
rect 637 228 648 262
rect 592 194 648 228
rect 592 160 603 194
rect 637 160 648 194
rect 592 126 648 160
rect 592 92 603 126
rect 637 92 648 126
rect 592 80 648 92
rect 768 262 824 280
rect 768 228 779 262
rect 813 228 824 262
rect 768 194 824 228
rect 768 160 779 194
rect 813 160 824 194
rect 768 126 824 160
rect 768 92 779 126
rect 813 92 824 126
rect 768 80 824 92
rect 944 262 1000 280
rect 944 228 955 262
rect 989 228 1000 262
rect 944 194 1000 228
rect 944 160 955 194
rect 989 160 1000 194
rect 944 126 1000 160
rect 944 92 955 126
rect 989 92 1000 126
rect 944 80 1000 92
rect 1120 262 1176 280
rect 1120 228 1131 262
rect 1165 228 1176 262
rect 1120 194 1176 228
rect 1120 160 1131 194
rect 1165 160 1176 194
rect 1120 126 1176 160
rect 1120 92 1131 126
rect 1165 92 1176 126
rect 1120 80 1176 92
rect 1296 262 1349 280
rect 1296 228 1307 262
rect 1341 228 1349 262
rect 1296 194 1349 228
rect 1296 160 1307 194
rect 1341 160 1349 194
rect 1296 126 1349 160
rect 1296 92 1307 126
rect 1341 92 1349 126
rect 1296 80 1349 92
<< mvndiffc >>
rect 75 651 109 685
rect 251 651 285 685
rect 427 651 461 685
rect 603 651 637 685
rect 779 651 813 685
rect 955 651 989 685
rect 1131 651 1165 685
rect 1307 651 1341 685
<< mvpdiffc >>
rect 75 228 109 262
rect 75 160 109 194
rect 75 92 109 126
rect 251 228 285 262
rect 251 160 285 194
rect 251 92 285 126
rect 427 228 461 262
rect 427 160 461 194
rect 427 92 461 126
rect 603 228 637 262
rect 603 160 637 194
rect 603 92 637 126
rect 779 228 813 262
rect 779 160 813 194
rect 779 92 813 126
rect 955 228 989 262
rect 955 160 989 194
rect 955 92 989 126
rect 1131 228 1165 262
rect 1131 160 1165 194
rect 1131 92 1165 126
rect 1307 228 1341 262
rect 1307 160 1341 194
rect 1307 92 1341 126
<< mvnsubdiff >>
rect 67 -35 91 -1
rect 125 -35 181 -1
rect 215 -35 270 -1
rect 304 -35 359 -1
rect 393 -35 417 -1
<< mvnsubdiffcont >>
rect 91 -35 125 -1
rect 181 -35 215 -1
rect 270 -35 304 -1
rect 359 -35 393 -1
<< poly >>
rect 120 723 240 755
rect 296 723 416 755
rect 472 723 592 755
rect 648 723 768 755
rect 824 723 944 755
rect 1000 723 1120 755
rect 1176 723 1296 755
rect 120 607 240 639
rect 296 607 416 639
rect 472 607 592 639
rect 648 607 768 639
rect 824 607 944 639
rect 1000 607 1120 639
rect 1176 607 1296 639
rect 120 582 768 607
rect 120 548 136 582
rect 170 548 213 582
rect 247 548 290 582
rect 324 548 366 582
rect 400 548 460 582
rect 494 548 543 582
rect 577 548 625 582
rect 659 548 707 582
rect 741 548 768 582
rect 120 527 768 548
rect 823 582 1296 607
rect 823 548 860 582
rect 894 548 938 582
rect 972 548 1015 582
rect 1049 548 1092 582
rect 1126 548 1169 582
rect 1203 548 1246 582
rect 1280 548 1296 582
rect 120 496 416 527
rect 120 462 136 496
rect 170 462 213 496
rect 247 462 290 496
rect 324 462 366 496
rect 400 462 416 496
rect 120 410 416 462
rect 120 376 136 410
rect 170 376 213 410
rect 247 376 290 410
rect 324 376 366 410
rect 400 376 416 410
rect 823 482 1296 548
rect 823 448 860 482
rect 894 448 938 482
rect 972 448 1015 482
rect 1049 448 1092 482
rect 1126 448 1169 482
rect 1203 448 1246 482
rect 1280 448 1296 482
rect 823 398 1296 448
rect 120 312 416 376
rect 120 280 240 312
rect 296 280 416 312
rect 472 382 1296 398
rect 472 348 494 382
rect 528 348 567 382
rect 601 348 640 382
rect 674 348 713 382
rect 747 348 786 382
rect 820 348 860 382
rect 894 348 938 382
rect 972 348 1015 382
rect 1049 348 1092 382
rect 1126 348 1169 382
rect 1203 348 1246 382
rect 1280 348 1296 382
rect 472 312 1296 348
rect 472 280 592 312
rect 648 280 768 312
rect 824 280 944 312
rect 1000 280 1120 312
rect 1176 280 1296 312
rect 120 48 240 80
rect 296 48 416 80
rect 472 48 592 80
rect 648 48 768 80
rect 824 48 944 80
rect 1000 48 1120 80
rect 1176 48 1296 80
<< polycont >>
rect 136 548 170 582
rect 213 548 247 582
rect 290 548 324 582
rect 366 548 400 582
rect 460 548 494 582
rect 543 548 577 582
rect 625 548 659 582
rect 707 548 741 582
rect 860 548 894 582
rect 938 548 972 582
rect 1015 548 1049 582
rect 1092 548 1126 582
rect 1169 548 1203 582
rect 1246 548 1280 582
rect 136 462 170 496
rect 213 462 247 496
rect 290 462 324 496
rect 366 462 400 496
rect 136 376 170 410
rect 213 376 247 410
rect 290 376 324 410
rect 366 376 400 410
rect 860 448 894 482
rect 938 448 972 482
rect 1015 448 1049 482
rect 1092 448 1126 482
rect 1169 448 1203 482
rect 1246 448 1280 482
rect 494 348 528 382
rect 567 348 601 382
rect 640 348 674 382
rect 713 348 747 382
rect 786 348 820 382
rect 860 348 894 382
rect 938 348 972 382
rect 1015 348 1049 382
rect 1092 348 1126 382
rect 1169 348 1203 382
rect 1246 348 1280 382
<< locali >>
rect 64 772 120 797
rect 416 772 472 797
rect 768 772 824 797
rect 1120 772 1173 797
rect 64 738 69 772
rect 103 738 143 772
rect 177 738 217 772
rect 251 738 290 772
rect 324 738 363 772
rect 397 738 436 772
rect 470 738 509 772
rect 543 738 582 772
rect 616 738 655 772
rect 689 738 728 772
rect 762 738 801 772
rect 835 738 874 772
rect 908 738 947 772
rect 981 738 1020 772
rect 1054 738 1093 772
rect 1127 738 1166 772
rect 1200 738 1239 772
rect 1273 738 1312 772
rect 64 685 120 738
rect 64 651 75 685
rect 109 651 120 685
rect 251 685 285 701
rect 416 685 472 738
rect 64 635 120 651
rect 245 651 251 669
rect 245 635 283 651
rect 416 651 427 685
rect 461 651 472 685
rect 603 685 637 701
rect 768 685 824 738
rect 416 619 472 651
rect 637 651 663 669
rect 625 635 663 651
rect 768 651 779 685
rect 813 651 824 685
rect 955 685 989 701
rect 768 635 824 651
rect 953 651 955 669
rect 1120 685 1173 738
rect 989 651 991 669
rect 953 635 991 651
rect 1120 651 1131 685
rect 1165 651 1173 685
rect 1307 685 1341 701
rect 1120 619 1173 651
rect 1264 635 1302 669
rect 1336 635 1341 651
rect 120 582 416 583
rect 120 548 136 582
rect 170 548 213 582
rect 247 548 290 582
rect 324 548 366 582
rect 400 548 460 582
rect 494 548 543 582
rect 577 548 625 582
rect 659 548 707 582
rect 741 548 757 582
rect 844 548 860 582
rect 894 548 938 582
rect 972 548 1015 582
rect 1049 548 1092 582
rect 1126 548 1169 582
rect 1203 548 1246 582
rect 1280 548 1296 582
rect 120 496 416 548
rect 120 481 136 496
rect 120 447 132 481
rect 170 462 213 496
rect 247 481 290 496
rect 324 481 366 496
rect 261 462 290 481
rect 356 462 366 481
rect 400 462 416 496
rect 166 447 227 462
rect 261 447 322 462
rect 356 447 416 462
rect 120 410 416 447
rect 120 409 136 410
rect 120 375 132 409
rect 170 376 213 410
rect 247 409 290 410
rect 324 409 366 410
rect 261 376 290 409
rect 356 376 366 409
rect 400 376 416 410
rect 844 482 1296 548
rect 844 448 860 482
rect 894 448 938 482
rect 972 448 1015 482
rect 1049 448 1092 482
rect 1126 448 1169 482
rect 1203 448 1246 482
rect 1280 448 1296 482
rect 524 382 575 383
rect 609 382 660 383
rect 694 382 745 383
rect 844 382 1296 448
rect 166 375 227 376
rect 261 375 322 376
rect 356 375 416 376
rect 478 349 490 382
rect 478 348 494 349
rect 528 348 567 382
rect 609 349 640 382
rect 694 349 713 382
rect 779 349 786 382
rect 601 348 640 349
rect 674 348 713 349
rect 747 348 786 349
rect 820 348 860 382
rect 894 348 938 382
rect 972 348 1015 382
rect 1049 348 1092 382
rect 1126 348 1169 382
rect 1203 348 1246 382
rect 1280 348 1296 382
rect 75 262 109 278
rect 75 194 109 228
rect 75 138 109 160
rect 75 66 109 92
rect 251 262 285 272
rect 251 194 285 200
rect 251 126 285 160
rect 251 76 285 92
rect 427 262 461 278
rect 603 262 637 278
rect 779 262 813 278
rect 427 194 461 228
rect 618 194 656 228
rect 779 194 813 228
rect 427 138 461 160
rect 427 66 461 92
rect 603 126 637 160
rect 603 76 637 92
rect 779 138 813 160
rect 779 66 813 92
rect 955 262 989 272
rect 955 194 989 200
rect 955 126 989 160
rect 955 76 989 92
rect 1131 262 1165 278
rect 1131 194 1165 228
rect 1131 138 1165 160
rect 1131 66 1165 92
rect 1307 272 1309 278
rect 1307 262 1343 272
rect 1341 234 1343 262
rect 1307 200 1309 228
rect 1307 194 1341 200
rect 1307 126 1341 160
rect 1307 76 1341 92
rect 75 -1 109 32
rect 67 -6 91 -1
rect 125 -6 181 -1
rect 215 -6 270 -1
rect 304 -6 359 -1
rect 393 -6 417 -1
rect 67 -35 79 -6
rect 125 -35 152 -6
rect 215 -35 225 -6
rect 113 -40 152 -35
rect 186 -40 225 -35
rect 259 -35 270 -6
rect 332 -35 359 -6
rect 405 -35 417 -6
rect 259 -40 298 -35
rect 332 -40 371 -35
<< viali >>
rect 69 738 103 772
rect 143 738 177 772
rect 217 738 251 772
rect 290 738 324 772
rect 363 738 397 772
rect 436 738 470 772
rect 509 738 543 772
rect 582 738 616 772
rect 655 738 689 772
rect 728 738 762 772
rect 801 738 835 772
rect 874 738 908 772
rect 947 738 981 772
rect 1020 738 1054 772
rect 1093 738 1127 772
rect 1166 738 1200 772
rect 1239 738 1273 772
rect 1312 738 1346 772
rect 211 635 245 669
rect 283 651 285 669
rect 285 651 317 669
rect 283 635 317 651
rect 591 651 603 669
rect 603 651 625 669
rect 591 635 625 651
rect 663 635 697 669
rect 919 635 953 669
rect 991 635 1025 669
rect 1230 635 1264 669
rect 1302 651 1307 669
rect 1307 651 1336 669
rect 1302 635 1336 651
rect 132 462 136 481
rect 136 462 166 481
rect 227 462 247 481
rect 247 462 261 481
rect 322 462 324 481
rect 324 462 356 481
rect 132 447 166 462
rect 227 447 261 462
rect 322 447 356 462
rect 132 376 136 409
rect 136 376 166 409
rect 227 376 247 409
rect 247 376 261 409
rect 322 376 324 409
rect 324 376 356 409
rect 490 382 524 383
rect 575 382 609 383
rect 660 382 694 383
rect 745 382 779 383
rect 132 375 166 376
rect 227 375 261 376
rect 322 375 356 376
rect 490 349 494 382
rect 494 349 524 382
rect 575 349 601 382
rect 601 349 609 382
rect 660 349 674 382
rect 674 349 694 382
rect 745 349 747 382
rect 747 349 779 382
rect 75 126 109 138
rect 75 104 109 126
rect 251 272 285 306
rect 251 228 285 234
rect 251 200 285 228
rect 584 194 618 228
rect 656 194 690 228
rect 427 126 461 138
rect 427 104 461 126
rect 75 32 109 66
rect 779 126 813 138
rect 779 104 813 126
rect 427 32 461 66
rect 955 272 989 306
rect 955 228 989 234
rect 955 200 989 228
rect 1131 126 1165 138
rect 1131 104 1165 126
rect 779 32 813 66
rect 1309 272 1343 306
rect 1309 228 1341 234
rect 1341 228 1343 234
rect 1309 200 1343 228
rect 1131 32 1165 66
rect 79 -35 91 -6
rect 91 -35 113 -6
rect 152 -35 181 -6
rect 181 -35 186 -6
rect 79 -40 113 -35
rect 152 -40 186 -35
rect 225 -40 259 -6
rect 298 -35 304 -6
rect 304 -35 332 -6
rect 371 -35 393 -6
rect 393 -35 405 -6
rect 298 -40 332 -35
rect 371 -40 405 -35
<< metal1 >>
rect 56 772 1358 792
rect 56 738 69 772
rect 103 738 143 772
rect 177 738 217 772
rect 251 738 290 772
rect 324 738 363 772
rect 397 738 436 772
rect 470 738 509 772
rect 543 738 582 772
rect 616 738 655 772
rect 689 738 728 772
rect 762 738 801 772
rect 835 738 874 772
rect 908 738 947 772
rect 981 738 1020 772
rect 1054 738 1093 772
rect 1127 738 1166 772
rect 1200 738 1239 772
rect 1273 738 1312 772
rect 1346 738 1358 772
rect 56 711 1358 738
rect 191 669 709 675
rect 191 635 211 669
rect 245 635 283 669
rect 317 635 591 669
rect 625 635 663 669
rect 697 635 709 669
rect 191 629 709 635
rect 873 669 1350 675
rect 873 635 919 669
rect 953 635 991 669
rect 1025 635 1230 669
rect 1264 635 1302 669
rect 1336 635 1350 669
rect 191 625 530 629
rect 120 481 368 487
rect 120 447 132 481
rect 166 447 227 481
rect 261 447 322 481
rect 356 447 368 481
rect 120 409 368 447
rect 120 375 132 409
rect 166 375 227 409
rect 261 375 322 409
rect 356 375 368 409
rect 120 369 368 375
rect 398 389 530 625
rect 398 383 791 389
rect 398 349 490 383
rect 524 349 575 383
rect 609 349 660 383
rect 694 349 745 383
rect 779 349 791 383
rect 398 343 791 349
rect 398 318 530 343
rect 67 306 530 318
rect 67 272 251 306
rect 285 272 530 306
rect 873 306 1350 635
rect 873 299 955 306
rect 67 234 530 272
rect 67 200 251 234
rect 285 200 530 234
rect 67 188 530 200
rect 572 272 955 299
rect 989 272 1309 306
rect 1343 272 1350 306
rect 572 234 1350 272
rect 572 228 955 234
rect 572 194 584 228
rect 618 194 656 228
rect 690 200 955 228
rect 989 200 1309 234
rect 1343 200 1350 234
rect 690 194 1350 200
rect 572 188 1350 194
rect 67 138 1349 151
rect 67 104 75 138
rect 109 104 427 138
rect 461 104 779 138
rect 813 104 1131 138
rect 1165 104 1349 138
rect 67 66 1349 104
rect 67 32 75 66
rect 109 32 427 66
rect 461 32 779 66
rect 813 32 1131 66
rect 1165 32 1349 66
rect 67 -6 1349 32
rect 67 -40 79 -6
rect 113 -40 152 -6
rect 186 -40 225 -6
rect 259 -40 298 -6
rect 332 -40 371 -6
rect 405 -40 1349 -6
rect 67 -41 1349 -40
rect 67 -46 417 -41
use sky130_fd_pr__nfet_01v8__example_55959141808487  sky130_fd_pr__nfet_01v8__example_55959141808487_0
timestamp 1640697850
transform 1 0 120 0 1 639
box -28 0 1204 29
use sky130_fd_pr__pfet_01v8__example_55959141808486  sky130_fd_pr__pfet_01v8__example_55959141808486_0
timestamp 1640697850
transform 1 0 120 0 1 80
box -28 0 1204 97
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 48538054
string GDS_START 48527122
<< end >>
