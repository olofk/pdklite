magic
tech sky130A
magscale 1 2
timestamp 1619729579
<< nwell >>
rect -66 1201 102 1251
rect -66 419 1204 1201
rect -66 377 102 419
rect 1778 409 2142 1219
<< pwell >>
rect 0 1611 2784 1645
rect 0 -17 2784 17
<< locali >>
rect 191 539 235 615
rect 151 481 235 539
rect 151 321 195 481
rect 151 263 235 321
rect 191 179 235 263
rect 946 366 1080 432
rect 1841 337 1979 403
<< obsli1 >>
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2143 1645
rect 2177 1611 2239 1645
rect 2273 1611 2335 1645
rect 2369 1611 2431 1645
rect 2465 1611 2527 1645
rect 2561 1611 2623 1645
rect 2657 1611 2719 1645
rect 2753 1611 2784 1645
rect 191 1525 980 1569
rect 191 1289 235 1525
rect 347 1255 391 1491
rect 503 1289 547 1525
rect 179 1211 391 1255
rect 72 831 106 1056
rect 179 959 223 1211
rect 659 1177 703 1491
rect 815 1289 859 1525
rect 936 1303 980 1525
rect 1941 1544 2059 1550
rect 1941 1510 1947 1544
rect 1981 1510 2019 1544
rect 2053 1510 2059 1544
rect 1941 1504 2059 1510
rect 1550 1415 1907 1481
rect 936 1259 1689 1303
rect 273 1133 1135 1177
rect 273 1111 407 1133
rect 179 915 556 959
rect 422 859 556 915
rect 635 926 679 1081
rect 1091 989 1135 1133
rect 635 882 729 926
rect 0 797 31 831
rect 65 797 103 831
rect 352 689 470 747
rect 352 481 386 689
rect 512 617 556 859
rect 685 747 729 882
rect 612 689 729 747
rect 452 572 556 617
rect 352 125 398 313
rect 452 129 496 572
rect 685 481 729 689
rect 841 432 885 751
rect 530 388 885 432
rect 530 366 664 388
rect 672 125 718 331
rect 841 129 885 388
rect 1293 261 1337 1259
rect 1468 125 1514 1211
rect 1645 261 1689 1259
rect 1841 955 1907 1415
rect 1941 1325 2007 1504
rect 1941 1225 2107 1291
rect 1941 847 2007 1161
rect 1820 781 2007 847
rect 1913 673 1979 781
rect 2041 673 2107 1225
rect 1861 650 1979 673
rect 1861 616 1867 650
rect 1901 616 1939 650
rect 1973 616 1979 650
rect 1861 604 1979 616
rect 1913 467 1979 604
rect 2013 607 2107 673
rect 1913 125 1979 303
rect 2013 147 2079 607
rect 280 79 398 125
rect 635 79 753 125
rect 1431 79 1549 125
rect 1861 79 1979 125
rect 0 -17 2784 17
<< obsli1c >>
rect 31 1611 65 1645
rect 127 1611 161 1645
rect 223 1611 257 1645
rect 319 1611 353 1645
rect 415 1611 449 1645
rect 511 1611 545 1645
rect 607 1611 641 1645
rect 703 1611 737 1645
rect 799 1611 833 1645
rect 895 1611 929 1645
rect 991 1611 1025 1645
rect 1087 1611 1121 1645
rect 1183 1611 1217 1645
rect 1279 1611 1313 1645
rect 1375 1611 1409 1645
rect 1471 1611 1505 1645
rect 1567 1611 1601 1645
rect 1663 1611 1697 1645
rect 1759 1611 1793 1645
rect 1855 1611 1889 1645
rect 1951 1611 1985 1645
rect 2047 1611 2081 1645
rect 2143 1611 2177 1645
rect 2239 1611 2273 1645
rect 2335 1611 2369 1645
rect 2431 1611 2465 1645
rect 2527 1611 2561 1645
rect 2623 1611 2657 1645
rect 2719 1611 2753 1645
rect 1947 1510 1981 1544
rect 2019 1510 2053 1544
rect 31 797 65 831
rect 103 797 137 831
rect 1867 616 1901 650
rect 1939 616 1973 650
<< metal1 >>
rect 0 1645 2784 1651
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2143 1645
rect 2177 1611 2239 1645
rect 2273 1611 2335 1645
rect 2369 1611 2431 1645
rect 2465 1611 2527 1645
rect 2561 1611 2623 1645
rect 2657 1611 2719 1645
rect 2753 1611 2784 1645
rect 0 1605 2784 1611
rect 0 1544 2784 1577
rect 0 1510 1947 1544
rect 1981 1510 2019 1544
rect 2053 1510 2784 1544
rect 0 1503 2784 1510
rect 0 865 2784 939
rect 0 831 2784 837
rect 0 797 31 831
rect 65 797 103 831
rect 137 797 2784 831
rect 0 791 2784 797
rect 14 650 2770 661
rect 14 616 1867 650
rect 1901 616 1939 650
rect 1973 616 2770 650
rect 14 604 2770 616
<< obsm1 >>
rect 0 689 2784 763
rect 0 51 2784 125
rect 0 -23 2784 23
<< labels >>
rlabel locali s 1841 337 1979 403 6 A
port 1 nsew signal input
rlabel locali s 946 366 1080 432 6 SLEEP_B
port 2 nsew signal input
rlabel locali s 191 539 235 615 6 X
port 8 nsew signal output
rlabel locali s 191 179 235 263 6 X
port 8 nsew signal output
rlabel locali s 151 481 235 539 6 X
port 8 nsew signal output
rlabel locali s 151 321 195 481 6 X
port 8 nsew signal output
rlabel locali s 151 263 235 321 6 X
port 8 nsew signal output
rlabel nwell s 1778 409 2142 1219 6 LVPWR
port 3 nsew power bidirectional
rlabel metal1 s 14 604 2770 661 6 LVPWR
port 3 nsew power bidirectional
rlabel metal1 s 0 1503 2784 1577 6 VGND
port 4 nsew ground bidirectional
rlabel pwell s 0 1611 2784 1645 6 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 1605 2784 1651 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -66 1201 102 1251 6 VPB
port 6 nsew power bidirectional
rlabel nwell s -66 419 1204 1201 6 VPB
port 6 nsew power bidirectional
rlabel nwell s -66 377 102 419 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 791 2784 837 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 865 2784 939 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithvdbl
string LEFclass CORE
string FIXED_BBOX 0 0 2784 1628
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_END 1067012
string GDS_START 1037752
<< end >>
