magic
tech sky130A
magscale 1 2
timestamp 1640697675
<< pwell >>
rect 0 1187 1340 1340
rect 0 153 153 1187
rect 1187 153 1340 1187
rect 0 0 1340 153
<< nbase >>
rect 153 153 1187 1187
<< pnp3p40 >>
rect 153 153 1187 1187
<< pdiff >>
rect 330 958 1010 1010
rect 330 924 384 958
rect 418 924 474 958
rect 508 924 564 958
rect 598 924 654 958
rect 688 924 744 958
rect 778 924 834 958
rect 868 924 924 958
rect 958 924 1010 958
rect 330 868 1010 924
rect 330 834 384 868
rect 418 834 474 868
rect 508 834 564 868
rect 598 834 654 868
rect 688 834 744 868
rect 778 834 834 868
rect 868 834 924 868
rect 958 834 1010 868
rect 330 778 1010 834
rect 330 744 384 778
rect 418 744 474 778
rect 508 744 564 778
rect 598 744 654 778
rect 688 744 744 778
rect 778 744 834 778
rect 868 744 924 778
rect 958 744 1010 778
rect 330 688 1010 744
rect 330 654 384 688
rect 418 654 474 688
rect 508 654 564 688
rect 598 654 654 688
rect 688 654 744 688
rect 778 654 834 688
rect 868 654 924 688
rect 958 654 1010 688
rect 330 598 1010 654
rect 330 564 384 598
rect 418 564 474 598
rect 508 564 564 598
rect 598 564 654 598
rect 688 564 744 598
rect 778 564 834 598
rect 868 564 924 598
rect 958 564 1010 598
rect 330 508 1010 564
rect 330 474 384 508
rect 418 474 474 508
rect 508 474 564 508
rect 598 474 654 508
rect 688 474 744 508
rect 778 474 834 508
rect 868 474 924 508
rect 958 474 1010 508
rect 330 418 1010 474
rect 330 384 384 418
rect 418 384 474 418
rect 508 384 564 418
rect 598 384 654 418
rect 688 384 744 418
rect 778 384 834 418
rect 868 384 924 418
rect 958 384 1010 418
rect 330 330 1010 384
<< pdiffc >>
rect 384 924 418 958
rect 474 924 508 958
rect 564 924 598 958
rect 654 924 688 958
rect 744 924 778 958
rect 834 924 868 958
rect 924 924 958 958
rect 384 834 418 868
rect 474 834 508 868
rect 564 834 598 868
rect 654 834 688 868
rect 744 834 778 868
rect 834 834 868 868
rect 924 834 958 868
rect 384 744 418 778
rect 474 744 508 778
rect 564 744 598 778
rect 654 744 688 778
rect 744 744 778 778
rect 834 744 868 778
rect 924 744 958 778
rect 384 654 418 688
rect 474 654 508 688
rect 564 654 598 688
rect 654 654 688 688
rect 744 654 778 688
rect 834 654 868 688
rect 924 654 958 688
rect 384 564 418 598
rect 474 564 508 598
rect 564 564 598 598
rect 654 564 688 598
rect 744 564 778 598
rect 834 564 868 598
rect 924 564 958 598
rect 384 474 418 508
rect 474 474 508 508
rect 564 474 598 508
rect 654 474 688 508
rect 744 474 778 508
rect 834 474 868 508
rect 924 474 958 508
rect 384 384 418 418
rect 474 384 508 418
rect 564 384 598 418
rect 654 384 688 418
rect 744 384 778 418
rect 834 384 868 418
rect 924 384 958 418
<< psubdiff >>
rect 26 1279 1314 1314
rect 26 1256 156 1279
rect 26 1222 60 1256
rect 94 1245 156 1256
rect 190 1245 246 1279
rect 280 1245 336 1279
rect 370 1245 426 1279
rect 460 1245 516 1279
rect 550 1245 606 1279
rect 640 1245 696 1279
rect 730 1245 786 1279
rect 820 1245 876 1279
rect 910 1245 966 1279
rect 1000 1245 1056 1279
rect 1090 1245 1146 1279
rect 1180 1256 1314 1279
rect 1180 1245 1247 1256
rect 94 1222 1247 1245
rect 1281 1222 1314 1256
rect 26 1213 1314 1222
rect 26 1166 127 1213
rect 26 1132 60 1166
rect 94 1132 127 1166
rect 1213 1166 1314 1213
rect 26 1076 127 1132
rect 26 1042 60 1076
rect 94 1042 127 1076
rect 26 986 127 1042
rect 26 952 60 986
rect 94 952 127 986
rect 26 896 127 952
rect 26 862 60 896
rect 94 862 127 896
rect 26 806 127 862
rect 26 772 60 806
rect 94 772 127 806
rect 26 716 127 772
rect 26 682 60 716
rect 94 682 127 716
rect 26 626 127 682
rect 26 592 60 626
rect 94 592 127 626
rect 26 536 127 592
rect 26 502 60 536
rect 94 502 127 536
rect 26 446 127 502
rect 26 412 60 446
rect 94 412 127 446
rect 26 356 127 412
rect 26 322 60 356
rect 94 322 127 356
rect 26 266 127 322
rect 26 232 60 266
rect 94 232 127 266
rect 26 176 127 232
rect 1213 1132 1247 1166
rect 1281 1132 1314 1166
rect 1213 1076 1314 1132
rect 1213 1042 1247 1076
rect 1281 1042 1314 1076
rect 1213 986 1314 1042
rect 1213 952 1247 986
rect 1281 952 1314 986
rect 1213 896 1314 952
rect 1213 862 1247 896
rect 1281 862 1314 896
rect 1213 806 1314 862
rect 1213 772 1247 806
rect 1281 772 1314 806
rect 1213 716 1314 772
rect 1213 682 1247 716
rect 1281 682 1314 716
rect 1213 626 1314 682
rect 1213 592 1247 626
rect 1281 592 1314 626
rect 1213 536 1314 592
rect 1213 502 1247 536
rect 1281 502 1314 536
rect 1213 446 1314 502
rect 1213 412 1247 446
rect 1281 412 1314 446
rect 1213 356 1314 412
rect 1213 322 1247 356
rect 1281 322 1314 356
rect 1213 266 1314 322
rect 1213 232 1247 266
rect 1281 232 1314 266
rect 26 142 60 176
rect 94 142 127 176
rect 26 127 127 142
rect 1213 176 1314 232
rect 1213 142 1247 176
rect 1281 142 1314 176
rect 1213 127 1314 142
rect 26 92 1314 127
rect 26 58 156 92
rect 190 58 246 92
rect 280 58 336 92
rect 370 58 426 92
rect 460 58 516 92
rect 550 58 606 92
rect 640 58 696 92
rect 730 58 786 92
rect 820 58 876 92
rect 910 58 966 92
rect 1000 58 1056 92
rect 1090 58 1146 92
rect 1180 58 1314 92
rect 26 26 1314 58
<< nsubdiff >>
rect 189 1132 1151 1151
rect 189 1098 320 1132
rect 354 1098 410 1132
rect 444 1098 500 1132
rect 534 1098 590 1132
rect 624 1098 680 1132
rect 714 1098 770 1132
rect 804 1098 860 1132
rect 894 1098 950 1132
rect 984 1098 1040 1132
rect 1074 1098 1151 1132
rect 189 1079 1151 1098
rect 189 1075 261 1079
rect 189 1041 208 1075
rect 242 1041 261 1075
rect 189 985 261 1041
rect 1079 1056 1151 1079
rect 1079 1022 1098 1056
rect 1132 1022 1151 1056
rect 189 951 208 985
rect 242 951 261 985
rect 189 895 261 951
rect 189 861 208 895
rect 242 861 261 895
rect 189 805 261 861
rect 189 771 208 805
rect 242 771 261 805
rect 189 715 261 771
rect 189 681 208 715
rect 242 681 261 715
rect 189 625 261 681
rect 189 591 208 625
rect 242 591 261 625
rect 189 535 261 591
rect 189 501 208 535
rect 242 501 261 535
rect 189 445 261 501
rect 189 411 208 445
rect 242 411 261 445
rect 189 355 261 411
rect 189 321 208 355
rect 242 321 261 355
rect 1079 966 1151 1022
rect 1079 932 1098 966
rect 1132 932 1151 966
rect 1079 876 1151 932
rect 1079 842 1098 876
rect 1132 842 1151 876
rect 1079 786 1151 842
rect 1079 752 1098 786
rect 1132 752 1151 786
rect 1079 696 1151 752
rect 1079 662 1098 696
rect 1132 662 1151 696
rect 1079 606 1151 662
rect 1079 572 1098 606
rect 1132 572 1151 606
rect 1079 516 1151 572
rect 1079 482 1098 516
rect 1132 482 1151 516
rect 1079 426 1151 482
rect 1079 392 1098 426
rect 1132 392 1151 426
rect 1079 336 1151 392
rect 189 261 261 321
rect 1079 302 1098 336
rect 1132 302 1151 336
rect 1079 261 1151 302
rect 189 242 1151 261
rect 189 208 286 242
rect 320 208 376 242
rect 410 208 466 242
rect 500 208 556 242
rect 590 208 646 242
rect 680 208 736 242
rect 770 208 826 242
rect 860 208 916 242
rect 950 208 1006 242
rect 1040 208 1151 242
rect 189 189 1151 208
<< psubdiffcont >>
rect 60 1222 94 1256
rect 156 1245 190 1279
rect 246 1245 280 1279
rect 336 1245 370 1279
rect 426 1245 460 1279
rect 516 1245 550 1279
rect 606 1245 640 1279
rect 696 1245 730 1279
rect 786 1245 820 1279
rect 876 1245 910 1279
rect 966 1245 1000 1279
rect 1056 1245 1090 1279
rect 1146 1245 1180 1279
rect 1247 1222 1281 1256
rect 60 1132 94 1166
rect 60 1042 94 1076
rect 60 952 94 986
rect 60 862 94 896
rect 60 772 94 806
rect 60 682 94 716
rect 60 592 94 626
rect 60 502 94 536
rect 60 412 94 446
rect 60 322 94 356
rect 60 232 94 266
rect 1247 1132 1281 1166
rect 1247 1042 1281 1076
rect 1247 952 1281 986
rect 1247 862 1281 896
rect 1247 772 1281 806
rect 1247 682 1281 716
rect 1247 592 1281 626
rect 1247 502 1281 536
rect 1247 412 1281 446
rect 1247 322 1281 356
rect 1247 232 1281 266
rect 60 142 94 176
rect 1247 142 1281 176
rect 156 58 190 92
rect 246 58 280 92
rect 336 58 370 92
rect 426 58 460 92
rect 516 58 550 92
rect 606 58 640 92
rect 696 58 730 92
rect 786 58 820 92
rect 876 58 910 92
rect 966 58 1000 92
rect 1056 58 1090 92
rect 1146 58 1180 92
<< nsubdiffcont >>
rect 320 1098 354 1132
rect 410 1098 444 1132
rect 500 1098 534 1132
rect 590 1098 624 1132
rect 680 1098 714 1132
rect 770 1098 804 1132
rect 860 1098 894 1132
rect 950 1098 984 1132
rect 1040 1098 1074 1132
rect 208 1041 242 1075
rect 1098 1022 1132 1056
rect 208 951 242 985
rect 208 861 242 895
rect 208 771 242 805
rect 208 681 242 715
rect 208 591 242 625
rect 208 501 242 535
rect 208 411 242 445
rect 208 321 242 355
rect 1098 932 1132 966
rect 1098 842 1132 876
rect 1098 752 1132 786
rect 1098 662 1132 696
rect 1098 572 1132 606
rect 1098 482 1132 516
rect 1098 392 1132 426
rect 1098 302 1132 336
rect 286 208 320 242
rect 376 208 410 242
rect 466 208 500 242
rect 556 208 590 242
rect 646 208 680 242
rect 736 208 770 242
rect 826 208 860 242
rect 916 208 950 242
rect 1006 208 1040 242
<< locali >>
rect 26 1279 1314 1314
rect 26 1256 156 1279
rect 26 1222 60 1256
rect 94 1245 156 1256
rect 190 1245 246 1279
rect 280 1245 336 1279
rect 370 1245 426 1279
rect 460 1245 516 1279
rect 550 1245 606 1279
rect 640 1245 696 1279
rect 730 1245 786 1279
rect 820 1245 876 1279
rect 910 1245 966 1279
rect 1000 1245 1056 1279
rect 1090 1245 1146 1279
rect 1180 1256 1314 1279
rect 1180 1245 1247 1256
rect 94 1222 1247 1245
rect 1281 1222 1314 1256
rect 26 1215 1314 1222
rect 26 1166 125 1215
rect 26 1132 60 1166
rect 94 1132 125 1166
rect 1215 1166 1314 1215
rect 26 1076 125 1132
rect 26 1042 60 1076
rect 94 1042 125 1076
rect 26 986 125 1042
rect 26 952 60 986
rect 94 952 125 986
rect 26 896 125 952
rect 26 862 60 896
rect 94 862 125 896
rect 26 806 125 862
rect 26 772 60 806
rect 94 772 125 806
rect 26 716 125 772
rect 26 682 60 716
rect 94 682 125 716
rect 26 626 125 682
rect 26 592 60 626
rect 94 592 125 626
rect 26 536 125 592
rect 26 502 60 536
rect 94 502 125 536
rect 26 446 125 502
rect 26 412 60 446
rect 94 412 125 446
rect 26 356 125 412
rect 26 322 60 356
rect 94 322 125 356
rect 26 266 125 322
rect 26 232 60 266
rect 94 232 125 266
rect 26 176 125 232
rect 189 1132 1151 1151
rect 189 1098 320 1132
rect 354 1098 410 1132
rect 444 1098 500 1132
rect 534 1098 590 1132
rect 624 1098 680 1132
rect 714 1098 770 1132
rect 804 1098 860 1132
rect 894 1098 950 1132
rect 984 1098 1040 1132
rect 1074 1098 1151 1132
rect 189 1079 1151 1098
rect 189 1075 261 1079
rect 189 1041 208 1075
rect 242 1041 261 1075
rect 189 985 261 1041
rect 1079 1056 1151 1079
rect 1079 1022 1098 1056
rect 1132 1022 1151 1056
rect 189 951 208 985
rect 242 951 261 985
rect 189 895 261 951
rect 189 861 208 895
rect 242 861 261 895
rect 189 805 261 861
rect 189 771 208 805
rect 242 771 261 805
rect 189 715 261 771
rect 189 681 208 715
rect 242 681 261 715
rect 189 625 261 681
rect 189 591 208 625
rect 242 591 261 625
rect 189 535 261 591
rect 189 501 208 535
rect 242 501 261 535
rect 189 445 261 501
rect 189 411 208 445
rect 242 411 261 445
rect 189 355 261 411
rect 189 321 208 355
rect 242 321 261 355
rect 323 958 1017 1017
rect 323 924 384 958
rect 418 930 474 958
rect 508 930 564 958
rect 598 930 654 958
rect 430 924 474 930
rect 530 924 564 930
rect 630 924 654 930
rect 688 930 744 958
rect 688 924 696 930
rect 323 896 396 924
rect 430 896 496 924
rect 530 896 596 924
rect 630 896 696 924
rect 730 924 744 930
rect 778 930 834 958
rect 778 924 796 930
rect 730 896 796 924
rect 830 924 834 930
rect 868 930 924 958
rect 868 924 896 930
rect 958 924 1017 958
rect 830 896 896 924
rect 930 896 1017 924
rect 323 868 1017 896
rect 323 834 384 868
rect 418 834 474 868
rect 508 834 564 868
rect 598 834 654 868
rect 688 834 744 868
rect 778 834 834 868
rect 868 834 924 868
rect 958 834 1017 868
rect 323 830 1017 834
rect 323 796 396 830
rect 430 796 496 830
rect 530 796 596 830
rect 630 796 696 830
rect 730 796 796 830
rect 830 796 896 830
rect 930 796 1017 830
rect 323 778 1017 796
rect 323 744 384 778
rect 418 744 474 778
rect 508 744 564 778
rect 598 744 654 778
rect 688 744 744 778
rect 778 744 834 778
rect 868 744 924 778
rect 958 744 1017 778
rect 323 730 1017 744
rect 323 696 396 730
rect 430 696 496 730
rect 530 696 596 730
rect 630 696 696 730
rect 730 696 796 730
rect 830 696 896 730
rect 930 696 1017 730
rect 323 688 1017 696
rect 323 654 384 688
rect 418 654 474 688
rect 508 654 564 688
rect 598 654 654 688
rect 688 654 744 688
rect 778 654 834 688
rect 868 654 924 688
rect 958 654 1017 688
rect 323 630 1017 654
rect 323 598 396 630
rect 430 598 496 630
rect 530 598 596 630
rect 630 598 696 630
rect 323 564 384 598
rect 430 596 474 598
rect 530 596 564 598
rect 630 596 654 598
rect 418 564 474 596
rect 508 564 564 596
rect 598 564 654 596
rect 688 596 696 598
rect 730 598 796 630
rect 730 596 744 598
rect 688 564 744 596
rect 778 596 796 598
rect 830 598 896 630
rect 930 598 1017 630
rect 830 596 834 598
rect 778 564 834 596
rect 868 596 896 598
rect 868 564 924 596
rect 958 564 1017 598
rect 323 530 1017 564
rect 323 508 396 530
rect 430 508 496 530
rect 530 508 596 530
rect 630 508 696 530
rect 323 474 384 508
rect 430 496 474 508
rect 530 496 564 508
rect 630 496 654 508
rect 418 474 474 496
rect 508 474 564 496
rect 598 474 654 496
rect 688 496 696 508
rect 730 508 796 530
rect 730 496 744 508
rect 688 474 744 496
rect 778 496 796 508
rect 830 508 896 530
rect 930 508 1017 530
rect 830 496 834 508
rect 778 474 834 496
rect 868 496 896 508
rect 868 474 924 496
rect 958 474 1017 508
rect 323 430 1017 474
rect 323 418 396 430
rect 430 418 496 430
rect 530 418 596 430
rect 630 418 696 430
rect 323 384 384 418
rect 430 396 474 418
rect 530 396 564 418
rect 630 396 654 418
rect 418 384 474 396
rect 508 384 564 396
rect 598 384 654 396
rect 688 396 696 418
rect 730 418 796 430
rect 730 396 744 418
rect 688 384 744 396
rect 778 396 796 418
rect 830 418 896 430
rect 930 418 1017 430
rect 830 396 834 418
rect 778 384 834 396
rect 868 396 896 418
rect 868 384 924 396
rect 958 384 1017 418
rect 323 323 1017 384
rect 1079 966 1151 1022
rect 1079 932 1098 966
rect 1132 932 1151 966
rect 1079 876 1151 932
rect 1079 842 1098 876
rect 1132 842 1151 876
rect 1079 786 1151 842
rect 1079 752 1098 786
rect 1132 752 1151 786
rect 1079 696 1151 752
rect 1079 662 1098 696
rect 1132 662 1151 696
rect 1079 606 1151 662
rect 1079 572 1098 606
rect 1132 572 1151 606
rect 1079 516 1151 572
rect 1079 482 1098 516
rect 1132 482 1151 516
rect 1079 426 1151 482
rect 1079 392 1098 426
rect 1132 392 1151 426
rect 1079 336 1151 392
rect 189 261 261 321
rect 1079 302 1098 336
rect 1132 302 1151 336
rect 1079 261 1151 302
rect 189 242 1151 261
rect 189 208 286 242
rect 320 208 376 242
rect 410 208 466 242
rect 500 208 556 242
rect 590 208 646 242
rect 680 208 736 242
rect 770 208 826 242
rect 860 208 916 242
rect 950 208 1006 242
rect 1040 208 1151 242
rect 189 189 1151 208
rect 1215 1132 1247 1166
rect 1281 1132 1314 1166
rect 1215 1076 1314 1132
rect 1215 1042 1247 1076
rect 1281 1042 1314 1076
rect 1215 986 1314 1042
rect 1215 952 1247 986
rect 1281 952 1314 986
rect 1215 896 1314 952
rect 1215 862 1247 896
rect 1281 862 1314 896
rect 1215 806 1314 862
rect 1215 772 1247 806
rect 1281 772 1314 806
rect 1215 716 1314 772
rect 1215 682 1247 716
rect 1281 682 1314 716
rect 1215 626 1314 682
rect 1215 592 1247 626
rect 1281 592 1314 626
rect 1215 536 1314 592
rect 1215 502 1247 536
rect 1281 502 1314 536
rect 1215 446 1314 502
rect 1215 412 1247 446
rect 1281 412 1314 446
rect 1215 356 1314 412
rect 1215 322 1247 356
rect 1281 322 1314 356
rect 1215 266 1314 322
rect 1215 232 1247 266
rect 1281 232 1314 266
rect 26 142 60 176
rect 94 142 125 176
rect 26 125 125 142
rect 1215 176 1314 232
rect 1215 142 1247 176
rect 1281 142 1314 176
rect 1215 125 1314 142
rect 26 92 1314 125
rect 26 58 156 92
rect 190 58 246 92
rect 280 58 336 92
rect 370 58 426 92
rect 460 58 516 92
rect 550 58 606 92
rect 640 58 696 92
rect 730 58 786 92
rect 820 58 876 92
rect 910 58 966 92
rect 1000 58 1056 92
rect 1090 58 1146 92
rect 1180 58 1314 92
rect 26 26 1314 58
<< viali >>
rect 396 924 418 930
rect 418 924 430 930
rect 496 924 508 930
rect 508 924 530 930
rect 596 924 598 930
rect 598 924 630 930
rect 396 896 430 924
rect 496 896 530 924
rect 596 896 630 924
rect 696 896 730 930
rect 796 896 830 930
rect 896 924 924 930
rect 924 924 930 930
rect 896 896 930 924
rect 396 796 430 830
rect 496 796 530 830
rect 596 796 630 830
rect 696 796 730 830
rect 796 796 830 830
rect 896 796 930 830
rect 396 696 430 730
rect 496 696 530 730
rect 596 696 630 730
rect 696 696 730 730
rect 796 696 830 730
rect 896 696 930 730
rect 396 598 430 630
rect 496 598 530 630
rect 596 598 630 630
rect 396 596 418 598
rect 418 596 430 598
rect 496 596 508 598
rect 508 596 530 598
rect 596 596 598 598
rect 598 596 630 598
rect 696 596 730 630
rect 796 596 830 630
rect 896 598 930 630
rect 896 596 924 598
rect 924 596 930 598
rect 396 508 430 530
rect 496 508 530 530
rect 596 508 630 530
rect 396 496 418 508
rect 418 496 430 508
rect 496 496 508 508
rect 508 496 530 508
rect 596 496 598 508
rect 598 496 630 508
rect 696 496 730 530
rect 796 496 830 530
rect 896 508 930 530
rect 896 496 924 508
rect 924 496 930 508
rect 396 418 430 430
rect 496 418 530 430
rect 596 418 630 430
rect 396 396 418 418
rect 418 396 430 418
rect 496 396 508 418
rect 508 396 530 418
rect 596 396 598 418
rect 598 396 630 418
rect 696 396 730 430
rect 796 396 830 430
rect 896 418 930 430
rect 896 396 924 418
rect 924 396 930 418
<< metal1 >>
rect 365 930 975 975
rect 365 896 396 930
rect 430 896 496 930
rect 530 896 596 930
rect 630 896 696 930
rect 730 896 796 930
rect 830 896 896 930
rect 930 896 975 930
rect 365 830 975 896
rect 365 796 396 830
rect 430 796 496 830
rect 530 796 596 830
rect 630 796 696 830
rect 730 796 796 830
rect 830 796 896 830
rect 930 796 975 830
rect 365 730 975 796
rect 365 696 396 730
rect 430 696 496 730
rect 530 696 596 730
rect 630 696 696 730
rect 730 696 796 730
rect 830 696 896 730
rect 930 696 975 730
rect 365 630 975 696
rect 365 596 396 630
rect 430 596 496 630
rect 530 596 596 630
rect 630 596 696 630
rect 730 596 796 630
rect 830 596 896 630
rect 930 596 975 630
rect 365 530 975 596
rect 365 496 396 530
rect 430 496 496 530
rect 530 496 596 530
rect 630 496 696 530
rect 730 496 796 530
rect 830 496 896 530
rect 930 496 975 530
rect 365 430 975 496
rect 365 396 396 430
rect 430 396 496 430
rect 530 396 596 430
rect 630 396 696 430
rect 730 396 796 430
rect 830 396 896 430
rect 930 396 975 430
rect 365 365 975 396
<< labels >>
flabel locali s 554 626 802 730 0 FreeSans 400 0 0 0 Emitter
port 1 nsew
flabel locali s 613 1252 714 1301 0 FreeSans 400 0 0 0 Collector
port 2 nsew
flabel locali s 590 1102 708 1142 0 FreeSans 400 0 0 0 Base
port 3 nsew
<< properties >>
string gencell sky130_fd_pr__rf_pnp_05v5_W3p40L3p40
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 10482778
string GDS_START 10454444
string parameter m=1
string library sky130
<< end >>
