magic
tech sky130A
magscale 1 2
timestamp 1640697996
<< nwell >>
rect -66 377 1698 897
<< pwell >>
rect 1191 217 1628 283
rect 45 43 1628 217
rect -26 -43 1658 43
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1632 831
rect 108 735 286 741
rect 142 701 180 735
rect 214 701 252 735
rect 108 451 286 701
rect 378 735 568 741
rect 378 701 384 735
rect 418 701 456 735
rect 490 701 528 735
rect 562 701 568 735
rect 378 599 568 701
rect 108 235 174 345
rect 505 359 620 493
rect 1054 735 1244 741
rect 1054 701 1060 735
rect 1094 701 1132 735
rect 1166 701 1204 735
rect 1238 701 1244 735
rect 1054 579 1244 701
rect 1307 735 1497 751
rect 1307 701 1313 735
rect 1347 701 1385 735
rect 1419 701 1457 735
rect 1491 701 1497 735
rect 169 113 359 199
rect 169 79 175 113
rect 209 79 247 113
rect 281 79 319 113
rect 353 79 359 113
rect 1307 507 1497 701
rect 481 113 599 195
rect 169 73 359 79
rect 481 79 487 113
rect 521 79 559 113
rect 593 79 599 113
rect 1054 113 1172 179
rect 481 73 599 79
rect 1054 79 1060 113
rect 1094 79 1132 113
rect 1166 79 1172 113
rect 1054 73 1172 79
rect 1311 113 1501 249
rect 1311 79 1317 113
rect 1351 79 1389 113
rect 1423 79 1461 113
rect 1495 79 1501 113
rect 1540 103 1610 751
rect 1311 73 1501 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 108 701 142 735
rect 180 701 214 735
rect 252 701 286 735
rect 384 701 418 735
rect 456 701 490 735
rect 528 701 562 735
rect 1060 701 1094 735
rect 1132 701 1166 735
rect 1204 701 1238 735
rect 1313 701 1347 735
rect 1385 701 1419 735
rect 1457 701 1491 735
rect 175 79 209 113
rect 247 79 281 113
rect 319 79 353 113
rect 487 79 521 113
rect 559 79 593 113
rect 1060 79 1094 113
rect 1132 79 1166 113
rect 1317 79 1351 113
rect 1389 79 1423 113
rect 1461 79 1495 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< obsli1 >>
rect 22 415 72 597
rect 604 727 810 761
rect 604 563 638 727
rect 322 529 638 563
rect 674 579 740 691
rect 322 415 356 529
rect 392 439 458 493
rect 22 403 356 415
rect 22 381 359 403
rect 22 199 72 381
rect 308 269 359 381
rect 395 323 458 439
rect 674 467 708 579
rect 776 543 810 727
rect 846 613 896 745
rect 846 579 1018 613
rect 744 503 948 543
rect 674 433 846 467
rect 710 323 776 397
rect 395 289 776 323
rect 22 99 133 199
rect 395 103 445 289
rect 812 253 846 433
rect 677 219 846 253
rect 882 219 948 503
rect 984 401 1018 579
rect 1205 471 1271 535
rect 1205 437 1406 471
rect 984 367 1336 401
rect 677 199 711 219
rect 645 99 711 199
rect 984 183 1018 367
rect 1270 355 1336 367
rect 1086 319 1152 331
rect 1372 319 1406 437
rect 1086 285 1406 319
rect 1086 215 1152 285
rect 801 149 1018 183
rect 801 99 867 149
rect 1209 169 1275 285
<< metal1 >>
rect 0 831 1632 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1632 831
rect 0 791 1632 797
rect 0 735 1632 763
rect 0 701 108 735
rect 142 701 180 735
rect 214 701 252 735
rect 286 701 384 735
rect 418 701 456 735
rect 490 701 528 735
rect 562 701 1060 735
rect 1094 701 1132 735
rect 1166 701 1204 735
rect 1238 701 1313 735
rect 1347 701 1385 735
rect 1419 701 1457 735
rect 1491 701 1632 735
rect 0 689 1632 701
rect 0 113 1632 125
rect 0 79 175 113
rect 209 79 247 113
rect 281 79 319 113
rect 353 79 487 113
rect 521 79 559 113
rect 593 79 1060 113
rect 1094 79 1132 113
rect 1166 79 1317 113
rect 1351 79 1389 113
rect 1423 79 1461 113
rect 1495 79 1632 113
rect 0 51 1632 79
rect 0 17 1632 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -23 1632 -17
<< labels >>
rlabel locali s 505 359 620 493 6 D
port 1 nsew signal input
rlabel locali s 108 235 174 345 6 GATE
port 2 nsew clock input
rlabel metal1 s 0 51 1632 125 6 VGND
port 3 nsew ground bidirectional
rlabel viali s 559 79 593 113 6 VGND
port 3 nsew ground bidirectional
rlabel viali s 487 79 521 113 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 481 73 599 195 6 VGND
port 3 nsew ground bidirectional
rlabel viali s 1132 79 1166 113 6 VGND
port 3 nsew ground bidirectional
rlabel viali s 1060 79 1094 113 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 1054 73 1172 179 6 VGND
port 3 nsew ground bidirectional
rlabel viali s 1461 79 1495 113 6 VGND
port 3 nsew ground bidirectional
rlabel viali s 1389 79 1423 113 6 VGND
port 3 nsew ground bidirectional
rlabel viali s 1317 79 1351 113 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 1311 73 1501 249 6 VGND
port 3 nsew ground bidirectional
rlabel viali s 319 79 353 113 6 VGND
port 3 nsew ground bidirectional
rlabel viali s 247 79 281 113 6 VGND
port 3 nsew ground bidirectional
rlabel viali s 175 79 209 113 6 VGND
port 3 nsew ground bidirectional
rlabel locali s 169 73 359 199 6 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 -23 1632 23 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s -26 -43 1658 43 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s 45 43 1628 217 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1191 217 1628 283 6 VNB
port 4 nsew ground bidirectional
rlabel viali s 1567 -17 1601 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 1471 -17 1505 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 1375 -17 1409 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 1279 -17 1313 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 1183 -17 1217 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 1087 -17 1121 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 991 -17 1025 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 895 -17 929 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 799 -17 833 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 703 -17 737 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 607 -17 641 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 511 -17 545 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 415 -17 449 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 319 -17 353 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 223 -17 257 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 127 -17 161 17 8 VNB
port 4 nsew ground bidirectional
rlabel viali s 31 -17 65 17 8 VNB
port 4 nsew ground bidirectional
rlabel locali s 0 -17 1632 17 8 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 791 1632 837 6 VPB
port 5 nsew power bidirectional
rlabel nwell s -66 377 1698 897 6 VPB
port 5 nsew power bidirectional
rlabel viali s 1567 797 1601 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 1471 797 1505 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 1375 797 1409 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 1279 797 1313 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 1183 797 1217 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 1087 797 1121 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 991 797 1025 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 895 797 929 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 799 797 833 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 703 797 737 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 607 797 641 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 511 797 545 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 415 797 449 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 319 797 353 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 223 797 257 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 127 797 161 831 6 VPB
port 5 nsew power bidirectional
rlabel viali s 31 797 65 831 6 VPB
port 5 nsew power bidirectional
rlabel locali s 0 797 1632 831 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 689 1632 763 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 528 701 562 735 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 456 701 490 735 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 384 701 418 735 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 378 599 568 741 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1204 701 1238 735 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1132 701 1166 735 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1060 701 1094 735 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 1054 579 1244 741 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1457 701 1491 735 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1385 701 1419 735 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 1313 701 1347 735 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 1307 507 1497 751 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 252 701 286 735 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 180 701 214 735 6 VPWR
port 6 nsew power bidirectional
rlabel viali s 108 701 142 735 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 108 451 286 741 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 1540 103 1610 751 6 Q
port 7 nsew signal output
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 1632 814
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_END 1220156
string GDS_START 1203716
<< end >>
