magic
tech sky130A
magscale 1 2
timestamp 1619729571
<< checkpaint >>
rect -1298 -1308 2770 1852
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 85 47 115 177
rect 169 47 199 177
rect 253 47 283 177
rect 337 47 367 177
rect 421 47 451 177
rect 505 47 535 177
rect 589 47 619 177
rect 673 47 703 177
rect 767 47 797 177
rect 851 47 881 177
rect 935 47 965 177
rect 1019 47 1049 177
rect 1103 47 1133 177
rect 1187 47 1217 177
rect 1271 47 1301 177
rect 1355 47 1385 177
<< scpmoshvt >>
rect 85 297 115 497
rect 169 297 199 497
rect 253 297 283 497
rect 337 297 367 497
rect 421 297 451 497
rect 505 297 535 497
rect 589 297 619 497
rect 673 297 703 497
rect 767 297 797 497
rect 851 297 881 497
rect 935 297 965 497
rect 1019 297 1049 497
rect 1103 297 1133 497
rect 1187 297 1217 497
rect 1271 297 1301 497
rect 1355 297 1385 497
<< ndiff >>
rect 33 163 85 177
rect 33 129 41 163
rect 75 129 85 163
rect 33 95 85 129
rect 33 61 41 95
rect 75 61 85 95
rect 33 47 85 61
rect 115 95 169 177
rect 115 61 125 95
rect 159 61 169 95
rect 115 47 169 61
rect 199 163 253 177
rect 199 129 209 163
rect 243 129 253 163
rect 199 95 253 129
rect 199 61 209 95
rect 243 61 253 95
rect 199 47 253 61
rect 283 95 337 177
rect 283 61 293 95
rect 327 61 337 95
rect 283 47 337 61
rect 367 163 421 177
rect 367 129 377 163
rect 411 129 421 163
rect 367 95 421 129
rect 367 61 377 95
rect 411 61 421 95
rect 367 47 421 61
rect 451 95 505 177
rect 451 61 461 95
rect 495 61 505 95
rect 451 47 505 61
rect 535 163 589 177
rect 535 129 545 163
rect 579 129 589 163
rect 535 95 589 129
rect 535 61 545 95
rect 579 61 589 95
rect 535 47 589 61
rect 619 95 673 177
rect 619 61 629 95
rect 663 61 673 95
rect 619 47 673 61
rect 703 163 767 177
rect 703 129 713 163
rect 747 129 767 163
rect 703 95 767 129
rect 703 61 713 95
rect 747 61 767 95
rect 703 47 767 61
rect 797 163 851 177
rect 797 129 807 163
rect 841 129 851 163
rect 797 47 851 129
rect 881 95 935 177
rect 881 61 891 95
rect 925 61 935 95
rect 881 47 935 61
rect 965 163 1019 177
rect 965 129 975 163
rect 1009 129 1019 163
rect 965 47 1019 129
rect 1049 95 1103 177
rect 1049 61 1059 95
rect 1093 61 1103 95
rect 1049 47 1103 61
rect 1133 163 1187 177
rect 1133 129 1143 163
rect 1177 129 1187 163
rect 1133 47 1187 129
rect 1217 95 1271 177
rect 1217 61 1227 95
rect 1261 61 1271 95
rect 1217 47 1271 61
rect 1301 163 1355 177
rect 1301 129 1311 163
rect 1345 129 1355 163
rect 1301 47 1355 129
rect 1385 95 1437 177
rect 1385 61 1395 95
rect 1429 61 1437 95
rect 1385 47 1437 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 41 477
rect 75 443 85 477
rect 27 409 85 443
rect 27 375 41 409
rect 75 375 85 409
rect 27 341 85 375
rect 27 307 41 341
rect 75 307 85 341
rect 27 297 85 307
rect 115 477 169 497
rect 115 443 125 477
rect 159 443 169 477
rect 115 409 169 443
rect 115 375 125 409
rect 159 375 169 409
rect 115 341 169 375
rect 115 307 125 341
rect 159 307 169 341
rect 115 297 169 307
rect 199 477 253 497
rect 199 443 209 477
rect 243 443 253 477
rect 199 297 253 443
rect 283 477 337 497
rect 283 443 293 477
rect 327 443 337 477
rect 283 409 337 443
rect 283 375 293 409
rect 327 375 337 409
rect 283 297 337 375
rect 367 409 421 497
rect 367 375 377 409
rect 411 375 421 409
rect 367 297 421 375
rect 451 477 505 497
rect 451 443 461 477
rect 495 443 505 477
rect 451 297 505 443
rect 535 409 589 497
rect 535 375 545 409
rect 579 375 589 409
rect 535 297 589 375
rect 619 477 673 497
rect 619 443 629 477
rect 663 443 673 477
rect 619 297 673 443
rect 703 477 767 497
rect 703 443 721 477
rect 755 443 767 477
rect 703 297 767 443
rect 797 477 851 497
rect 797 443 807 477
rect 841 443 851 477
rect 797 297 851 443
rect 881 477 935 497
rect 881 443 891 477
rect 925 443 935 477
rect 881 297 935 443
rect 965 477 1019 497
rect 965 443 975 477
rect 1009 443 1019 477
rect 965 409 1019 443
rect 965 375 975 409
rect 1009 375 1019 409
rect 965 297 1019 375
rect 1049 409 1103 497
rect 1049 375 1059 409
rect 1093 375 1103 409
rect 1049 297 1103 375
rect 1133 477 1187 497
rect 1133 443 1143 477
rect 1177 443 1187 477
rect 1133 297 1187 443
rect 1217 409 1271 497
rect 1217 375 1227 409
rect 1261 375 1271 409
rect 1217 297 1271 375
rect 1301 477 1355 497
rect 1301 443 1311 477
rect 1345 443 1355 477
rect 1301 297 1355 443
rect 1385 477 1437 497
rect 1385 443 1395 477
rect 1429 443 1437 477
rect 1385 297 1437 443
<< ndiffc >>
rect 41 129 75 163
rect 41 61 75 95
rect 125 61 159 95
rect 209 129 243 163
rect 209 61 243 95
rect 293 61 327 95
rect 377 129 411 163
rect 377 61 411 95
rect 461 61 495 95
rect 545 129 579 163
rect 545 61 579 95
rect 629 61 663 95
rect 713 129 747 163
rect 713 61 747 95
rect 807 129 841 163
rect 891 61 925 95
rect 975 129 1009 163
rect 1059 61 1093 95
rect 1143 129 1177 163
rect 1227 61 1261 95
rect 1311 129 1345 163
rect 1395 61 1429 95
<< pdiffc >>
rect 41 443 75 477
rect 41 375 75 409
rect 41 307 75 341
rect 125 443 159 477
rect 125 375 159 409
rect 125 307 159 341
rect 209 443 243 477
rect 293 443 327 477
rect 293 375 327 409
rect 377 375 411 409
rect 461 443 495 477
rect 545 375 579 409
rect 629 443 663 477
rect 721 443 755 477
rect 807 443 841 477
rect 891 443 925 477
rect 975 443 1009 477
rect 975 375 1009 409
rect 1059 375 1093 409
rect 1143 443 1177 477
rect 1227 375 1261 409
rect 1311 443 1345 477
rect 1395 443 1429 477
<< poly >>
rect 85 497 115 523
rect 169 497 199 523
rect 253 497 283 523
rect 337 497 367 523
rect 421 497 451 523
rect 505 497 535 523
rect 589 497 619 523
rect 673 497 703 523
rect 767 497 797 523
rect 851 497 881 523
rect 935 497 965 523
rect 1019 497 1049 523
rect 1103 497 1133 523
rect 1187 497 1217 523
rect 1271 497 1301 523
rect 1355 497 1385 523
rect 85 265 115 297
rect 169 265 199 297
rect 253 265 283 297
rect 76 249 283 265
rect 76 215 97 249
rect 131 215 165 249
rect 199 215 233 249
rect 267 215 283 249
rect 76 199 283 215
rect 85 177 115 199
rect 169 177 199 199
rect 253 177 283 199
rect 337 265 367 297
rect 421 265 451 297
rect 505 265 535 297
rect 589 265 619 297
rect 673 265 703 297
rect 767 265 797 297
rect 851 265 881 297
rect 935 265 965 297
rect 1019 265 1049 297
rect 1103 265 1133 297
rect 1187 265 1217 297
rect 1271 265 1301 297
rect 1355 265 1385 297
rect 337 249 619 265
rect 337 215 365 249
rect 399 215 433 249
rect 467 215 501 249
rect 535 215 569 249
rect 603 215 619 249
rect 337 199 619 215
rect 661 249 715 265
rect 661 215 671 249
rect 705 215 715 249
rect 661 199 715 215
rect 767 249 977 265
rect 767 215 859 249
rect 893 215 927 249
rect 961 215 977 249
rect 767 199 977 215
rect 1019 249 1301 265
rect 1019 215 1038 249
rect 1072 215 1106 249
rect 1140 215 1174 249
rect 1208 215 1242 249
rect 1276 215 1301 249
rect 1019 199 1301 215
rect 1343 249 1403 265
rect 1343 215 1353 249
rect 1387 215 1403 249
rect 1343 199 1403 215
rect 337 177 367 199
rect 421 177 451 199
rect 505 177 535 199
rect 589 177 619 199
rect 673 177 703 199
rect 767 177 797 199
rect 851 177 881 199
rect 935 177 965 199
rect 1019 177 1049 199
rect 1103 177 1133 199
rect 1187 177 1217 199
rect 1271 177 1301 199
rect 1355 177 1385 199
rect 85 21 115 47
rect 169 21 199 47
rect 253 21 283 47
rect 337 21 367 47
rect 421 21 451 47
rect 505 21 535 47
rect 589 21 619 47
rect 673 21 703 47
rect 767 21 797 47
rect 851 21 881 47
rect 935 21 965 47
rect 1019 21 1049 47
rect 1103 21 1133 47
rect 1187 21 1217 47
rect 1271 21 1301 47
rect 1355 21 1385 47
<< polycont >>
rect 97 215 131 249
rect 165 215 199 249
rect 233 215 267 249
rect 365 215 399 249
rect 433 215 467 249
rect 501 215 535 249
rect 569 215 603 249
rect 671 215 705 249
rect 859 215 893 249
rect 927 215 961 249
rect 1038 215 1072 249
rect 1106 215 1140 249
rect 1174 215 1208 249
rect 1242 215 1276 249
rect 1353 215 1387 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 33 477 83 527
rect 33 443 41 477
rect 75 443 83 477
rect 33 409 83 443
rect 33 375 41 409
rect 75 375 83 409
rect 33 341 83 375
rect 33 307 41 341
rect 75 307 83 341
rect 33 289 83 307
rect 117 477 167 493
rect 117 443 125 477
rect 159 443 167 477
rect 117 409 167 443
rect 201 477 251 527
rect 201 443 209 477
rect 243 443 251 477
rect 201 425 251 443
rect 285 477 679 493
rect 285 443 293 477
rect 327 459 461 477
rect 327 443 335 459
rect 117 375 125 409
rect 159 391 167 409
rect 285 409 335 443
rect 453 443 461 459
rect 495 459 629 477
rect 495 443 503 459
rect 453 425 503 443
rect 621 443 629 459
rect 663 443 679 477
rect 621 425 679 443
rect 713 477 757 527
rect 713 443 721 477
rect 755 443 757 477
rect 713 425 757 443
rect 791 477 851 493
rect 791 443 807 477
rect 841 443 851 477
rect 791 425 851 443
rect 885 477 933 527
rect 885 443 891 477
rect 925 443 933 477
rect 885 425 933 443
rect 967 477 1353 493
rect 967 443 975 477
rect 1009 459 1143 477
rect 1009 443 1017 459
rect 285 391 293 409
rect 159 375 293 391
rect 327 375 335 409
rect 117 357 335 375
rect 369 409 419 425
rect 369 375 377 409
rect 411 391 419 409
rect 537 409 587 425
rect 537 391 545 409
rect 411 375 545 391
rect 579 391 587 409
rect 817 391 851 425
rect 967 409 1017 443
rect 1135 443 1143 459
rect 1177 459 1311 477
rect 1177 443 1185 459
rect 1135 425 1185 443
rect 1303 443 1311 459
rect 1345 443 1353 477
rect 1303 427 1353 443
rect 1387 477 1443 527
rect 1387 443 1395 477
rect 1429 443 1443 477
rect 1387 425 1443 443
rect 967 391 975 409
rect 579 375 783 391
rect 369 357 783 375
rect 817 375 975 391
rect 1009 375 1017 409
rect 817 357 1017 375
rect 1051 409 1101 425
rect 1051 375 1059 409
rect 1093 391 1101 409
rect 1219 409 1269 425
rect 1219 391 1227 409
rect 1093 375 1227 391
rect 1261 391 1269 409
rect 1261 375 1455 391
rect 1051 357 1455 375
rect 117 341 167 357
rect 117 307 125 341
rect 159 307 167 341
rect 749 323 783 357
rect 117 289 167 307
rect 230 289 715 323
rect 749 289 825 323
rect 230 255 283 289
rect 17 249 283 255
rect 17 215 97 249
rect 131 215 165 249
rect 199 215 233 249
rect 267 215 283 249
rect 337 249 619 255
rect 337 215 365 249
rect 399 215 433 249
rect 467 215 501 249
rect 535 215 569 249
rect 603 215 619 249
rect 655 249 715 289
rect 655 215 671 249
rect 705 215 721 249
rect 25 163 757 181
rect 25 129 41 163
rect 75 145 209 163
rect 75 129 91 145
rect 25 95 91 129
rect 193 129 209 145
rect 243 147 377 163
rect 243 129 259 147
rect 25 61 41 95
rect 75 61 91 95
rect 25 51 91 61
rect 125 95 159 111
rect 125 17 159 61
rect 193 95 259 129
rect 361 129 377 147
rect 411 145 545 163
rect 411 129 427 145
rect 193 61 209 95
rect 243 61 259 95
rect 193 51 259 61
rect 293 95 327 111
rect 293 17 327 61
rect 361 95 427 129
rect 529 129 545 145
rect 579 147 713 163
rect 579 129 595 147
rect 361 61 377 95
rect 411 61 427 95
rect 361 51 427 61
rect 461 95 495 111
rect 461 17 495 61
rect 529 95 595 129
rect 697 129 713 147
rect 747 129 757 163
rect 791 164 825 289
rect 859 289 1387 323
rect 859 249 988 289
rect 893 215 927 249
rect 961 215 988 249
rect 1022 249 1292 255
rect 1022 215 1038 249
rect 1072 215 1106 249
rect 1140 215 1174 249
rect 1208 215 1242 249
rect 1276 215 1292 249
rect 1343 249 1387 289
rect 1343 215 1353 249
rect 859 199 988 215
rect 1343 199 1387 215
rect 1421 164 1455 357
rect 791 163 1455 164
rect 791 129 807 163
rect 841 129 975 163
rect 1009 129 1143 163
rect 1177 129 1311 163
rect 1345 129 1455 163
rect 529 61 545 95
rect 579 61 595 95
rect 529 51 595 61
rect 629 95 663 111
rect 629 17 663 61
rect 697 95 757 129
rect 697 61 713 95
rect 747 61 891 95
rect 925 61 1059 95
rect 1093 61 1227 95
rect 1261 61 1395 95
rect 1429 61 1449 95
rect 697 51 1449 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 581 357 615 391 0 FreeSans 400 0 0 0 Y
port 9 nsew signal output
flabel locali s 489 221 523 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 949 221 983 255 0 FreeSans 400 180 0 0 B1
port 3 nsew signal input
flabel locali s 1225 221 1259 255 0 FreeSans 400 180 0 0 B2
port 4 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o22ai_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 2943764
string GDS_START 2933160
string path 0.000 0.000 36.800 0.000 
<< end >>
