magic
tech sky130A
timestamp 1619729433
<< properties >>
string gencell sky130_fd_pr__rf_test_coil2
string parameter m=1
string library sky130
<< end >>
