magic
tech sky130A
magscale 1 2
timestamp 1640697977
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 643 203
rect 27 -17 61 21
<< scnmos >>
rect 80 47 110 177
rect 270 47 300 177
rect 356 47 386 177
rect 442 47 472 177
rect 534 47 564 177
<< scpmoshvt >>
rect 80 297 110 497
rect 270 297 300 497
rect 356 297 386 497
rect 442 297 472 497
rect 534 297 564 497
<< ndiff >>
rect 27 165 80 177
rect 27 131 35 165
rect 69 131 80 165
rect 27 97 80 131
rect 27 63 35 97
rect 69 63 80 97
rect 27 47 80 63
rect 110 89 270 177
rect 110 55 137 89
rect 171 55 209 89
rect 243 55 270 89
rect 110 47 270 55
rect 300 47 356 177
rect 386 123 442 177
rect 386 89 397 123
rect 431 89 442 123
rect 386 47 442 89
rect 472 89 534 177
rect 472 55 486 89
rect 520 55 534 89
rect 472 47 534 55
rect 564 123 617 177
rect 564 89 575 123
rect 609 89 617 123
rect 564 47 617 89
<< pdiff >>
rect 27 475 80 497
rect 27 441 35 475
rect 69 441 80 475
rect 27 347 80 441
rect 27 313 35 347
rect 69 313 80 347
rect 27 297 80 313
rect 110 485 163 497
rect 110 451 121 485
rect 155 451 163 485
rect 110 417 163 451
rect 110 383 121 417
rect 155 383 163 417
rect 110 297 163 383
rect 217 475 270 497
rect 217 441 225 475
rect 259 441 270 475
rect 217 407 270 441
rect 217 373 225 407
rect 259 373 270 407
rect 217 297 270 373
rect 300 489 356 497
rect 300 455 311 489
rect 345 455 356 489
rect 300 297 356 455
rect 386 475 442 497
rect 386 441 397 475
rect 431 441 442 475
rect 386 407 442 441
rect 386 373 397 407
rect 431 373 442 407
rect 386 297 442 373
rect 472 297 534 497
rect 564 461 617 497
rect 564 427 575 461
rect 609 427 617 461
rect 564 387 617 427
rect 564 353 575 387
rect 609 353 617 387
rect 564 297 617 353
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 137 55 171 89
rect 209 55 243 89
rect 397 89 431 123
rect 486 55 520 89
rect 575 89 609 123
<< pdiffc >>
rect 35 441 69 475
rect 35 313 69 347
rect 121 451 155 485
rect 121 383 155 417
rect 225 441 259 475
rect 225 373 259 407
rect 311 455 345 489
rect 397 441 431 475
rect 397 373 431 407
rect 575 427 609 461
rect 575 353 609 387
<< poly >>
rect 80 497 110 523
rect 270 497 300 523
rect 356 497 386 523
rect 442 497 472 523
rect 534 497 564 523
rect 80 265 110 297
rect 270 265 300 297
rect 356 265 386 297
rect 442 265 472 297
rect 534 265 564 297
rect 80 249 164 265
rect 80 215 120 249
rect 154 215 164 249
rect 80 199 164 215
rect 216 249 300 265
rect 216 215 226 249
rect 260 215 300 249
rect 216 199 300 215
rect 342 249 396 265
rect 342 215 352 249
rect 386 215 396 249
rect 342 199 396 215
rect 438 249 492 265
rect 438 215 448 249
rect 482 215 492 249
rect 438 199 492 215
rect 534 249 618 265
rect 534 215 574 249
rect 608 215 618 249
rect 534 199 618 215
rect 80 177 110 199
rect 270 177 300 199
rect 356 177 386 199
rect 442 177 472 199
rect 534 177 564 199
rect 80 21 110 47
rect 270 21 300 47
rect 356 21 386 47
rect 442 21 472 47
rect 534 21 564 47
<< polycont >>
rect 120 215 154 249
rect 226 215 260 249
rect 352 215 386 249
rect 448 215 482 249
rect 574 215 608 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 18 475 71 491
rect 18 441 35 475
rect 69 441 71 475
rect 18 347 71 441
rect 105 485 171 527
rect 105 451 121 485
rect 155 451 171 485
rect 105 417 171 451
rect 105 383 121 417
rect 155 383 171 417
rect 209 475 261 491
rect 209 441 225 475
rect 259 441 261 475
rect 295 489 361 527
rect 295 455 311 489
rect 345 455 361 489
rect 295 453 361 455
rect 395 475 447 491
rect 209 419 261 441
rect 395 441 397 475
rect 431 441 447 475
rect 395 419 447 441
rect 209 407 447 419
rect 209 373 225 407
rect 259 373 397 407
rect 431 373 447 407
rect 561 461 619 491
rect 561 427 575 461
rect 609 427 619 461
rect 561 387 619 427
rect 18 313 35 347
rect 69 337 71 347
rect 561 353 575 387
rect 609 353 619 387
rect 561 337 619 353
rect 69 313 85 337
rect 18 165 85 313
rect 18 131 35 165
rect 69 131 85 165
rect 18 97 85 131
rect 120 301 619 337
rect 120 249 165 301
rect 154 215 165 249
rect 120 163 165 215
rect 205 249 261 265
rect 205 215 226 249
rect 260 215 261 249
rect 205 199 261 215
rect 297 249 412 265
rect 297 215 352 249
rect 386 215 412 249
rect 297 199 412 215
rect 448 249 535 265
rect 482 215 535 249
rect 448 199 535 215
rect 571 249 625 265
rect 571 215 574 249
rect 608 215 625 249
rect 571 199 625 215
rect 120 125 617 163
rect 18 63 35 97
rect 69 63 85 97
rect 383 123 434 125
rect 18 53 85 63
rect 121 89 270 91
rect 121 55 137 89
rect 171 55 209 89
rect 243 55 270 89
rect 121 17 270 55
rect 383 89 397 123
rect 431 89 434 123
rect 572 123 617 125
rect 383 53 434 89
rect 470 89 536 91
rect 470 55 486 89
rect 520 55 536 89
rect 470 17 536 55
rect 572 89 575 123
rect 609 89 617 123
rect 572 53 617 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel pwell s 27 -17 61 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 27 527 61 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 27 -17 61 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 27 527 61 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 27 425 61 459 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 27 85 61 119 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 215 221 249 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 27 357 61 391 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 491 221 525 255 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 27 221 61 255 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 307 221 341 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 27 153 61 187 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 27 289 61 323 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 583 221 617 255 0 FreeSans 200 0 0 0 C1
port 4 nsew signal input
rlabel comment s 0 0 0 0 4 a211o_1
rlabel metal1 s 0 -48 644 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 3634700
string GDS_START 3628354
string path 0.000 0.000 16.100 0.000 
<< end >>
