magic
tech sky130A
magscale 1 2
timestamp 1619729571
<< checkpaint >>
rect -1298 -1308 2402 1852
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 85 47 115 177
rect 171 47 201 177
rect 257 47 287 177
rect 365 47 395 177
rect 460 47 490 177
rect 568 47 598 177
rect 654 47 684 177
rect 794 47 824 177
rect 893 47 923 177
rect 979 47 1009 177
<< scpmoshvt >>
rect 85 297 115 497
rect 171 297 201 497
rect 257 297 287 497
rect 343 297 373 497
rect 437 297 467 497
rect 523 297 553 497
rect 713 297 743 497
rect 799 297 829 497
rect 885 297 915 497
rect 979 297 1009 497
<< ndiff >>
rect 28 169 85 177
rect 28 135 40 169
rect 74 135 85 169
rect 28 101 85 135
rect 28 67 40 101
rect 74 67 85 101
rect 28 47 85 67
rect 115 89 171 177
rect 115 55 126 89
rect 160 55 171 89
rect 115 47 171 55
rect 201 169 257 177
rect 201 135 212 169
rect 246 135 257 169
rect 201 101 257 135
rect 201 67 212 101
rect 246 67 257 101
rect 201 47 257 67
rect 287 89 365 177
rect 287 55 309 89
rect 343 55 365 89
rect 287 47 365 55
rect 395 165 460 177
rect 395 131 409 165
rect 443 131 460 165
rect 395 97 460 131
rect 395 63 409 97
rect 443 63 460 97
rect 395 47 460 63
rect 490 89 568 177
rect 490 55 509 89
rect 543 55 568 89
rect 490 47 568 55
rect 598 165 654 177
rect 598 131 609 165
rect 643 131 654 165
rect 598 92 654 131
rect 598 58 609 92
rect 643 58 654 92
rect 598 47 654 58
rect 684 47 794 177
rect 824 89 893 177
rect 824 55 841 89
rect 875 55 893 89
rect 824 47 893 55
rect 923 47 979 177
rect 1009 161 1062 177
rect 1009 127 1020 161
rect 1054 127 1062 161
rect 1009 93 1062 127
rect 1009 59 1020 93
rect 1054 59 1062 93
rect 1009 47 1062 59
<< pdiff >>
rect 28 489 85 497
rect 28 455 40 489
rect 74 455 85 489
rect 28 421 85 455
rect 28 387 40 421
rect 74 387 85 421
rect 28 297 85 387
rect 115 297 171 497
rect 201 413 257 497
rect 201 379 212 413
rect 246 379 257 413
rect 201 297 257 379
rect 287 297 343 497
rect 373 489 437 497
rect 373 455 384 489
rect 418 455 437 489
rect 373 297 437 455
rect 467 412 523 497
rect 467 378 478 412
rect 512 378 523 412
rect 467 297 523 378
rect 553 477 605 497
rect 553 443 563 477
rect 597 443 605 477
rect 553 297 605 443
rect 661 477 713 497
rect 661 443 669 477
rect 703 443 713 477
rect 661 409 713 443
rect 661 375 669 409
rect 703 375 713 409
rect 661 297 713 375
rect 743 489 799 497
rect 743 455 754 489
rect 788 455 799 489
rect 743 297 799 455
rect 829 477 885 497
rect 829 443 840 477
rect 874 443 885 477
rect 829 409 885 443
rect 829 375 840 409
rect 874 375 885 409
rect 829 297 885 375
rect 915 489 979 497
rect 915 455 930 489
rect 964 455 979 489
rect 915 297 979 455
rect 1009 489 1076 497
rect 1009 455 1030 489
rect 1064 455 1076 489
rect 1009 421 1076 455
rect 1009 387 1030 421
rect 1064 387 1076 421
rect 1009 297 1076 387
<< ndiffc >>
rect 40 135 74 169
rect 40 67 74 101
rect 126 55 160 89
rect 212 135 246 169
rect 212 67 246 101
rect 309 55 343 89
rect 409 131 443 165
rect 409 63 443 97
rect 509 55 543 89
rect 609 131 643 165
rect 609 58 643 92
rect 841 55 875 89
rect 1020 127 1054 161
rect 1020 59 1054 93
<< pdiffc >>
rect 40 455 74 489
rect 40 387 74 421
rect 212 379 246 413
rect 384 455 418 489
rect 478 378 512 412
rect 563 443 597 477
rect 669 443 703 477
rect 669 375 703 409
rect 754 455 788 489
rect 840 443 874 477
rect 840 375 874 409
rect 930 455 964 489
rect 1030 455 1064 489
rect 1030 387 1064 421
<< poly >>
rect 85 497 115 523
rect 171 497 201 523
rect 257 497 287 523
rect 343 497 373 523
rect 437 497 467 523
rect 523 497 553 523
rect 713 497 743 523
rect 799 497 829 523
rect 885 497 915 523
rect 979 497 1009 523
rect 85 265 115 297
rect 171 265 201 297
rect 257 265 287 297
rect 343 265 373 297
rect 437 265 467 297
rect 523 265 553 297
rect 713 265 743 297
rect 799 265 829 297
rect 885 265 915 297
rect 979 265 1009 297
rect 25 249 115 265
rect 25 215 41 249
rect 75 215 115 249
rect 25 199 115 215
rect 157 249 287 265
rect 157 215 167 249
rect 201 215 235 249
rect 269 215 287 249
rect 157 199 287 215
rect 329 249 395 265
rect 329 215 339 249
rect 373 215 395 249
rect 329 199 395 215
rect 437 249 598 265
rect 437 215 453 249
rect 487 215 521 249
rect 555 215 598 249
rect 437 199 598 215
rect 85 177 115 199
rect 171 177 201 199
rect 257 177 287 199
rect 365 177 395 199
rect 460 177 490 199
rect 568 177 598 199
rect 654 249 743 265
rect 654 215 693 249
rect 727 215 743 249
rect 654 199 743 215
rect 794 249 937 265
rect 794 215 819 249
rect 853 215 887 249
rect 921 215 937 249
rect 654 177 684 199
rect 794 198 937 215
rect 979 249 1045 265
rect 979 215 995 249
rect 1029 215 1045 249
rect 979 199 1045 215
rect 794 177 824 198
rect 893 177 923 198
rect 979 177 1009 199
rect 85 21 115 47
rect 171 21 201 47
rect 257 21 287 47
rect 365 21 395 47
rect 460 21 490 47
rect 568 21 598 47
rect 654 21 684 47
rect 794 21 824 47
rect 893 21 923 47
rect 979 21 1009 47
<< polycont >>
rect 41 215 75 249
rect 167 215 201 249
rect 235 215 269 249
rect 339 215 373 249
rect 453 215 487 249
rect 521 215 555 249
rect 693 215 727 249
rect 819 215 853 249
rect 887 215 921 249
rect 995 215 1029 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 20 489 597 493
rect 20 455 40 489
rect 74 455 384 489
rect 418 477 597 489
rect 418 459 563 477
rect 418 455 437 459
rect 20 421 92 455
rect 563 427 597 443
rect 631 477 704 493
rect 631 443 669 477
rect 703 443 704 477
rect 738 489 804 527
rect 738 455 754 489
rect 788 455 804 489
rect 838 477 880 493
rect 20 387 40 421
rect 74 387 92 421
rect 20 374 92 387
rect 180 413 428 421
rect 180 379 212 413
rect 246 379 428 413
rect 631 419 704 443
rect 838 443 840 477
rect 874 443 880 477
rect 914 489 980 527
rect 914 455 930 489
rect 964 455 980 489
rect 1014 489 1080 493
rect 1014 455 1030 489
rect 1064 455 1080 489
rect 838 421 880 443
rect 1014 421 1080 455
rect 838 419 1030 421
rect 180 370 428 379
rect 25 289 360 336
rect 394 325 428 370
rect 462 378 478 412
rect 512 393 528 412
rect 631 409 1030 419
rect 631 393 669 409
rect 512 378 669 393
rect 462 375 669 378
rect 703 375 840 409
rect 874 387 1030 409
rect 1064 387 1080 421
rect 874 375 1080 387
rect 462 369 1080 375
rect 462 359 667 369
rect 394 289 651 325
rect 25 249 91 289
rect 323 255 360 289
rect 25 215 41 249
rect 75 215 91 249
rect 151 249 285 255
rect 151 215 167 249
rect 201 215 235 249
rect 269 215 285 249
rect 323 249 395 255
rect 323 215 339 249
rect 373 215 395 249
rect 25 209 91 215
rect 323 206 395 215
rect 437 249 571 255
rect 437 215 453 249
rect 487 215 521 249
rect 555 215 571 249
rect 437 206 571 215
rect 605 169 651 289
rect 693 289 1058 335
rect 693 249 743 289
rect 727 215 743 249
rect 693 197 743 215
rect 794 249 945 255
rect 794 215 819 249
rect 853 215 887 249
rect 921 215 945 249
rect 794 203 945 215
rect 979 249 1058 289
rect 979 215 995 249
rect 1029 215 1058 249
rect 979 199 1058 215
rect 24 135 40 169
rect 74 135 212 169
rect 246 165 651 169
rect 246 135 409 165
rect 24 131 409 135
rect 443 131 609 165
rect 643 161 651 165
rect 643 131 1020 161
rect 24 127 1020 131
rect 1054 127 1071 161
rect 24 123 1071 127
rect 24 101 76 123
rect 24 67 40 101
rect 74 67 76 101
rect 210 101 259 123
rect 24 51 76 67
rect 110 55 126 89
rect 160 55 176 89
rect 110 17 176 55
rect 210 67 212 101
rect 246 67 259 101
rect 393 97 459 123
rect 210 51 259 67
rect 293 55 309 89
rect 343 55 359 89
rect 293 17 359 55
rect 393 63 409 97
rect 443 63 459 97
rect 593 92 659 123
rect 393 51 459 63
rect 493 55 509 89
rect 543 55 559 89
rect 593 58 609 92
rect 643 58 659 92
rect 1004 93 1071 123
rect 593 55 659 58
rect 825 55 841 89
rect 875 55 891 89
rect 1004 59 1020 93
rect 1054 59 1071 93
rect 493 17 559 55
rect 825 17 891 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 D1
port 5 nsew signal input
flabel locali s 305 289 339 323 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel locali s 857 221 891 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 765 289 799 323 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 581 289 615 323 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 489 221 523 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a2111oi_2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 2449558
string GDS_START 2441330
string path 0.000 0.000 27.600 0.000 
<< end >>
