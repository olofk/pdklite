magic
tech sky130A
magscale 1 2
timestamp 1640697977
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 189 157 1085 203
rect 1 21 1085 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 267 47 297 177
rect 351 47 381 177
rect 435 47 465 177
rect 519 47 549 177
rect 707 47 737 177
rect 791 47 821 177
rect 893 47 923 177
rect 977 47 1007 177
<< scpmoshvt >>
rect 79 413 109 497
rect 267 297 297 497
rect 351 297 381 497
rect 435 297 465 497
rect 519 297 549 497
rect 697 297 727 497
rect 781 297 811 497
rect 883 297 913 497
rect 967 297 997 497
<< ndiff >>
rect 215 161 267 177
rect 27 103 79 131
rect 27 69 35 103
rect 69 69 79 103
rect 27 47 79 69
rect 109 93 161 131
rect 109 59 119 93
rect 153 59 161 93
rect 109 47 161 59
rect 215 127 223 161
rect 257 127 267 161
rect 215 93 267 127
rect 215 59 223 93
rect 257 59 267 93
rect 215 47 267 59
rect 297 161 351 177
rect 297 127 307 161
rect 341 127 351 161
rect 297 47 351 127
rect 381 127 435 177
rect 381 93 391 127
rect 425 93 435 127
rect 381 47 435 93
rect 465 93 519 177
rect 465 59 475 93
rect 509 59 519 93
rect 465 47 519 59
rect 549 161 601 177
rect 549 127 559 161
rect 593 127 601 161
rect 549 47 601 127
rect 655 161 707 177
rect 655 127 663 161
rect 697 127 707 161
rect 655 47 707 127
rect 737 93 791 177
rect 737 59 747 93
rect 781 59 791 93
rect 737 47 791 59
rect 821 169 893 177
rect 821 135 840 169
rect 874 135 893 169
rect 821 101 893 135
rect 821 67 840 101
rect 874 67 893 101
rect 821 47 893 67
rect 923 93 977 177
rect 923 59 933 93
rect 967 59 977 93
rect 923 47 977 59
rect 1007 161 1059 177
rect 1007 127 1017 161
rect 1051 127 1059 161
rect 1007 93 1059 127
rect 1007 59 1017 93
rect 1051 59 1059 93
rect 1007 47 1059 59
<< pdiff >>
rect 27 475 79 497
rect 27 441 35 475
rect 69 441 79 475
rect 27 413 79 441
rect 109 485 161 497
rect 109 451 119 485
rect 153 451 161 485
rect 109 413 161 451
rect 215 485 267 497
rect 215 451 223 485
rect 257 451 267 485
rect 215 417 267 451
rect 215 383 223 417
rect 257 383 267 417
rect 215 349 267 383
rect 215 315 223 349
rect 257 315 267 349
rect 215 297 267 315
rect 297 485 351 497
rect 297 451 307 485
rect 341 451 351 485
rect 297 417 351 451
rect 297 383 307 417
rect 341 383 351 417
rect 297 349 351 383
rect 297 315 307 349
rect 341 315 351 349
rect 297 297 351 315
rect 381 485 435 497
rect 381 451 391 485
rect 425 451 435 485
rect 381 417 435 451
rect 381 383 391 417
rect 425 383 435 417
rect 381 297 435 383
rect 465 485 519 497
rect 465 451 475 485
rect 509 451 519 485
rect 465 417 519 451
rect 465 383 475 417
rect 509 383 519 417
rect 465 349 519 383
rect 465 315 475 349
rect 509 315 519 349
rect 465 297 519 315
rect 549 485 697 497
rect 549 451 559 485
rect 593 451 637 485
rect 671 451 697 485
rect 549 417 697 451
rect 549 383 559 417
rect 593 383 637 417
rect 671 383 697 417
rect 549 297 697 383
rect 727 485 781 497
rect 727 451 737 485
rect 771 451 781 485
rect 727 417 781 451
rect 727 383 737 417
rect 771 383 781 417
rect 727 349 781 383
rect 727 315 737 349
rect 771 315 781 349
rect 727 297 781 315
rect 811 485 883 497
rect 811 451 828 485
rect 862 451 883 485
rect 811 417 883 451
rect 811 383 828 417
rect 862 383 883 417
rect 811 297 883 383
rect 913 485 967 497
rect 913 451 923 485
rect 957 451 967 485
rect 913 417 967 451
rect 913 383 923 417
rect 957 383 967 417
rect 913 297 967 383
rect 997 485 1077 497
rect 997 451 1023 485
rect 1057 451 1077 485
rect 997 417 1077 451
rect 997 383 1023 417
rect 1057 383 1077 417
rect 997 349 1077 383
rect 997 315 1023 349
rect 1057 315 1077 349
rect 997 297 1077 315
<< ndiffc >>
rect 35 69 69 103
rect 119 59 153 93
rect 223 127 257 161
rect 223 59 257 93
rect 307 127 341 161
rect 391 93 425 127
rect 475 59 509 93
rect 559 127 593 161
rect 663 127 697 161
rect 747 59 781 93
rect 840 135 874 169
rect 840 67 874 101
rect 933 59 967 93
rect 1017 127 1051 161
rect 1017 59 1051 93
<< pdiffc >>
rect 35 441 69 475
rect 119 451 153 485
rect 223 451 257 485
rect 223 383 257 417
rect 223 315 257 349
rect 307 451 341 485
rect 307 383 341 417
rect 307 315 341 349
rect 391 451 425 485
rect 391 383 425 417
rect 475 451 509 485
rect 475 383 509 417
rect 475 315 509 349
rect 559 451 593 485
rect 637 451 671 485
rect 559 383 593 417
rect 637 383 671 417
rect 737 451 771 485
rect 737 383 771 417
rect 737 315 771 349
rect 828 451 862 485
rect 828 383 862 417
rect 923 451 957 485
rect 923 383 957 417
rect 1023 451 1057 485
rect 1023 383 1057 417
rect 1023 315 1057 349
<< poly >>
rect 79 497 109 523
rect 267 497 297 523
rect 351 497 381 523
rect 435 497 465 523
rect 519 497 549 523
rect 697 497 727 523
rect 781 497 811 523
rect 883 497 913 523
rect 967 497 997 523
rect 79 265 109 413
rect 267 265 297 297
rect 351 265 381 297
rect 22 249 109 265
rect 22 215 32 249
rect 66 215 109 249
rect 22 199 109 215
rect 210 249 381 265
rect 210 215 226 249
rect 260 215 381 249
rect 210 199 381 215
rect 79 131 109 199
rect 267 177 297 199
rect 351 177 381 199
rect 435 265 465 297
rect 519 265 549 297
rect 697 265 727 297
rect 781 265 811 297
rect 883 265 913 297
rect 967 265 997 297
rect 435 249 606 265
rect 435 215 455 249
rect 489 215 556 249
rect 590 215 606 249
rect 435 199 606 215
rect 697 249 841 265
rect 697 215 713 249
rect 747 215 787 249
rect 821 215 841 249
rect 697 199 841 215
rect 883 261 1054 265
rect 883 249 1082 261
rect 883 215 940 249
rect 974 215 1032 249
rect 1066 215 1082 249
rect 883 203 1082 215
rect 883 199 1054 203
rect 435 177 465 199
rect 519 177 549 199
rect 707 177 737 199
rect 791 177 821 199
rect 893 177 923 199
rect 977 177 1007 199
rect 79 21 109 47
rect 267 21 297 47
rect 351 21 381 47
rect 435 21 465 47
rect 519 21 549 47
rect 707 21 737 47
rect 791 21 821 47
rect 893 21 923 47
rect 977 21 1007 47
<< polycont >>
rect 32 215 66 249
rect 226 215 260 249
rect 455 215 489 249
rect 556 215 590 249
rect 713 215 747 249
rect 787 215 821 249
rect 940 215 974 249
rect 1032 215 1066 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 18 475 69 493
rect 18 441 35 475
rect 103 485 257 527
rect 103 451 119 485
rect 153 451 223 485
rect 18 417 69 441
rect 207 417 257 451
rect 18 383 134 417
rect 18 249 66 323
rect 18 215 32 249
rect 18 199 66 215
rect 100 249 134 383
rect 207 383 223 417
rect 207 349 257 383
rect 207 315 223 349
rect 207 289 257 315
rect 291 485 357 493
rect 291 451 307 485
rect 341 451 357 485
rect 291 417 357 451
rect 291 383 307 417
rect 341 383 357 417
rect 291 349 357 383
rect 391 485 425 527
rect 391 417 425 451
rect 391 367 425 383
rect 459 485 525 493
rect 459 451 475 485
rect 509 451 525 485
rect 459 417 525 451
rect 459 383 475 417
rect 509 383 525 417
rect 291 315 307 349
rect 341 333 357 349
rect 459 349 525 383
rect 559 485 687 527
rect 593 451 637 485
rect 671 451 687 485
rect 559 417 687 451
rect 593 383 637 417
rect 671 383 687 417
rect 559 367 687 383
rect 721 485 787 493
rect 721 451 737 485
rect 771 451 787 485
rect 721 417 787 451
rect 721 383 737 417
rect 771 383 787 417
rect 459 333 475 349
rect 341 315 475 333
rect 509 333 525 349
rect 721 349 787 383
rect 821 485 873 527
rect 821 451 828 485
rect 862 451 873 485
rect 821 417 873 451
rect 821 383 828 417
rect 862 383 873 417
rect 821 367 873 383
rect 907 485 973 493
rect 907 451 923 485
rect 957 451 973 485
rect 907 417 973 451
rect 907 383 923 417
rect 957 383 973 417
rect 721 333 737 349
rect 509 315 737 333
rect 771 333 787 349
rect 907 333 973 383
rect 771 315 973 333
rect 291 289 973 315
rect 1007 485 1086 527
rect 1007 451 1023 485
rect 1057 451 1086 485
rect 1007 417 1086 451
rect 1007 383 1023 417
rect 1057 383 1086 417
rect 1007 349 1086 383
rect 1007 315 1023 349
rect 1057 315 1086 349
rect 1007 299 1086 315
rect 100 215 226 249
rect 260 215 276 249
rect 100 161 134 215
rect 18 127 134 161
rect 207 161 257 181
rect 310 165 357 289
rect 402 249 620 255
rect 402 215 455 249
rect 489 215 556 249
rect 590 215 620 249
rect 672 249 890 255
rect 672 215 713 249
rect 747 215 787 249
rect 821 215 890 249
rect 924 249 1086 255
rect 924 215 940 249
rect 974 215 1032 249
rect 1066 215 1086 249
rect 207 127 223 161
rect 291 161 357 165
rect 291 127 307 161
rect 341 127 357 161
rect 391 161 609 181
rect 391 127 559 161
rect 593 127 609 161
rect 647 169 1068 181
rect 647 161 840 169
rect 647 127 663 161
rect 697 135 840 161
rect 874 161 1068 169
rect 874 143 1017 161
rect 874 135 891 143
rect 697 127 891 135
rect 18 103 69 127
rect 18 69 35 103
rect 207 93 257 127
rect 831 123 891 127
rect 1001 127 1017 143
rect 1051 127 1068 161
rect 831 101 883 123
rect 18 51 69 69
rect 103 59 119 93
rect 153 59 169 93
rect 103 17 169 59
rect 207 59 223 93
rect 257 59 425 93
rect 207 51 425 59
rect 459 59 475 93
rect 509 59 747 93
rect 781 59 797 93
rect 459 51 797 59
rect 831 67 840 101
rect 874 67 883 101
rect 831 51 883 67
rect 933 93 967 109
rect 933 17 967 59
rect 1001 93 1068 127
rect 1001 59 1017 93
rect 1051 59 1068 93
rect 1001 51 1068 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel locali s 1040 221 1074 255 0 FreeSans 250 0 0 0 D
port 4 nsew signal input
flabel locali s 948 221 982 255 0 FreeSans 250 0 0 0 D
port 4 nsew signal input
flabel locali s 856 221 890 255 0 FreeSans 250 0 0 0 C
port 3 nsew signal input
flabel locali s 764 221 798 255 0 FreeSans 250 0 0 0 C
port 3 nsew signal input
flabel locali s 672 221 706 255 0 FreeSans 250 0 0 0 C
port 3 nsew signal input
flabel locali s 586 221 620 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 494 221 528 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 402 221 436 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 310 153 344 187 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel locali s 310 221 344 255 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel locali s 310 289 344 323 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 250 0 0 0 A_N
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 250 0 0 0 A_N
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nand4b_2
rlabel metal1 s 0 -48 1104 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 1920460
string GDS_START 1910404
string path 0.000 0.000 27.600 0.000 
<< end >>
