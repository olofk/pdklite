magic
tech sky130A
magscale 1 2
timestamp 1640697850
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_0
timestamp 1640697850
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_1
timestamp 1640697850
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_2
timestamp 1640697850
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_3
timestamp 1640697850
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_4
timestamp 1640697850
transform 1 0 724 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_5
timestamp 1640697850
transform 1 0 880 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_6
timestamp 1640697850
transform 1 0 1036 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_7
timestamp 1640697850
transform 1 0 1192 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_8
timestamp 1640697850
transform 1 0 1348 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_9
timestamp 1640697850
transform 1 0 1504 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_10
timestamp 1640697850
transform 1 0 1660 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_11
timestamp 1640697850
transform 1 0 1816 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_12
timestamp 1640697850
transform 1 0 1972 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_13
timestamp 1640697850
transform 1 0 2128 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_14
timestamp 1640697850
transform 1 0 2284 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_15
timestamp 1640697850
transform 1 0 2440 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_16
timestamp 1640697850
transform 1 0 2596 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_17
timestamp 1640697850
transform 1 0 2752 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_18
timestamp 1640697850
transform 1 0 2908 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_19
timestamp 1640697850
transform 1 0 3064 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_20
timestamp 1640697850
transform 1 0 3220 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_21
timestamp 1640697850
transform 1 0 3376 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_22
timestamp 1640697850
transform 1 0 3532 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_23
timestamp 1640697850
transform 1 0 3688 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_24
timestamp 1640697850
transform 1 0 3844 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_25
timestamp 1640697850
transform 1 0 4000 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_26
timestamp 1640697850
transform 1 0 4156 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_27
timestamp 1640697850
transform 1 0 4312 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_28
timestamp 1640697850
transform 1 0 4468 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_29
timestamp 1640697850
transform 1 0 4624 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_30
timestamp 1640697850
transform 1 0 4780 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_31
timestamp 1640697850
transform 1 0 4936 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_32
timestamp 1640697850
transform 1 0 5092 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_33
timestamp 1640697850
transform 1 0 5248 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_34
timestamp 1640697850
transform 1 0 5404 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_35
timestamp 1640697850
transform 1 0 5560 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_36
timestamp 1640697850
transform 1 0 5716 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_37
timestamp 1640697850
transform 1 0 5872 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_38
timestamp 1640697850
transform 1 0 6028 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_39
timestamp 1640697850
transform 1 0 6184 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_40
timestamp 1640697850
transform 1 0 6340 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_41
timestamp 1640697850
transform 1 0 6496 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_42
timestamp 1640697850
transform 1 0 6652 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_43
timestamp 1640697850
transform 1 0 6808 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_44
timestamp 1640697850
transform 1 0 6964 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_45
timestamp 1640697850
transform 1 0 7120 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_46
timestamp 1640697850
transform 1 0 7276 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_47
timestamp 1640697850
transform 1 0 7432 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_48
timestamp 1640697850
transform 1 0 7588 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808336  sky130_fd_pr__dfl1sd__example_55959141808336_0
timestamp 1640697850
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808336  sky130_fd_pr__dfl1sd__example_55959141808336_1
timestamp 1640697850
transform 1 0 7744 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 7772 675 7772 675 0 FreeSans 300 0 0 0 S
flabel comment s 7616 675 7616 675 0 FreeSans 300 0 0 0 D
flabel comment s 7460 675 7460 675 0 FreeSans 300 0 0 0 S
flabel comment s 7304 675 7304 675 0 FreeSans 300 0 0 0 D
flabel comment s 7148 675 7148 675 0 FreeSans 300 0 0 0 S
flabel comment s 6992 675 6992 675 0 FreeSans 300 0 0 0 D
flabel comment s 6836 675 6836 675 0 FreeSans 300 0 0 0 S
flabel comment s 6680 675 6680 675 0 FreeSans 300 0 0 0 D
flabel comment s 6524 675 6524 675 0 FreeSans 300 0 0 0 S
flabel comment s 6368 675 6368 675 0 FreeSans 300 0 0 0 D
flabel comment s 6212 675 6212 675 0 FreeSans 300 0 0 0 S
flabel comment s 6056 675 6056 675 0 FreeSans 300 0 0 0 D
flabel comment s 5900 675 5900 675 0 FreeSans 300 0 0 0 S
flabel comment s 5744 675 5744 675 0 FreeSans 300 0 0 0 D
flabel comment s 5588 675 5588 675 0 FreeSans 300 0 0 0 S
flabel comment s 5432 675 5432 675 0 FreeSans 300 0 0 0 D
flabel comment s 5276 675 5276 675 0 FreeSans 300 0 0 0 S
flabel comment s 5120 675 5120 675 0 FreeSans 300 0 0 0 D
flabel comment s 4964 675 4964 675 0 FreeSans 300 0 0 0 S
flabel comment s 4808 675 4808 675 0 FreeSans 300 0 0 0 D
flabel comment s 4652 675 4652 675 0 FreeSans 300 0 0 0 S
flabel comment s 4496 675 4496 675 0 FreeSans 300 0 0 0 D
flabel comment s 4340 675 4340 675 0 FreeSans 300 0 0 0 S
flabel comment s 4184 675 4184 675 0 FreeSans 300 0 0 0 D
flabel comment s 4028 675 4028 675 0 FreeSans 300 0 0 0 S
flabel comment s 3872 675 3872 675 0 FreeSans 300 0 0 0 D
flabel comment s 3716 675 3716 675 0 FreeSans 300 0 0 0 S
flabel comment s 3560 675 3560 675 0 FreeSans 300 0 0 0 D
flabel comment s 3404 675 3404 675 0 FreeSans 300 0 0 0 S
flabel comment s 3248 675 3248 675 0 FreeSans 300 0 0 0 D
flabel comment s 3092 675 3092 675 0 FreeSans 300 0 0 0 S
flabel comment s 2936 675 2936 675 0 FreeSans 300 0 0 0 D
flabel comment s 2780 675 2780 675 0 FreeSans 300 0 0 0 S
flabel comment s 2624 675 2624 675 0 FreeSans 300 0 0 0 D
flabel comment s 2468 675 2468 675 0 FreeSans 300 0 0 0 S
flabel comment s 2312 675 2312 675 0 FreeSans 300 0 0 0 D
flabel comment s 2156 675 2156 675 0 FreeSans 300 0 0 0 S
flabel comment s 2000 675 2000 675 0 FreeSans 300 0 0 0 D
flabel comment s 1844 675 1844 675 0 FreeSans 300 0 0 0 S
flabel comment s 1688 675 1688 675 0 FreeSans 300 0 0 0 D
flabel comment s 1532 675 1532 675 0 FreeSans 300 0 0 0 S
flabel comment s 1376 675 1376 675 0 FreeSans 300 0 0 0 D
flabel comment s 1220 675 1220 675 0 FreeSans 300 0 0 0 S
flabel comment s 1064 675 1064 675 0 FreeSans 300 0 0 0 D
flabel comment s 908 675 908 675 0 FreeSans 300 0 0 0 S
flabel comment s 752 675 752 675 0 FreeSans 300 0 0 0 D
flabel comment s 596 675 596 675 0 FreeSans 300 0 0 0 S
flabel comment s 440 675 440 675 0 FreeSans 300 0 0 0 D
flabel comment s 284 675 284 675 0 FreeSans 300 0 0 0 S
flabel comment s 128 675 128 675 0 FreeSans 300 0 0 0 D
flabel comment s -28 675 -28 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 11317482
string GDS_START 11291148
<< end >>
