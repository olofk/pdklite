magic
tech sky130A
magscale 1 2
timestamp 1619729571
<< checkpaint >>
rect -1298 -1308 3230 1852
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 355 47 385 131
rect 453 47 483 131
rect 531 47 561 131
rect 627 47 657 131
rect 703 47 733 131
rect 904 47 934 119
rect 1000 47 1030 119
rect 1098 47 1128 131
rect 1244 47 1274 175
rect 1345 47 1375 119
rect 1448 47 1478 119
rect 1543 47 1573 131
rect 1731 47 1761 177
rect 1822 47 1852 177
<< scpmoshvt >>
rect 80 363 110 491
rect 164 363 194 491
rect 352 369 382 497
rect 437 369 467 497
rect 526 369 556 497
rect 610 369 640 497
rect 704 369 734 497
rect 903 413 933 497
rect 996 413 1026 497
rect 1092 413 1122 497
rect 1224 347 1254 497
rect 1319 413 1349 497
rect 1403 413 1433 497
rect 1520 413 1550 497
rect 1731 297 1761 497
rect 1822 297 1852 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 93 355 131
rect 299 59 308 93
rect 342 59 355 93
rect 299 47 355 59
rect 385 89 453 131
rect 385 55 408 89
rect 442 55 453 89
rect 385 47 453 55
rect 483 47 531 131
rect 561 89 627 131
rect 561 55 582 89
rect 616 55 627 89
rect 561 47 627 55
rect 657 47 703 131
rect 733 93 795 131
rect 1194 131 1244 175
rect 1048 119 1098 131
rect 733 59 753 93
rect 787 59 795 93
rect 733 47 795 59
rect 849 107 904 119
rect 849 73 857 107
rect 891 73 904 107
rect 849 47 904 73
rect 934 107 1000 119
rect 934 73 956 107
rect 990 73 1000 107
rect 934 47 1000 73
rect 1030 47 1098 119
rect 1128 101 1244 131
rect 1128 67 1172 101
rect 1206 67 1244 101
rect 1128 47 1244 67
rect 1274 119 1324 175
rect 1679 162 1731 177
rect 1493 119 1543 131
rect 1274 107 1345 119
rect 1274 73 1290 107
rect 1324 73 1345 107
rect 1274 47 1345 73
rect 1375 107 1448 119
rect 1375 73 1402 107
rect 1436 73 1448 107
rect 1375 47 1448 73
rect 1478 47 1543 119
rect 1573 107 1625 131
rect 1573 73 1583 107
rect 1617 73 1625 107
rect 1573 47 1625 73
rect 1679 128 1687 162
rect 1721 128 1731 162
rect 1679 94 1731 128
rect 1679 60 1687 94
rect 1721 60 1731 94
rect 1679 47 1731 60
rect 1761 123 1822 177
rect 1761 89 1775 123
rect 1809 89 1822 123
rect 1761 47 1822 89
rect 1852 164 1904 177
rect 1852 130 1862 164
rect 1896 130 1904 164
rect 1852 96 1904 130
rect 1852 62 1862 96
rect 1896 62 1904 96
rect 1852 47 1904 62
<< pdiff >>
rect 28 477 80 491
rect 28 443 36 477
rect 70 443 80 477
rect 28 409 80 443
rect 28 375 36 409
rect 70 375 80 409
rect 28 363 80 375
rect 110 461 164 491
rect 110 427 120 461
rect 154 427 164 461
rect 110 363 164 427
rect 194 477 246 491
rect 194 443 204 477
rect 238 443 246 477
rect 194 409 246 443
rect 194 375 204 409
rect 238 375 246 409
rect 194 363 246 375
rect 300 452 352 497
rect 300 418 308 452
rect 342 418 352 452
rect 300 369 352 418
rect 382 483 437 497
rect 382 449 392 483
rect 426 449 437 483
rect 382 369 437 449
rect 467 369 526 497
rect 556 483 610 497
rect 556 449 566 483
rect 600 449 610 483
rect 556 369 610 449
rect 640 369 704 497
rect 734 483 788 497
rect 734 449 746 483
rect 780 449 788 483
rect 734 369 788 449
rect 842 472 903 497
rect 842 438 850 472
rect 884 438 903 472
rect 842 413 903 438
rect 933 472 996 497
rect 933 438 948 472
rect 982 438 996 472
rect 933 413 996 438
rect 1026 413 1092 497
rect 1122 485 1224 497
rect 1122 451 1180 485
rect 1214 451 1224 485
rect 1122 417 1224 451
rect 1122 413 1180 417
rect 1137 383 1180 413
rect 1214 383 1224 417
rect 1137 347 1224 383
rect 1254 477 1319 497
rect 1254 443 1264 477
rect 1298 443 1319 477
rect 1254 413 1319 443
rect 1349 467 1403 497
rect 1349 433 1359 467
rect 1393 433 1403 467
rect 1349 413 1403 433
rect 1433 413 1520 497
rect 1550 477 1625 497
rect 1550 443 1582 477
rect 1616 443 1625 477
rect 1550 413 1625 443
rect 1679 475 1731 497
rect 1679 441 1687 475
rect 1721 441 1731 475
rect 1254 347 1304 413
rect 1679 353 1731 441
rect 1679 319 1687 353
rect 1721 319 1731 353
rect 1679 297 1731 319
rect 1761 455 1822 497
rect 1761 421 1775 455
rect 1809 421 1822 455
rect 1761 375 1822 421
rect 1761 341 1775 375
rect 1809 341 1822 375
rect 1761 297 1822 341
rect 1852 479 1904 497
rect 1852 445 1862 479
rect 1896 445 1904 479
rect 1852 411 1904 445
rect 1852 377 1862 411
rect 1896 377 1904 411
rect 1852 343 1904 377
rect 1852 309 1862 343
rect 1896 309 1904 343
rect 1852 297 1904 309
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 308 59 342 93
rect 408 55 442 89
rect 582 55 616 89
rect 753 59 787 93
rect 857 73 891 107
rect 956 73 990 107
rect 1172 67 1206 101
rect 1290 73 1324 107
rect 1402 73 1436 107
rect 1583 73 1617 107
rect 1687 128 1721 162
rect 1687 60 1721 94
rect 1775 89 1809 123
rect 1862 130 1896 164
rect 1862 62 1896 96
<< pdiffc >>
rect 36 443 70 477
rect 36 375 70 409
rect 120 427 154 461
rect 204 443 238 477
rect 204 375 238 409
rect 308 418 342 452
rect 392 449 426 483
rect 566 449 600 483
rect 746 449 780 483
rect 850 438 884 472
rect 948 438 982 472
rect 1180 451 1214 485
rect 1180 383 1214 417
rect 1264 443 1298 477
rect 1359 433 1393 467
rect 1582 443 1616 477
rect 1687 441 1721 475
rect 1687 319 1721 353
rect 1775 421 1809 455
rect 1775 341 1809 375
rect 1862 445 1896 479
rect 1862 377 1896 411
rect 1862 309 1896 343
<< poly >>
rect 80 491 110 517
rect 164 491 194 517
rect 352 497 382 523
rect 437 497 467 523
rect 526 497 556 523
rect 610 497 640 523
rect 704 497 734 523
rect 903 497 933 523
rect 996 497 1026 523
rect 1092 497 1122 523
rect 1224 497 1254 523
rect 1319 497 1349 523
rect 1403 497 1433 523
rect 1520 497 1550 523
rect 1731 497 1761 523
rect 1822 497 1852 523
rect 903 375 933 413
rect 996 381 1026 413
rect 80 348 110 363
rect 47 318 110 348
rect 47 265 77 318
rect 164 274 194 363
rect 352 331 382 369
rect 437 331 467 369
rect 526 337 556 369
rect 340 321 467 331
rect 340 287 352 321
rect 386 301 467 321
rect 514 321 568 337
rect 386 287 402 301
rect 340 277 402 287
rect 514 287 524 321
rect 558 287 568 321
rect 23 249 77 265
rect 23 215 33 249
rect 67 215 77 249
rect 119 264 194 274
rect 119 230 135 264
rect 169 230 194 264
rect 119 220 194 230
rect 23 199 77 215
rect 47 176 77 199
rect 47 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 351 163 381 277
rect 514 271 568 287
rect 610 327 640 369
rect 704 354 734 369
rect 888 365 954 375
rect 704 343 736 354
rect 610 311 664 327
rect 610 277 620 311
rect 654 277 664 311
rect 423 226 489 236
rect 423 192 439 226
rect 473 192 489 226
rect 423 182 489 192
rect 351 146 385 163
rect 355 131 385 146
rect 453 131 483 182
rect 531 131 561 271
rect 610 261 664 277
rect 706 304 736 343
rect 888 331 904 365
rect 938 331 954 365
rect 888 321 954 331
rect 996 365 1050 381
rect 996 331 1006 365
rect 1040 331 1050 365
rect 996 315 1050 331
rect 706 288 760 304
rect 706 254 716 288
rect 750 254 760 288
rect 996 279 1026 315
rect 706 238 760 254
rect 703 220 760 238
rect 904 249 1026 279
rect 603 203 657 219
rect 603 169 613 203
rect 647 169 657 203
rect 603 153 657 169
rect 627 131 657 153
rect 703 131 733 220
rect 904 119 934 249
rect 1092 213 1122 413
rect 1224 309 1254 347
rect 1319 315 1349 413
rect 1403 375 1433 413
rect 1520 381 1550 413
rect 1402 365 1468 375
rect 1402 331 1418 365
rect 1452 331 1468 365
rect 1402 321 1468 331
rect 1520 365 1598 381
rect 1520 331 1554 365
rect 1588 331 1598 365
rect 1520 315 1598 331
rect 1164 299 1254 309
rect 1164 265 1180 299
rect 1214 265 1254 299
rect 1164 255 1254 265
rect 1224 220 1254 255
rect 1306 299 1360 315
rect 1306 265 1316 299
rect 1350 279 1360 299
rect 1350 265 1478 279
rect 1306 249 1478 265
rect 976 191 1030 207
rect 976 157 986 191
rect 1020 157 1030 191
rect 1092 203 1172 213
rect 1092 183 1122 203
rect 976 141 1030 157
rect 1000 119 1030 141
rect 1098 169 1122 183
rect 1156 169 1172 203
rect 1224 190 1274 220
rect 1244 175 1274 190
rect 1345 191 1406 207
rect 1098 159 1172 169
rect 1098 131 1128 159
rect 1345 157 1362 191
rect 1396 157 1406 191
rect 1345 141 1406 157
rect 1345 119 1375 141
rect 1448 119 1478 249
rect 1543 131 1573 315
rect 1731 265 1761 297
rect 1822 265 1852 297
rect 1629 249 1761 265
rect 1629 215 1639 249
rect 1673 215 1761 249
rect 1629 199 1761 215
rect 1803 249 1867 265
rect 1803 215 1813 249
rect 1847 215 1867 249
rect 1803 199 1867 215
rect 1731 177 1761 199
rect 1822 177 1852 199
rect 79 21 109 47
rect 163 21 193 47
rect 355 21 385 47
rect 453 21 483 47
rect 531 21 561 47
rect 627 21 657 47
rect 703 21 733 47
rect 904 21 934 47
rect 1000 21 1030 47
rect 1098 21 1128 47
rect 1244 21 1274 47
rect 1345 21 1375 47
rect 1448 21 1478 47
rect 1543 21 1573 47
rect 1731 21 1761 47
rect 1822 21 1852 47
<< polycont >>
rect 352 287 386 321
rect 524 287 558 321
rect 33 215 67 249
rect 135 230 169 264
rect 620 277 654 311
rect 439 192 473 226
rect 904 331 938 365
rect 1006 331 1040 365
rect 716 254 750 288
rect 613 169 647 203
rect 1418 331 1452 365
rect 1554 331 1588 365
rect 1180 265 1214 299
rect 1316 265 1350 299
rect 986 157 1020 191
rect 1122 169 1156 203
rect 1362 157 1396 191
rect 1639 215 1673 249
rect 1813 215 1847 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 36 477 70 493
rect 36 409 70 443
rect 104 461 170 527
rect 104 427 120 461
rect 154 427 170 461
rect 204 477 246 493
rect 238 443 246 477
rect 204 409 246 443
rect 70 391 169 393
rect 70 375 128 391
rect 36 359 128 375
rect 123 357 128 359
rect 162 357 169 391
rect 19 249 89 325
rect 19 215 33 249
rect 67 215 89 249
rect 19 195 89 215
rect 123 264 169 357
rect 123 230 135 264
rect 123 194 169 230
rect 238 375 246 409
rect 123 161 162 194
rect 35 127 162 161
rect 204 187 246 375
rect 204 153 208 187
rect 242 153 246 187
rect 204 143 246 153
rect 35 119 69 127
rect 203 119 246 143
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 246 119
rect 203 69 246 85
rect 284 452 342 489
rect 284 418 308 452
rect 376 483 442 527
rect 746 483 785 527
rect 376 449 392 483
rect 426 449 442 483
rect 538 449 566 483
rect 600 449 712 483
rect 284 415 342 418
rect 284 372 644 415
rect 284 93 318 372
rect 352 321 386 337
rect 352 167 386 287
rect 423 226 458 372
rect 492 321 558 337
rect 492 287 524 321
rect 492 271 558 287
rect 610 327 644 372
rect 678 399 712 449
rect 780 449 785 483
rect 746 433 785 449
rect 836 472 884 488
rect 1180 485 1214 527
rect 836 438 850 472
rect 932 438 948 472
rect 982 438 1146 472
rect 836 413 884 438
rect 836 399 870 413
rect 678 365 870 399
rect 990 391 1078 402
rect 610 311 654 327
rect 610 277 620 311
rect 610 261 654 277
rect 706 288 798 331
rect 706 254 716 288
rect 750 254 798 288
rect 423 192 439 226
rect 473 192 492 226
rect 613 203 650 219
rect 706 211 798 254
rect 647 169 650 203
rect 836 177 870 365
rect 352 157 398 167
rect 613 157 650 169
rect 352 127 650 157
rect 374 123 650 127
rect 684 143 870 177
rect 904 365 952 381
rect 938 331 952 365
rect 990 365 1041 391
rect 990 331 1006 365
rect 1040 357 1041 365
rect 1075 357 1078 391
rect 1040 331 1078 357
rect 904 207 952 331
rect 1112 315 1146 438
rect 1180 417 1214 451
rect 1180 367 1214 383
rect 1248 477 1298 493
rect 1248 443 1264 477
rect 1558 477 1619 527
rect 1248 427 1298 443
rect 1343 433 1359 467
rect 1393 433 1520 467
rect 1112 299 1214 315
rect 1112 297 1180 299
rect 1054 265 1180 297
rect 1054 263 1214 265
rect 904 191 1020 207
rect 904 187 986 191
rect 904 156 949 187
rect 103 17 169 59
rect 284 59 308 93
rect 342 59 358 93
rect 284 52 358 59
rect 392 55 408 89
rect 442 55 461 89
rect 495 61 530 123
rect 684 89 718 143
rect 836 123 870 143
rect 926 153 949 156
rect 983 157 986 187
rect 983 153 1020 157
rect 926 141 1020 153
rect 564 55 582 89
rect 616 55 718 89
rect 752 93 792 109
rect 752 59 753 93
rect 787 59 792 93
rect 392 17 461 55
rect 752 17 792 59
rect 836 107 892 123
rect 1054 107 1088 263
rect 1180 249 1214 263
rect 1122 213 1156 219
rect 1248 213 1282 427
rect 1316 391 1354 393
rect 1316 357 1318 391
rect 1352 357 1354 391
rect 1316 299 1354 357
rect 1350 265 1354 299
rect 1316 249 1354 265
rect 1388 365 1452 381
rect 1388 331 1418 365
rect 1388 315 1452 331
rect 1122 203 1282 213
rect 1388 207 1426 315
rect 1486 281 1520 433
rect 1558 443 1582 477
rect 1616 443 1619 477
rect 1558 427 1619 443
rect 1687 475 1741 491
rect 1721 441 1741 475
rect 1687 381 1741 441
rect 1554 365 1741 381
rect 1588 353 1741 365
rect 1588 331 1687 353
rect 1554 319 1687 331
rect 1721 319 1741 353
rect 1775 455 1809 527
rect 1775 375 1809 421
rect 1775 325 1809 341
rect 1846 445 1862 479
rect 1896 445 1915 479
rect 1846 411 1915 445
rect 1846 377 1862 411
rect 1896 377 1915 411
rect 1846 343 1915 377
rect 1554 315 1741 319
rect 1156 169 1282 203
rect 1122 153 1282 169
rect 836 73 857 107
rect 891 73 892 107
rect 940 73 956 107
rect 990 73 1088 107
rect 1138 101 1212 117
rect 836 57 892 73
rect 1138 67 1172 101
rect 1206 67 1212 101
rect 1248 107 1282 153
rect 1316 191 1426 207
rect 1316 187 1362 191
rect 1316 153 1326 187
rect 1360 157 1362 187
rect 1396 157 1426 191
rect 1360 153 1426 157
rect 1316 141 1426 153
rect 1460 265 1520 281
rect 1707 265 1741 315
rect 1846 309 1862 343
rect 1896 309 1915 343
rect 1846 301 1915 309
rect 1460 249 1673 265
rect 1460 215 1639 249
rect 1460 199 1673 215
rect 1707 249 1847 265
rect 1707 215 1813 249
rect 1707 199 1847 215
rect 1460 107 1494 199
rect 1707 165 1741 199
rect 1671 162 1741 165
rect 1881 164 1915 301
rect 1671 128 1687 162
rect 1721 128 1741 162
rect 1248 73 1290 107
rect 1324 73 1340 107
rect 1386 73 1402 107
rect 1436 73 1494 107
rect 1543 107 1617 123
rect 1543 73 1583 107
rect 1138 17 1212 67
rect 1543 17 1617 73
rect 1671 94 1741 128
rect 1671 60 1687 94
rect 1721 60 1741 94
rect 1775 123 1809 139
rect 1775 17 1809 89
rect 1846 130 1862 164
rect 1896 130 1915 164
rect 1846 96 1915 130
rect 1846 62 1862 96
rect 1896 62 1915 96
rect 1846 61 1915 62
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 128 357 162 391
rect 208 153 242 187
rect 1041 357 1075 391
rect 949 153 983 187
rect 1318 357 1352 391
rect 1326 153 1360 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 116 391 174 397
rect 116 357 128 391
rect 162 388 174 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 162 360 1041 388
rect 162 357 174 360
rect 116 351 174 357
rect 1029 357 1041 360
rect 1075 388 1087 391
rect 1306 391 1364 397
rect 1306 388 1318 391
rect 1075 360 1318 388
rect 1075 357 1087 360
rect 1029 351 1087 357
rect 1306 357 1318 360
rect 1352 357 1364 391
rect 1306 351 1364 357
rect 196 187 254 193
rect 196 153 208 187
rect 242 184 254 187
rect 937 187 995 193
rect 937 184 949 187
rect 242 156 949 184
rect 242 153 254 156
rect 196 147 254 153
rect 937 153 949 156
rect 983 184 995 187
rect 1314 187 1372 193
rect 1314 184 1326 187
rect 983 156 1326 184
rect 983 153 995 156
rect 937 147 995 153
rect 1314 153 1326 156
rect 1360 153 1372 187
rect 1314 147 1372 153
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfxtp_1
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel locali s 1869 425 1903 459 0 FreeSans 200 0 0 0 Q
port 9 nsew signal output
flabel locali s 1869 357 1903 391 0 FreeSans 200 0 0 0 Q
port 9 nsew signal output
flabel locali s 1869 85 1903 119 0 FreeSans 200 0 0 0 Q
port 9 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 495 85 529 119 0 FreeSans 300 0 0 0 SCE
port 4 nsew signal input
flabel locali s 501 289 535 323 0 FreeSans 300 0 0 0 D
port 2 nsew signal input
flabel locali s 749 221 783 255 0 FreeSans 300 0 0 0 SCD
port 3 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 1344940
string GDS_START 1329734
string path 0.000 13.600 48.300 13.600 
<< end >>
