magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1326 -1253 8538 3892
<< nwell >>
rect 811 2228 831 2514
rect 224 1496 934 2228
rect 4464 1464 4504 2596
<< mvnmos >>
rect 363 1179 483 1379
rect 539 1179 659 1379
rect 715 1179 835 1379
<< mvpmos >>
rect 343 1562 463 2162
rect 519 1562 639 2162
rect 695 1562 815 2162
<< mvndiff >>
rect 310 1367 363 1379
rect 310 1333 318 1367
rect 352 1333 363 1367
rect 310 1299 363 1333
rect 310 1265 318 1299
rect 352 1265 363 1299
rect 310 1231 363 1265
rect 310 1197 318 1231
rect 352 1197 363 1231
rect 310 1179 363 1197
rect 483 1179 539 1379
rect 659 1367 715 1379
rect 659 1333 670 1367
rect 704 1333 715 1367
rect 659 1299 715 1333
rect 659 1265 670 1299
rect 704 1265 715 1299
rect 659 1231 715 1265
rect 659 1197 670 1231
rect 704 1197 715 1231
rect 659 1179 715 1197
rect 835 1367 888 1379
rect 835 1333 846 1367
rect 880 1333 888 1367
rect 835 1299 888 1333
rect 835 1265 846 1299
rect 880 1265 888 1299
rect 835 1231 888 1265
rect 835 1197 846 1231
rect 880 1197 888 1231
rect 835 1179 888 1197
<< mvpdiff >>
rect 290 2150 343 2162
rect 290 2116 298 2150
rect 332 2116 343 2150
rect 290 2082 343 2116
rect 290 2048 298 2082
rect 332 2048 343 2082
rect 290 2014 343 2048
rect 290 1980 298 2014
rect 332 1980 343 2014
rect 290 1946 343 1980
rect 290 1912 298 1946
rect 332 1912 343 1946
rect 290 1878 343 1912
rect 290 1844 298 1878
rect 332 1844 343 1878
rect 290 1810 343 1844
rect 290 1776 298 1810
rect 332 1776 343 1810
rect 290 1742 343 1776
rect 290 1708 298 1742
rect 332 1708 343 1742
rect 290 1674 343 1708
rect 290 1640 298 1674
rect 332 1640 343 1674
rect 290 1562 343 1640
rect 463 2150 519 2162
rect 463 2116 474 2150
rect 508 2116 519 2150
rect 463 2082 519 2116
rect 463 2048 474 2082
rect 508 2048 519 2082
rect 463 2014 519 2048
rect 463 1980 474 2014
rect 508 1980 519 2014
rect 463 1946 519 1980
rect 463 1912 474 1946
rect 508 1912 519 1946
rect 463 1878 519 1912
rect 463 1844 474 1878
rect 508 1844 519 1878
rect 463 1810 519 1844
rect 463 1776 474 1810
rect 508 1776 519 1810
rect 463 1742 519 1776
rect 463 1708 474 1742
rect 508 1708 519 1742
rect 463 1674 519 1708
rect 463 1640 474 1674
rect 508 1640 519 1674
rect 463 1562 519 1640
rect 639 2150 695 2162
rect 639 2116 650 2150
rect 684 2116 695 2150
rect 639 2082 695 2116
rect 639 2048 650 2082
rect 684 2048 695 2082
rect 639 2014 695 2048
rect 639 1980 650 2014
rect 684 1980 695 2014
rect 639 1946 695 1980
rect 639 1912 650 1946
rect 684 1912 695 1946
rect 639 1878 695 1912
rect 639 1844 650 1878
rect 684 1844 695 1878
rect 639 1810 695 1844
rect 639 1776 650 1810
rect 684 1776 695 1810
rect 639 1742 695 1776
rect 639 1708 650 1742
rect 684 1708 695 1742
rect 639 1674 695 1708
rect 639 1640 650 1674
rect 684 1640 695 1674
rect 639 1562 695 1640
rect 815 2150 868 2162
rect 815 2116 826 2150
rect 860 2116 868 2150
rect 815 2082 868 2116
rect 815 2048 826 2082
rect 860 2048 868 2082
rect 815 2014 868 2048
rect 815 1980 826 2014
rect 860 1980 868 2014
rect 815 1946 868 1980
rect 815 1912 826 1946
rect 860 1912 868 1946
rect 815 1878 868 1912
rect 815 1844 826 1878
rect 860 1844 868 1878
rect 815 1810 868 1844
rect 815 1776 826 1810
rect 860 1776 868 1810
rect 815 1742 868 1776
rect 815 1708 826 1742
rect 860 1708 868 1742
rect 815 1674 868 1708
rect 815 1640 826 1674
rect 860 1640 868 1674
rect 815 1562 868 1640
<< mvndiffc >>
rect 318 1333 352 1367
rect 318 1265 352 1299
rect 318 1197 352 1231
rect 670 1333 704 1367
rect 670 1265 704 1299
rect 670 1197 704 1231
rect 846 1333 880 1367
rect 846 1265 880 1299
rect 846 1197 880 1231
<< mvpdiffc >>
rect 298 2116 332 2150
rect 298 2048 332 2082
rect 298 1980 332 2014
rect 298 1912 332 1946
rect 298 1844 332 1878
rect 298 1776 332 1810
rect 298 1708 332 1742
rect 298 1640 332 1674
rect 474 2116 508 2150
rect 474 2048 508 2082
rect 474 1980 508 2014
rect 474 1912 508 1946
rect 474 1844 508 1878
rect 474 1776 508 1810
rect 474 1708 508 1742
rect 474 1640 508 1674
rect 650 2116 684 2150
rect 650 2048 684 2082
rect 650 1980 684 2014
rect 650 1912 684 1946
rect 650 1844 684 1878
rect 650 1776 684 1810
rect 650 1708 684 1742
rect 650 1640 684 1674
rect 826 2116 860 2150
rect 826 2048 860 2082
rect 826 1980 860 2014
rect 826 1912 860 1946
rect 826 1844 860 1878
rect 826 1776 860 1810
rect 826 1708 860 1742
rect 826 1640 860 1674
<< poly >>
rect 343 2162 463 2188
rect 519 2162 639 2188
rect 695 2162 815 2188
rect 343 1536 463 1562
rect 519 1536 639 1562
rect 695 1536 815 1562
rect 322 1472 463 1536
rect 322 1438 338 1472
rect 372 1438 406 1472
rect 440 1438 463 1472
rect 322 1405 463 1438
rect 526 1475 639 1536
rect 526 1455 660 1475
rect 526 1421 542 1455
rect 576 1421 610 1455
rect 644 1421 660 1455
rect 526 1405 660 1421
rect 704 1472 838 1536
rect 704 1438 720 1472
rect 754 1438 788 1472
rect 822 1438 838 1472
rect 704 1405 838 1438
rect 363 1379 483 1405
rect 539 1379 659 1405
rect 715 1379 835 1405
rect 5059 1386 5113 1462
rect 363 1153 483 1179
rect 539 1153 659 1179
rect 715 1153 835 1179
rect 4857 1012 5313 1034
rect 4857 978 4893 1012
rect 4927 978 4961 1012
rect 4995 978 5029 1012
rect 5063 978 5097 1012
rect 5131 978 5165 1012
rect 5199 978 5233 1012
rect 5267 978 5313 1012
rect 4857 958 5313 978
<< polycont >>
rect 338 1438 372 1472
rect 406 1438 440 1472
rect 542 1421 576 1455
rect 610 1421 644 1455
rect 720 1438 754 1472
rect 788 1438 822 1472
rect 4893 978 4927 1012
rect 4961 978 4995 1012
rect 5029 978 5063 1012
rect 5097 978 5131 1012
rect 5165 978 5199 1012
rect 5233 978 5267 1012
<< locali >>
rect 298 2150 332 2166
rect 298 2082 332 2116
rect 298 2014 332 2048
rect 298 1946 332 1980
rect 298 1878 332 1912
rect 298 1810 332 1844
rect 298 1760 332 1776
rect 298 1688 332 1708
rect 298 1616 332 1640
rect 474 2150 508 2166
rect 650 2150 684 2166
rect 474 2082 508 2116
rect 474 2014 508 2048
rect 474 1946 508 1980
rect 474 1878 508 1912
rect 474 1810 508 1844
rect 474 1742 508 1776
rect 474 1674 508 1708
rect 368 1502 406 1536
rect 334 1472 440 1502
rect 334 1438 338 1472
rect 372 1438 406 1472
rect 334 1422 440 1438
rect 474 1386 508 1640
rect 542 2100 564 2134
rect 598 2100 616 2134
rect 542 2062 616 2100
rect 542 2028 564 2062
rect 598 2028 616 2062
rect 542 1471 616 2028
rect 650 2082 684 2116
rect 650 2014 684 2048
rect 650 1946 684 1980
rect 650 1878 684 1912
rect 650 1810 684 1844
rect 650 1760 684 1776
rect 650 1688 684 1708
rect 650 1616 684 1640
rect 826 2150 890 2166
rect 860 2116 890 2150
rect 826 2082 890 2116
rect 860 2048 890 2082
rect 826 2014 890 2048
rect 860 1954 890 2014
rect 1121 1954 1159 1988
rect 826 1946 890 1954
rect 860 1882 890 1946
rect 826 1878 890 1882
rect 860 1844 890 1878
rect 826 1810 890 1844
rect 860 1776 890 1810
rect 826 1742 890 1776
rect 860 1708 890 1742
rect 826 1674 890 1708
rect 860 1640 890 1674
rect 826 1624 890 1640
rect 720 1472 822 1488
rect 542 1455 644 1471
rect 576 1421 610 1455
rect 754 1438 788 1472
rect 720 1422 822 1438
rect 542 1405 644 1421
rect 318 1367 474 1383
rect 352 1352 474 1367
rect 738 1386 812 1422
rect 352 1333 508 1352
rect 318 1314 508 1333
rect 318 1299 474 1314
rect 352 1280 474 1299
rect 670 1367 704 1383
rect 670 1299 704 1333
rect 318 1231 352 1265
rect 318 1181 352 1197
rect 738 1352 750 1386
rect 784 1352 812 1386
rect 856 1383 890 1624
rect 738 1314 812 1352
rect 738 1280 750 1314
rect 784 1280 812 1314
rect 846 1367 890 1383
rect 880 1333 890 1367
rect 846 1299 890 1333
rect 670 1234 704 1265
rect 670 1162 704 1197
rect 880 1265 890 1299
rect 846 1231 890 1265
rect 880 1197 890 1231
rect 846 1181 890 1197
rect 4869 1432 5034 1433
rect 5059 1432 5113 1442
rect 4869 1398 4895 1432
rect 4929 1398 4967 1432
rect 5001 1398 5039 1432
rect 5073 1398 5111 1432
rect 5145 1398 5183 1432
rect 5217 1398 5255 1432
rect 5289 1398 5315 1408
rect 4869 1342 5034 1398
rect 4869 1308 4901 1342
rect 4935 1308 4973 1342
rect 5007 1308 5034 1342
rect 670 1090 704 1128
rect 4869 1012 5034 1308
rect 5136 1342 5315 1398
rect 5136 1308 5167 1342
rect 5201 1308 5239 1342
rect 5273 1308 5315 1342
rect 6311 1357 6417 1408
rect 6345 1323 6383 1357
rect 6567 1357 6673 1408
rect 6601 1323 6639 1357
rect 5136 1012 5315 1308
rect 4869 978 4893 1012
rect 4927 978 4961 1012
rect 4995 978 5029 1012
rect 5063 978 5097 1012
rect 5131 978 5165 1012
rect 5199 978 5233 1012
rect 5267 978 5315 1012
rect 4869 924 5034 978
rect 4869 890 4895 924
rect 4929 890 4967 924
rect 5001 890 5034 924
rect 4869 875 5034 890
rect 5136 924 5315 978
rect 5136 890 5169 924
rect 5203 890 5241 924
rect 5275 890 5315 924
rect 5136 875 5315 890
rect 6311 527 6349 561
rect 6567 527 6605 561
rect 3184 305 3222 339
<< viali >>
rect 298 1742 332 1760
rect 298 1726 332 1742
rect 298 1674 332 1688
rect 298 1654 332 1674
rect 298 1582 332 1616
rect 334 1502 368 1536
rect 406 1502 440 1536
rect 564 2100 598 2134
rect 564 2028 598 2062
rect 650 1742 684 1760
rect 650 1726 684 1742
rect 650 1674 684 1688
rect 650 1654 684 1674
rect 826 1980 860 1988
rect 826 1954 860 1980
rect 1087 1954 1121 1988
rect 1159 1954 1193 1988
rect 826 1912 860 1916
rect 826 1882 860 1912
rect 650 1582 684 1616
rect 474 1352 508 1386
rect 474 1280 508 1314
rect 750 1352 784 1386
rect 750 1280 784 1314
rect 670 1231 704 1234
rect 670 1200 704 1231
rect 4895 1398 4929 1432
rect 4967 1398 5001 1432
rect 5039 1398 5073 1432
rect 5111 1398 5145 1432
rect 5183 1398 5217 1432
rect 5255 1398 5289 1432
rect 4901 1308 4935 1342
rect 4973 1308 5007 1342
rect 670 1128 704 1162
rect 670 1056 704 1090
rect 5167 1308 5201 1342
rect 5239 1308 5273 1342
rect 6311 1323 6345 1357
rect 6383 1323 6417 1357
rect 6567 1323 6601 1357
rect 6639 1323 6673 1357
rect 4895 890 4929 924
rect 4967 890 5001 924
rect 5169 890 5203 924
rect 5241 890 5275 924
rect 6277 527 6311 561
rect 6349 527 6383 561
rect 6533 527 6567 561
rect 6605 527 6639 561
rect 3150 305 3184 339
rect 3222 305 3256 339
<< metal1 >>
rect -66 2284 7072 2430
rect 4464 2250 6774 2256
rect 4464 2228 4715 2250
tri 4690 2204 4714 2228 ne
rect 4714 2204 4715 2228
tri 4714 2203 4715 2204 ne
rect 4464 2180 4562 2200
tri 4562 2180 4582 2200 sw
rect 4767 2228 6774 2250
rect 4767 2204 4768 2228
tri 4768 2204 4792 2228 nw
tri 6743 2204 6767 2228 ne
rect 6767 2204 6774 2228
rect 6826 2204 6838 2256
rect 6890 2228 7072 2256
rect 6890 2204 6897 2228
tri 6897 2204 6921 2228 nw
tri 4767 2203 4768 2204 nw
rect 4715 2186 4767 2198
rect 4464 2172 4582 2180
tri 4550 2140 4582 2172 ne
tri 4582 2140 4622 2180 sw
rect 552 2134 610 2140
rect 552 2100 564 2134
rect 598 2100 610 2134
tri 4582 2105 4617 2140 ne
rect 4617 2124 4622 2140
tri 4622 2124 4638 2140 sw
rect 4715 2128 4767 2134
rect 4617 2105 4638 2124
tri 527 2068 552 2093 se
rect 552 2068 610 2100
tri 610 2068 635 2093 sw
tri 1295 2068 1320 2093 se
rect 1320 2068 1366 2105
tri 4617 2100 4622 2105 ne
rect 4622 2100 4638 2105
tri 4638 2100 4662 2124 sw
tri 5382 2100 5406 2124 se
rect 5406 2100 5412 2124
tri 4622 2072 4650 2100 ne
rect 4650 2072 5412 2100
rect 5464 2072 5476 2124
rect 5528 2100 5534 2124
tri 5534 2100 5558 2124 sw
tri 6027 2100 6051 2124 se
rect 6051 2100 6057 2124
rect 5528 2072 6057 2100
rect 6109 2072 6121 2124
rect 6173 2100 6179 2124
tri 6179 2100 6203 2124 sw
rect 6173 2072 7072 2100
rect 0 2062 1366 2068
rect 0 2028 564 2062
rect 598 2028 1366 2062
rect 0 2022 1366 2028
rect 439 1942 518 1994
rect 570 1988 1205 1994
rect 570 1954 826 1988
rect 860 1954 1087 1988
rect 1121 1954 1159 1988
rect 1193 1954 1205 1988
rect 570 1948 1205 1954
rect 570 1942 878 1948
rect 439 1930 878 1942
rect 439 1878 518 1930
rect 570 1916 878 1930
tri 878 1923 903 1948 nw
rect 570 1882 826 1916
rect 860 1882 878 1916
rect 570 1878 878 1882
rect 439 1876 878 1878
rect 4464 1800 4560 1846
rect 5700 1800 5740 1846
rect 5836 1800 5877 1846
rect 7016 1800 7072 1846
rect -66 1760 7072 1772
rect -66 1726 298 1760
rect 332 1726 650 1760
rect 684 1726 7072 1760
rect -66 1688 7072 1726
rect -66 1654 298 1688
rect 332 1654 650 1688
rect 684 1654 7072 1688
rect -66 1616 7072 1654
rect -66 1582 298 1616
rect 332 1582 650 1616
rect 684 1606 7072 1616
rect 684 1582 1445 1606
rect -66 1570 1445 1582
tri 1445 1570 1481 1606 nw
tri 1595 1570 1631 1606 ne
rect 1631 1570 7072 1606
rect 318 1536 452 1542
rect 318 1502 334 1536
rect 368 1502 406 1536
rect 440 1502 452 1536
rect 318 1496 452 1502
tri 4468 1468 4493 1493 se
rect 4493 1468 4654 1519
rect 4656 1518 4692 1519
rect 4655 1468 4693 1518
rect 4450 1467 4654 1468
rect 4656 1467 4692 1468
rect 4694 1467 5301 1519
rect 4450 1461 4607 1467
rect 4450 1416 4555 1461
tri 4468 1402 4482 1416 ne
rect 4482 1409 4555 1416
tri 4607 1442 4632 1467 nw
tri 4858 1442 4883 1467 ne
rect 4482 1402 4607 1409
rect 4883 1432 5301 1467
rect 461 1398 1157 1402
tri 1157 1398 1161 1402 sw
tri 4482 1398 4486 1402 ne
rect 4486 1398 4607 1402
rect 461 1391 1161 1398
tri 1161 1391 1168 1398 sw
tri 4486 1391 4493 1398 ne
rect 4493 1397 4607 1398
rect 4493 1391 4555 1397
rect 461 1386 1168 1391
rect 461 1352 474 1386
rect 508 1352 750 1386
rect 784 1377 1168 1386
tri 1168 1377 1182 1391 sw
tri 4529 1377 4543 1391 ne
rect 4543 1377 4555 1391
rect 784 1357 1182 1377
tri 1182 1357 1202 1377 sw
tri 4543 1365 4555 1377 ne
rect 784 1352 1202 1357
rect 461 1349 1202 1352
tri 1202 1349 1210 1357 sw
rect 461 1333 1338 1349
rect 4555 1339 4607 1345
rect 4635 1398 4687 1402
tri 4687 1398 4691 1402 sw
tri 4879 1398 4883 1402 se
rect 4883 1398 4895 1432
rect 4929 1398 4967 1432
rect 5001 1398 5039 1432
rect 5073 1398 5111 1432
rect 5145 1398 5183 1432
rect 5217 1398 5255 1432
rect 5289 1398 5301 1432
rect 4635 1396 4691 1398
rect 4687 1391 4691 1396
tri 4691 1391 4698 1398 sw
tri 4872 1391 4879 1398 se
rect 4879 1391 5301 1398
rect 4687 1377 4698 1391
tri 4698 1377 4712 1391 sw
tri 4858 1377 4872 1391 se
rect 4872 1377 5301 1391
rect 4687 1344 4739 1377
rect 461 1314 1216 1333
rect 461 1280 474 1314
rect 508 1280 750 1314
rect 784 1281 1216 1314
rect 1268 1281 1280 1333
rect 1332 1281 1338 1333
rect 784 1280 1338 1281
rect 461 1274 1338 1280
rect 4635 1332 4739 1344
rect 4687 1325 4739 1332
rect 4740 1326 4741 1376
rect 4777 1326 4778 1376
rect 4779 1342 5301 1377
rect 5786 1475 6685 1481
rect 5838 1429 6685 1475
rect 5786 1411 5838 1423
tri 5838 1404 5863 1429 nw
tri 6274 1404 6299 1429 ne
rect 6299 1404 6429 1429
tri 6429 1404 6454 1429 nw
tri 6530 1404 6555 1429 ne
rect 6555 1404 6685 1429
rect 6300 1402 6428 1403
rect 6556 1402 6684 1403
rect 5786 1353 5838 1359
rect 6300 1365 6428 1366
rect 6299 1357 6429 1364
rect 4779 1325 4901 1342
rect 4687 1308 4695 1325
tri 4695 1308 4712 1325 nw
tri 4858 1308 4875 1325 ne
rect 4875 1308 4901 1325
rect 4935 1308 4973 1342
rect 5007 1308 5167 1342
rect 5201 1308 5239 1342
rect 5273 1308 5301 1342
tri 4687 1300 4695 1308 nw
tri 4875 1300 4883 1308 ne
rect 4635 1274 4687 1280
rect 4883 1274 5301 1308
rect 6299 1323 6311 1357
rect 6345 1323 6383 1357
rect 6417 1323 6429 1357
rect 6299 1311 6429 1323
rect 6300 1309 6428 1310
rect 6299 1273 6429 1309
rect 6300 1272 6428 1273
rect 6556 1365 6684 1366
rect 6555 1357 6685 1364
rect 6555 1323 6567 1357
rect 6601 1323 6639 1357
rect 6673 1323 6685 1357
rect 6555 1311 6685 1323
rect 6556 1309 6684 1310
rect 6555 1273 6685 1309
rect 6556 1272 6684 1273
tri 6274 1246 6299 1271 se
rect 6299 1246 6429 1271
tri 6429 1246 6454 1271 sw
tri 6530 1246 6555 1271 se
rect 6555 1246 6685 1271
tri 6685 1246 6710 1271 sw
rect 594 1234 7006 1246
rect 594 1200 670 1234
rect 704 1200 7006 1234
rect 594 1162 7006 1200
rect 594 1128 670 1162
rect 704 1128 7006 1162
rect 594 1090 7006 1128
rect 594 1056 670 1090
rect 704 1056 7006 1090
rect 594 1044 7006 1056
rect 7036 1044 7072 1246
rect 4889 924 5007 936
rect 512 866 518 918
rect 570 866 1000 918
rect 1052 866 1058 918
rect 4889 890 4895 924
rect 4929 890 4967 924
rect 5001 890 5007 924
rect 4889 878 5007 890
rect 5163 924 5281 936
rect 5163 890 5169 924
rect 5203 890 5241 924
rect 5275 890 5281 924
rect 5163 878 5281 890
rect 512 854 1058 866
rect 512 802 518 854
rect 570 802 1000 854
rect 1052 802 1058 854
rect 578 632 7072 762
tri 6240 607 6265 632 ne
rect 6265 607 6395 632
tri 6395 607 6420 632 nw
rect 6266 605 6394 606
rect 5786 598 5838 604
tri 5780 579 5786 585 se
rect 994 527 1000 579
rect 1052 527 1064 579
rect 1116 573 1122 579
tri 1122 573 1128 579 sw
tri 5774 573 5780 579 se
rect 5780 573 5786 579
rect 1116 567 4017 573
tri 4017 567 4023 573 sw
tri 5768 567 5774 573 se
rect 5774 567 5786 573
rect 1116 561 4023 567
tri 4023 561 4029 567 sw
tri 5762 561 5768 567 se
rect 5768 561 5786 567
rect 1116 560 4029 561
tri 4029 560 4030 561 sw
tri 5761 560 5762 561 se
rect 5762 560 5786 561
rect 1116 557 4030 560
tri 4030 557 4033 560 sw
rect 1116 527 4033 557
tri 4033 527 4063 557 sw
rect 4635 554 5721 560
tri 3997 499 4025 527 ne
rect 4025 508 4063 527
tri 4063 508 4082 527 sw
tri 4627 508 4635 516 se
rect 4025 499 4082 508
rect 1210 493 1262 499
tri 4025 491 4033 499 ne
rect 4033 491 4082 499
tri 4082 491 4099 508 sw
tri 4610 491 4627 508 se
rect 4627 502 4635 508
rect 4687 508 5721 554
rect 5722 509 5723 559
rect 5759 509 5760 559
rect 5761 546 5786 560
rect 6266 568 6394 569
rect 6265 561 6395 567
rect 5761 534 5838 546
rect 5761 508 5786 534
rect 4687 502 4695 508
rect 4627 491 4695 502
tri 4695 491 4712 508 nw
tri 5761 491 5778 508 ne
rect 5778 491 5786 508
tri 4033 484 4040 491 ne
rect 4040 490 4688 491
rect 4040 484 4635 490
tri 4040 483 4041 484 ne
rect 4041 483 4635 484
tri 4041 475 4049 483 ne
rect 4049 475 4635 483
tri 1262 450 1287 475 sw
tri 4049 459 4065 475 ne
rect 4065 459 4635 475
tri 4065 450 4074 459 ne
rect 4074 450 4635 459
rect 1262 441 1287 450
rect 1210 429 1287 441
rect 1262 417 1287 429
tri 1287 417 1320 450 sw
tri 4074 445 4079 450 ne
rect 4079 445 4635 450
tri 4622 432 4635 445 ne
rect 4687 484 4688 490
tri 4688 484 4695 491 nw
tri 5778 484 5785 491 ne
rect 5785 484 5786 491
tri 4687 483 4688 484 nw
tri 5785 483 5786 484 ne
rect 4635 432 4687 438
tri 5838 527 5860 549 sw
rect 6265 527 6277 561
rect 6311 527 6349 561
rect 6383 527 6395 561
rect 5838 524 5860 527
tri 5860 524 5863 527 sw
rect 5838 508 5987 524
tri 5987 508 6003 524 sw
rect 6265 515 6395 527
rect 6266 513 6394 514
rect 5838 484 6003 508
tri 6003 484 6027 508 sw
rect 5838 482 5854 484
rect 5786 475 5854 482
tri 5854 475 5863 484 nw
tri 5969 475 5978 484 ne
rect 5978 475 6027 484
tri 6027 475 6036 484 sw
rect 6265 477 6395 513
rect 6266 476 6394 477
rect 6521 561 6653 567
rect 6521 527 6533 561
rect 6567 527 6605 561
rect 6639 527 6653 561
rect 5786 459 5838 475
tri 5838 459 5854 475 nw
tri 5978 459 5994 475 ne
rect 5994 459 6036 475
tri 6036 459 6052 475 sw
tri 6249 459 6265 475 se
rect 6265 459 6395 475
tri 6395 459 6411 475 sw
tri 6505 459 6521 475 se
rect 6521 459 6653 527
tri 5994 458 5995 459 ne
rect 5995 458 6052 459
rect 5787 457 5837 458
tri 5995 457 5996 458 ne
rect 5996 457 6052 458
rect 5786 421 5838 457
tri 5996 450 6003 457 ne
rect 6003 450 6052 457
tri 6052 450 6061 459 sw
tri 6240 450 6249 459 se
rect 6249 450 6411 459
tri 6411 450 6420 459 sw
tri 6496 450 6505 459 se
rect 6505 450 6653 459
tri 6003 421 6032 450 ne
rect 6032 421 6653 450
rect 5787 420 5837 421
tri 6032 420 6033 421 ne
rect 6033 420 6653 421
tri 6033 419 6034 420 ne
rect 6034 419 6653 420
rect 1262 377 3268 417
rect 1210 371 3268 377
tri 3113 346 3138 371 ne
rect 3138 339 3268 371
rect 3138 305 3150 339
rect 3184 305 3222 339
rect 3256 305 3268 339
tri 5761 311 5786 336 se
rect 5786 311 5838 419
tri 6034 417 6036 419 ne
rect 6036 417 6653 419
tri 6036 409 6044 417 ne
rect 6044 409 6653 417
rect 3138 299 3268 305
rect 4555 259 4561 311
rect 4613 259 4625 311
rect 4677 259 5838 311
<< rmetal1 >>
rect 4654 1518 4656 1519
rect 4692 1518 4694 1519
rect 4654 1468 4655 1518
rect 4693 1468 4694 1518
rect 4654 1467 4656 1468
rect 4692 1467 4694 1468
rect 4739 1376 4741 1377
rect 4739 1326 4740 1376
rect 4739 1325 4741 1326
rect 4777 1376 4779 1377
rect 4778 1326 4779 1376
rect 6299 1403 6429 1404
rect 6299 1402 6300 1403
rect 6428 1402 6429 1403
rect 6555 1403 6685 1404
rect 6555 1402 6556 1403
rect 6684 1402 6685 1403
rect 6299 1365 6300 1366
rect 6428 1365 6429 1366
rect 6299 1364 6429 1365
rect 4777 1325 4779 1326
rect 6299 1310 6429 1311
rect 6299 1309 6300 1310
rect 6428 1309 6429 1310
rect 6299 1272 6300 1273
rect 6428 1272 6429 1273
rect 6299 1271 6429 1272
rect 6555 1365 6556 1366
rect 6684 1365 6685 1366
rect 6555 1364 6685 1365
rect 6555 1310 6685 1311
rect 6555 1309 6556 1310
rect 6684 1309 6685 1310
rect 6555 1272 6556 1273
rect 6684 1272 6685 1273
rect 6555 1271 6685 1272
rect 6265 606 6395 607
rect 6265 605 6266 606
rect 6394 605 6395 606
rect 5721 559 5723 560
rect 5721 509 5722 559
rect 5721 508 5723 509
rect 5759 559 5761 560
rect 5760 509 5761 559
rect 6265 568 6266 569
rect 6394 568 6395 569
rect 6265 567 6395 568
rect 5759 508 5761 509
rect 6265 514 6395 515
rect 6265 513 6266 514
rect 6394 513 6395 514
rect 6265 476 6266 477
rect 6394 476 6395 477
rect 6265 475 6395 476
rect 5786 458 5838 459
rect 5786 457 5787 458
rect 5837 457 5838 458
rect 5786 420 5787 421
rect 5837 420 5838 421
rect 5786 419 5838 420
<< via1 >>
rect 4715 2198 4767 2250
rect 6774 2204 6826 2256
rect 6838 2204 6890 2256
rect 4715 2134 4767 2186
rect 5412 2072 5464 2124
rect 5476 2072 5528 2124
rect 6057 2072 6109 2124
rect 6121 2072 6173 2124
rect 518 1942 570 1994
rect 518 1878 570 1930
rect 4555 1409 4607 1461
rect 4555 1345 4607 1397
rect 4635 1344 4687 1396
rect 1216 1281 1268 1333
rect 1280 1281 1332 1333
rect 4635 1280 4687 1332
rect 5786 1423 5838 1475
rect 5786 1359 5838 1411
rect 518 866 570 918
rect 1000 866 1052 918
rect 518 802 570 854
rect 1000 802 1052 854
rect 1000 527 1052 579
rect 1064 527 1116 579
rect 1210 441 1262 493
rect 4635 502 4687 554
rect 5786 546 5838 598
rect 1210 377 1262 429
rect 4635 438 4687 490
rect 5786 482 5838 534
rect 4561 259 4613 311
rect 4625 259 4677 311
<< metal2 >>
tri 6804 2292 6809 2297 se
tri 6768 2256 6804 2292 se
rect 6804 2256 6809 2292
tri 6860 2256 6896 2292 sw
rect 4715 2250 4767 2256
rect 4715 2186 4767 2198
rect 6768 2204 6774 2256
rect 6826 2204 6838 2256
rect 6890 2204 6896 2256
tri 6768 2168 6804 2204 ne
rect 6804 2168 6809 2204
tri 6860 2168 6896 2204 nw
tri 6804 2164 6808 2168 ne
rect 6808 2164 6809 2168
tri 6139 2163 6140 2164 sw
tri 6808 2163 6809 2164 ne
tri 6082 2155 6087 2160 se
rect 4715 2128 4767 2134
tri 5410 2128 5437 2155 se
tri 5406 2124 5410 2128 se
rect 5410 2124 5437 2128
tri 5489 2124 5520 2155 sw
tri 6051 2124 6082 2155 se
rect 6082 2124 6087 2155
rect 6139 2124 6140 2163
tri 6140 2124 6179 2163 sw
rect 5406 2072 5412 2124
rect 5464 2072 5476 2124
rect 5528 2072 5534 2124
rect 6051 2072 6057 2124
rect 6109 2072 6121 2124
rect 6173 2072 6179 2124
tri 5406 2041 5437 2072 ne
tri 5489 2041 5520 2072 nw
tri 6052 2041 6083 2072 ne
rect 6083 2041 6087 2072
tri 6083 2037 6087 2041 ne
rect 6139 2037 6144 2072
tri 6144 2037 6179 2072 nw
tri 6139 2032 6144 2037 nw
rect 512 1942 518 1994
rect 570 1942 576 1994
rect 512 1930 576 1942
rect 512 1878 518 1930
rect 570 1878 576 1930
rect 512 918 576 1878
rect 5786 1475 5838 1481
rect 4555 1461 4607 1467
rect 4555 1397 4607 1409
rect 5786 1411 5838 1423
rect 1210 1281 1216 1333
rect 1268 1281 1280 1333
rect 1332 1281 1338 1333
rect 1210 1280 1337 1281
tri 1337 1280 1338 1281 nw
rect 512 866 518 918
rect 570 866 576 918
rect 512 854 576 866
rect 512 802 518 854
rect 570 802 576 854
rect 994 866 1000 918
rect 1052 866 1058 918
rect 994 854 1058 866
rect 994 802 1000 854
rect 1052 802 1058 854
rect 994 598 1058 802
tri 1058 598 1079 619 sw
rect 994 579 1079 598
tri 1079 579 1098 598 sw
rect 994 527 1000 579
rect 1052 527 1064 579
rect 1116 527 1122 579
rect 1210 493 1262 1280
tri 1262 1205 1337 1280 nw
rect 1210 429 1262 441
rect 1210 371 1262 377
rect 4555 311 4607 1345
rect 4635 1396 4687 1402
rect 4635 1332 4687 1344
rect 4635 554 4687 1280
rect 4635 490 4687 502
rect 5786 598 5838 1359
rect 5786 534 5838 546
rect 5786 476 5838 482
rect 4635 432 4687 438
tri 4607 311 4651 355 sw
rect 4555 259 4561 311
rect 4613 259 4625 311
rect 4677 259 4683 311
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1619729480
transform 1 0 526 0 -1 1471
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1619729480
transform 1 0 322 0 -1 1488
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_2
timestamp 1619729480
transform 1 0 704 0 1 1422
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808272  sky130_fd_pr__via_pol1__example_55959141808272_0
timestamp 1619729480
transform 0 1 4877 1 0 962
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808271  sky130_fd_pr__via_m1m2__example_55959141808271_0
timestamp 1619729480
transform 1 0 512 0 -1 1994
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808271  sky130_fd_pr__via_m1m2__example_55959141808271_1
timestamp 1619729480
transform 1 0 512 0 -1 918
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808271  sky130_fd_pr__via_m1m2__example_55959141808271_2
timestamp 1619729480
transform 1 0 994 0 -1 918
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1619729480
transform 0 1 1210 -1 0 499
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1619729480
transform 0 1 5786 -1 0 1481
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1619729480
transform 1 0 4555 0 -1 311
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1619729480
transform 0 -1 4607 -1 0 1467
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_4
timestamp 1619729480
transform 0 -1 5838 -1 0 604
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_5
timestamp 1619729480
transform 0 -1 4687 -1 0 1402
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_6
timestamp 1619729480
transform 0 -1 4687 1 0 432
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_7
timestamp 1619729480
transform 1 0 6768 0 -1 2256
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_8
timestamp 1619729480
transform 1 0 5406 0 -1 2124
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_9
timestamp 1619729480
transform 1 0 6051 0 -1 2124
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_10
timestamp 1619729480
transform 0 1 4715 1 0 2128
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1619729480
transform 0 -1 684 -1 0 1760
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1619729480
transform 0 -1 704 -1 0 1234
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_2
timestamp 1619729480
transform 0 -1 332 -1 0 1760
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808270  sky130_fd_pr__via_l1m1__example_55959141808270_0
timestamp 1619729480
transform 1 0 4895 0 1 1398
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_0
timestamp 1619729480
transform -1 0 598 0 1 2028
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_1
timestamp 1619729480
transform -1 0 860 0 1 1882
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_2
timestamp 1619729480
transform -1 0 508 0 1 1280
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_3
timestamp 1619729480
transform -1 0 784 0 1 1280
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_4
timestamp 1619729480
transform 0 1 4895 1 0 890
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_5
timestamp 1619729480
transform 0 1 5169 1 0 890
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_6
timestamp 1619729480
transform 0 1 4901 1 0 1308
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_7
timestamp 1619729480
transform 0 1 5167 1 0 1308
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1619729480
transform -1 0 440 0 -1 1536
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1619729480
transform -1 0 6417 0 1 1323
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1619729480
transform 1 0 6277 0 1 527
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1619729480
transform -1 0 6673 0 1 1323
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1619729480
transform 1 0 6533 0 1 527
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1619729480
transform -1 0 1193 0 1 1954
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1619729480
transform -1 0 3256 0 1 305
box 0 0 1 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808101  sky130_fd_pr__model__pfet_highvoltage__example_55959141808101_0
timestamp 1619729480
transform 1 0 695 0 -1 2162
box -28 0 148 267
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808142  sky130_fd_pr__model__pfet_highvoltage__example_55959141808142_0
timestamp 1619729480
transform 1 0 343 0 -1 2162
box -28 0 324 267
use sky130_fd_pr__model__nfet_highvoltage__example_5595914180899  sky130_fd_pr__model__nfet_highvoltage__example_5595914180899_0
timestamp 1619729480
transform 1 0 715 0 -1 1379
box -28 0 148 97
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808144  sky130_fd_pr__model__nfet_highvoltage__example_55959141808144_0
timestamp 1619729480
transform 1 0 363 0 -1 1379
box -28 0 145 100
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808144  sky130_fd_pr__model__nfet_highvoltage__example_55959141808144_1
timestamp 1619729480
transform -1 0 659 0 -1 1379
box -28 0 145 100
use sky130_fd_io__tk_em1o_cdns_55959141808289  sky130_fd_io__tk_em1o_cdns_55959141808289_0
timestamp 1619729480
transform 0 -1 6685 1 0 1312
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_55959141808289  sky130_fd_io__tk_em1o_cdns_55959141808289_1
timestamp 1619729480
transform 0 -1 6395 1 0 515
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_55959141808289  sky130_fd_io__tk_em1o_cdns_55959141808289_2
timestamp 1619729480
transform 0 -1 6429 1 0 1312
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_0
timestamp 1619729480
transform 1 0 4687 0 1 1325
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_1
timestamp 1619729480
transform 1 0 5669 0 1 508
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_55959141808288  sky130_fd_io__tk_em1s_cdns_55959141808288_0
timestamp 1619729480
transform 0 -1 6685 1 0 1219
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_55959141808288  sky130_fd_io__tk_em1s_cdns_55959141808288_1
timestamp 1619729480
transform 0 -1 6429 1 0 1219
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_55959141808288  sky130_fd_io__tk_em1s_cdns_55959141808288_2
timestamp 1619729480
transform 0 1 6265 -1 0 567
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_0
timestamp 1619729480
transform -1 0 4746 0 1 1467
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_1
timestamp 1619729480
transform 0 1 5786 -1 0 511
box 0 24 144 28
use sky130_fd_io__feascom_pupredrvr_nbiasv2  sky130_fd_io__feascom_pupredrvr_nbiasv2_0
timestamp 1619729480
transform 1 0 831 0 1 165
box 0 36 3633 2349
use sky130_fd_io__gpiov2_pupredrvr_strong_nd2  sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0
timestamp 1619729480
transform -1 0 7072 0 1 0
box 0 7 1284 2632
use sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a  sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0
timestamp 1619729480
transform 1 0 4504 0 1 0
box 0 16 1284 2632
<< labels >>
flabel metal1 s -66 2284 -29 2430 3 FreeSans 300 0 0 0 VCC_IO
flabel metal1 s -66 1570 -24 1772 3 FreeSans 300 0 0 0 VCC_IO
flabel metal1 s 594 1044 636 1246 3 FreeSans 300 0 0 0 VGND_IO
flabel metal1 s 615 632 657 762 3 FreeSans 300 0 0 0 VGND_IO
flabel metal1 s 7036 2284 7072 2430 7 FreeSans 300 180 0 0 VCC_IO
flabel metal1 s 7036 1570 7072 1772 7 FreeSans 300 180 0 0 VCC_IO
flabel metal1 s 7036 1044 7072 1246 7 FreeSans 300 180 0 0 VGND_IO
flabel metal1 s 7036 632 7072 762 7 FreeSans 300 180 0 0 VGND_IO
flabel metal1 s 7036 2228 7072 2256 7 FreeSans 300 180 0 0 DRVHI_H
flabel metal1 s 7036 1800 7072 1846 7 FreeSans 300 180 0 0 PU_H_N[3]
flabel metal1 s 7036 2072 7072 2100 7 FreeSans 300 180 0 0 PUEN_H
flabel metal1 s 4504 1800 4540 1846 1 FreeSans 300 0 0 0 PU_H_N[2]
flabel metal1 s 5700 1800 5740 1846 2 FreeSans 300 180 0 0 PU_H_N[2]
flabel metal1 s 5836 1800 5877 1846 2 FreeSans 300 0 0 0 PU_H_N[3]
flabel metal1 s 0 2022 36 2068 7 FreeSans 300 180 0 0 PUEN_H
flabel metal1 s 318 1496 355 1542 7 FreeSans 300 180 0 0 SLOW_H_N
flabel comment s 678 397 678 397 0 FreeSans 300 0 0 0 EN_FAST_H_N
flabel comment s 884 1978 884 1978 0 FreeSans 300 0 0 0 EN_FAST_H
flabel comment s 947 469 947 469 0 FreeSans 300 0 0 0 EN_FAST_H
flabel comment s 5153 521 5153 521 0 FreeSans 300 180 0 0 EN_FAST_H
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 17502000
string GDS_START 17487592
<< end >>
