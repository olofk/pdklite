magic
tech sky130A
magscale 1 2
timestamp 1640697850
<< dnwell >>
rect -56 -102 4164 3162
<< nwell >>
rect 5197 1909 7274 2075
rect 18258 1213 19829 2127
rect 22582 1913 23468 2225
rect 23537 1913 23774 2225
rect 22582 1893 23820 1913
rect 22706 1581 23820 1893
rect 5192 -303 8093 583
rect 15799 -263 17119 -97
rect 6560 -322 6992 -303
rect 7039 -313 7601 -303
<< pwell >>
rect 3772 1847 4024 2654
rect 22798 2305 23252 2497
rect 3268 1495 4024 1847
rect 3772 1481 4024 1495
rect 3270 1094 3997 1296
rect 23980 1744 24066 2513
rect 22746 1265 23024 1502
rect 23502 1265 23780 1502
rect 22601 1177 23870 1265
rect 22395 1143 23870 1177
rect 3392 871 3742 1094
rect 3392 531 3990 871
rect 21825 839 23870 1143
rect 21825 765 22447 839
rect 3854 65 3990 531
rect 21586 187 22447 765
<< mvnmos >>
rect 3798 2475 3998 2575
rect 22877 2331 22997 2471
rect 23053 2331 23173 2471
rect 3798 2196 3998 2296
rect 3798 2040 3998 2140
rect 3347 1521 3447 1821
rect 3503 1521 3603 1821
rect 3798 1716 3998 1816
rect 3798 1560 3998 1660
rect 22825 1336 22945 1476
rect 23581 1336 23701 1476
rect 3349 1120 3449 1270
rect 3662 1120 3762 1270
rect 3818 1120 3918 1270
rect 3418 786 3502 906
rect 3632 786 3716 906
rect 3418 610 3502 730
rect 3632 610 3716 730
rect 3880 672 3964 792
rect 3880 496 3964 616
rect 3880 320 3964 440
rect 3880 144 3964 264
<< mvpmos >>
rect 22701 1959 22821 2159
rect 22877 1959 22997 2159
rect 23053 1959 23173 2159
rect 23229 1959 23349 2159
rect 22825 1647 22945 1847
rect 23025 1647 23145 1847
rect 23405 1647 23525 1847
rect 23581 1647 23701 1847
rect 5258 344 5458 464
rect 5258 168 5458 288
rect 6211 344 6411 464
rect 6211 168 6411 288
rect 6626 233 6926 333
rect 5258 -8 5458 112
rect 5258 -184 5458 -64
rect 6211 -8 6411 112
rect 6626 -47 6926 53
rect 6211 -184 6411 -64
rect 6626 -203 6926 -103
rect 7105 -194 7255 206
rect 7385 -194 7535 206
<< mvndiff >>
rect 3798 2620 3998 2628
rect 3798 2586 3816 2620
rect 3850 2586 3884 2620
rect 3918 2586 3952 2620
rect 3986 2586 3998 2620
rect 3798 2575 3998 2586
rect 3798 2464 3998 2475
rect 3798 2430 3816 2464
rect 3850 2430 3884 2464
rect 3918 2430 3952 2464
rect 3986 2430 3998 2464
rect 3798 2422 3998 2430
rect 22824 2459 22877 2471
rect 22824 2425 22832 2459
rect 22866 2425 22877 2459
rect 22824 2391 22877 2425
rect 22824 2357 22832 2391
rect 22866 2357 22877 2391
rect 3798 2341 3998 2349
rect 3798 2307 3816 2341
rect 3850 2307 3884 2341
rect 3918 2307 3952 2341
rect 3986 2307 3998 2341
rect 22824 2331 22877 2357
rect 22997 2459 23053 2471
rect 22997 2425 23008 2459
rect 23042 2425 23053 2459
rect 22997 2391 23053 2425
rect 22997 2357 23008 2391
rect 23042 2357 23053 2391
rect 22997 2331 23053 2357
rect 23173 2459 23226 2471
rect 23173 2425 23184 2459
rect 23218 2425 23226 2459
rect 23173 2391 23226 2425
rect 23173 2357 23184 2391
rect 23218 2357 23226 2391
rect 23173 2331 23226 2357
rect 3798 2296 3998 2307
rect 3798 2185 3998 2196
rect 3798 2151 3816 2185
rect 3850 2151 3884 2185
rect 3918 2151 3952 2185
rect 3986 2151 3998 2185
rect 3798 2140 3998 2151
rect 3798 2029 3998 2040
rect 3798 1995 3816 2029
rect 3850 1995 3884 2029
rect 3918 1995 3952 2029
rect 3986 1995 3998 2029
rect 3798 1987 3998 1995
rect 3798 1861 3998 1869
rect 3798 1827 3810 1861
rect 3844 1827 3878 1861
rect 3912 1827 3946 1861
rect 3980 1827 3998 1861
rect 3294 1771 3347 1821
rect 3294 1737 3302 1771
rect 3336 1737 3347 1771
rect 3294 1703 3347 1737
rect 3294 1669 3302 1703
rect 3336 1669 3347 1703
rect 3294 1635 3347 1669
rect 3294 1601 3302 1635
rect 3336 1601 3347 1635
rect 3294 1567 3347 1601
rect 3294 1533 3302 1567
rect 3336 1533 3347 1567
rect 3294 1521 3347 1533
rect 3447 1771 3503 1821
rect 3447 1737 3458 1771
rect 3492 1737 3503 1771
rect 3447 1703 3503 1737
rect 3447 1669 3458 1703
rect 3492 1669 3503 1703
rect 3447 1635 3503 1669
rect 3447 1601 3458 1635
rect 3492 1601 3503 1635
rect 3447 1567 3503 1601
rect 3447 1533 3458 1567
rect 3492 1533 3503 1567
rect 3447 1521 3503 1533
rect 3603 1771 3656 1821
rect 3798 1816 3998 1827
rect 3603 1737 3614 1771
rect 3648 1737 3656 1771
rect 3603 1703 3656 1737
rect 3603 1669 3614 1703
rect 3648 1669 3656 1703
rect 3603 1635 3656 1669
rect 3798 1705 3998 1716
rect 3798 1671 3810 1705
rect 3844 1671 3878 1705
rect 3912 1671 3946 1705
rect 3980 1671 3998 1705
rect 3798 1660 3998 1671
rect 3603 1601 3614 1635
rect 3648 1601 3656 1635
rect 3603 1567 3656 1601
rect 3603 1533 3614 1567
rect 3648 1533 3656 1567
rect 3603 1521 3656 1533
rect 3798 1549 3998 1560
rect 3798 1515 3810 1549
rect 3844 1515 3878 1549
rect 3912 1515 3946 1549
rect 3980 1515 3998 1549
rect 3798 1507 3998 1515
rect 22772 1450 22825 1476
rect 22772 1416 22780 1450
rect 22814 1416 22825 1450
rect 22772 1382 22825 1416
rect 22772 1348 22780 1382
rect 22814 1348 22825 1382
rect 22772 1336 22825 1348
rect 22945 1450 22998 1476
rect 22945 1416 22956 1450
rect 22990 1416 22998 1450
rect 22945 1382 22998 1416
rect 22945 1348 22956 1382
rect 22990 1348 22998 1382
rect 22945 1336 22998 1348
rect 23528 1450 23581 1476
rect 23528 1416 23536 1450
rect 23570 1416 23581 1450
rect 23528 1382 23581 1416
rect 23528 1348 23536 1382
rect 23570 1348 23581 1382
rect 23528 1336 23581 1348
rect 23701 1450 23754 1476
rect 23701 1416 23712 1450
rect 23746 1416 23754 1450
rect 23701 1382 23754 1416
rect 23701 1348 23712 1382
rect 23746 1348 23754 1382
rect 23701 1336 23754 1348
rect 3296 1234 3349 1270
rect 3296 1200 3304 1234
rect 3338 1200 3349 1234
rect 3296 1166 3349 1200
rect 3296 1132 3304 1166
rect 3338 1132 3349 1166
rect 3296 1120 3349 1132
rect 3449 1234 3502 1270
rect 3449 1200 3460 1234
rect 3494 1200 3502 1234
rect 3449 1166 3502 1200
rect 3449 1132 3460 1166
rect 3494 1132 3502 1166
rect 3449 1120 3502 1132
rect 3609 1258 3662 1270
rect 3609 1224 3617 1258
rect 3651 1224 3662 1258
rect 3609 1190 3662 1224
rect 3609 1156 3617 1190
rect 3651 1156 3662 1190
rect 3609 1120 3662 1156
rect 3762 1258 3818 1270
rect 3762 1224 3773 1258
rect 3807 1224 3818 1258
rect 3762 1190 3818 1224
rect 3762 1156 3773 1190
rect 3807 1156 3818 1190
rect 3762 1120 3818 1156
rect 3918 1258 3971 1270
rect 3918 1224 3929 1258
rect 3963 1224 3971 1258
rect 3918 1190 3971 1224
rect 3918 1156 3929 1190
rect 3963 1156 3971 1190
rect 3918 1120 3971 1156
rect 3418 951 3502 959
rect 3418 917 3430 951
rect 3464 917 3502 951
rect 3418 906 3502 917
rect 3632 951 3716 959
rect 3632 917 3644 951
rect 3678 917 3716 951
rect 3632 906 3716 917
rect 3418 775 3502 786
rect 3418 741 3430 775
rect 3464 741 3502 775
rect 3418 730 3502 741
rect 3880 837 3964 845
rect 3880 803 3892 837
rect 3926 803 3964 837
rect 3880 792 3964 803
rect 3632 775 3716 786
rect 3632 741 3644 775
rect 3678 741 3716 775
rect 3632 730 3716 741
rect 3880 661 3964 672
rect 3880 627 3892 661
rect 3926 627 3964 661
rect 3880 616 3964 627
rect 3418 599 3502 610
rect 3418 565 3430 599
rect 3464 565 3502 599
rect 3418 557 3502 565
rect 3632 599 3716 610
rect 3632 565 3644 599
rect 3678 565 3716 599
rect 3632 557 3716 565
rect 3880 485 3964 496
rect 3880 451 3892 485
rect 3926 451 3964 485
rect 3880 440 3964 451
rect 3880 309 3964 320
rect 3880 275 3892 309
rect 3926 275 3964 309
rect 3880 264 3964 275
rect 3880 133 3964 144
rect 3880 99 3892 133
rect 3926 99 3964 133
rect 3880 91 3964 99
<< mvpdiff >>
rect 22648 2141 22701 2159
rect 22648 2107 22656 2141
rect 22690 2107 22701 2141
rect 22648 2073 22701 2107
rect 22648 2039 22656 2073
rect 22690 2039 22701 2073
rect 22648 2005 22701 2039
rect 22648 1971 22656 2005
rect 22690 1971 22701 2005
rect 22648 1959 22701 1971
rect 22821 2141 22877 2159
rect 22821 2107 22832 2141
rect 22866 2107 22877 2141
rect 22821 2073 22877 2107
rect 22821 2039 22832 2073
rect 22866 2039 22877 2073
rect 22821 2005 22877 2039
rect 22821 1971 22832 2005
rect 22866 1971 22877 2005
rect 22821 1959 22877 1971
rect 22997 2141 23053 2159
rect 22997 2107 23008 2141
rect 23042 2107 23053 2141
rect 22997 2073 23053 2107
rect 22997 2039 23008 2073
rect 23042 2039 23053 2073
rect 22997 2005 23053 2039
rect 22997 1971 23008 2005
rect 23042 1971 23053 2005
rect 22997 1959 23053 1971
rect 23173 2141 23229 2159
rect 23173 2107 23184 2141
rect 23218 2107 23229 2141
rect 23173 2073 23229 2107
rect 23173 2039 23184 2073
rect 23218 2039 23229 2073
rect 23173 2005 23229 2039
rect 23173 1971 23184 2005
rect 23218 1971 23229 2005
rect 23173 1959 23229 1971
rect 23349 2141 23402 2159
rect 23349 2107 23360 2141
rect 23394 2107 23402 2141
rect 23349 2073 23402 2107
rect 23349 2039 23360 2073
rect 23394 2039 23402 2073
rect 23349 2005 23402 2039
rect 23349 1971 23360 2005
rect 23394 1971 23402 2005
rect 23349 1959 23402 1971
rect 22772 1829 22825 1847
rect 22772 1795 22780 1829
rect 22814 1795 22825 1829
rect 22772 1761 22825 1795
rect 22772 1727 22780 1761
rect 22814 1727 22825 1761
rect 22772 1693 22825 1727
rect 22772 1659 22780 1693
rect 22814 1659 22825 1693
rect 22772 1647 22825 1659
rect 22945 1829 23025 1847
rect 22945 1795 22968 1829
rect 23002 1795 23025 1829
rect 22945 1761 23025 1795
rect 22945 1727 22968 1761
rect 23002 1727 23025 1761
rect 22945 1693 23025 1727
rect 22945 1659 22968 1693
rect 23002 1659 23025 1693
rect 22945 1647 23025 1659
rect 23145 1829 23205 1847
rect 23345 1829 23405 1847
rect 23145 1795 23156 1829
rect 23190 1795 23205 1829
rect 23345 1795 23360 1829
rect 23394 1795 23405 1829
rect 23145 1761 23205 1795
rect 23345 1761 23405 1795
rect 23145 1727 23156 1761
rect 23190 1727 23205 1761
rect 23345 1727 23360 1761
rect 23394 1727 23405 1761
rect 23145 1693 23205 1727
rect 23345 1693 23405 1727
rect 23145 1659 23156 1693
rect 23190 1659 23205 1693
rect 23345 1659 23360 1693
rect 23394 1659 23405 1693
rect 23145 1647 23205 1659
rect 23345 1647 23405 1659
rect 23525 1829 23581 1847
rect 23525 1795 23536 1829
rect 23570 1795 23581 1829
rect 23525 1761 23581 1795
rect 23525 1727 23536 1761
rect 23570 1727 23581 1761
rect 23525 1693 23581 1727
rect 23525 1659 23536 1693
rect 23570 1659 23581 1693
rect 23525 1647 23581 1659
rect 23701 1829 23754 1847
rect 23701 1795 23712 1829
rect 23746 1795 23754 1829
rect 23701 1761 23754 1795
rect 23701 1727 23712 1761
rect 23746 1727 23754 1761
rect 23701 1693 23754 1727
rect 23701 1659 23712 1693
rect 23746 1659 23754 1693
rect 23701 1647 23754 1659
rect 5258 509 5458 517
rect 5258 475 5270 509
rect 5304 475 5338 509
rect 5372 475 5406 509
rect 5440 475 5458 509
rect 5258 464 5458 475
rect 6211 509 6411 517
rect 6211 475 6229 509
rect 6263 475 6297 509
rect 6331 475 6365 509
rect 6399 475 6411 509
rect 6211 464 6411 475
rect 5258 333 5458 344
rect 5258 299 5270 333
rect 5304 299 5338 333
rect 5372 299 5406 333
rect 5440 299 5458 333
rect 5258 288 5458 299
rect 6626 378 6926 386
rect 6211 333 6411 344
rect 6211 299 6229 333
rect 6263 299 6297 333
rect 6331 299 6365 333
rect 6399 299 6411 333
rect 6211 288 6411 299
rect 6626 344 6638 378
rect 6672 344 6706 378
rect 6740 344 6774 378
rect 6808 344 6842 378
rect 6876 344 6926 378
rect 6626 333 6926 344
rect 7105 251 7255 259
rect 6626 222 6926 233
rect 6626 188 6638 222
rect 6672 188 6706 222
rect 6740 188 6774 222
rect 6808 188 6842 222
rect 6876 188 6926 222
rect 7105 217 7117 251
rect 7151 217 7185 251
rect 7219 217 7255 251
rect 7105 206 7255 217
rect 7385 251 7535 259
rect 7385 217 7397 251
rect 7431 217 7465 251
rect 7499 217 7535 251
rect 7385 206 7535 217
rect 6626 180 6926 188
rect 5258 157 5458 168
rect 5258 123 5270 157
rect 5304 123 5338 157
rect 5372 123 5406 157
rect 5440 123 5458 157
rect 5258 112 5458 123
rect 6211 157 6411 168
rect 6211 123 6229 157
rect 6263 123 6297 157
rect 6331 123 6365 157
rect 6399 123 6411 157
rect 6211 112 6411 123
rect 5258 -19 5458 -8
rect 5258 -53 5270 -19
rect 5304 -53 5338 -19
rect 5372 -53 5406 -19
rect 5440 -53 5458 -19
rect 5258 -64 5458 -53
rect 6626 98 6926 106
rect 6626 64 6638 98
rect 6672 64 6706 98
rect 6740 64 6774 98
rect 6808 64 6842 98
rect 6876 64 6926 98
rect 6626 53 6926 64
rect 6211 -19 6411 -8
rect 6211 -53 6229 -19
rect 6263 -53 6297 -19
rect 6331 -53 6365 -19
rect 6399 -53 6411 -19
rect 6211 -64 6411 -53
rect 6626 -58 6926 -47
rect 6626 -92 6638 -58
rect 6672 -92 6706 -58
rect 6740 -92 6774 -58
rect 6808 -92 6842 -58
rect 6876 -92 6926 -58
rect 6626 -103 6926 -92
rect 5258 -195 5458 -184
rect 5258 -229 5270 -195
rect 5304 -229 5338 -195
rect 5372 -229 5406 -195
rect 5440 -229 5458 -195
rect 6211 -195 6411 -184
rect 5258 -237 5458 -229
rect 6211 -229 6229 -195
rect 6263 -229 6297 -195
rect 6331 -229 6365 -195
rect 6399 -229 6411 -195
rect 6211 -237 6411 -229
rect 6626 -214 6926 -203
rect 6626 -248 6638 -214
rect 6672 -248 6706 -214
rect 6740 -248 6774 -214
rect 6808 -248 6842 -214
rect 6876 -248 6926 -214
rect 7105 -205 7255 -194
rect 7105 -239 7117 -205
rect 7151 -239 7185 -205
rect 7219 -239 7255 -205
rect 7105 -247 7255 -239
rect 7385 -205 7535 -194
rect 7385 -239 7397 -205
rect 7431 -239 7465 -205
rect 7499 -239 7535 -205
rect 7385 -247 7535 -239
rect 6626 -256 6926 -248
<< mvndiffc >>
rect 3816 2586 3850 2620
rect 3884 2586 3918 2620
rect 3952 2586 3986 2620
rect 3816 2430 3850 2464
rect 3884 2430 3918 2464
rect 3952 2430 3986 2464
rect 22832 2425 22866 2459
rect 22832 2357 22866 2391
rect 3816 2307 3850 2341
rect 3884 2307 3918 2341
rect 3952 2307 3986 2341
rect 23008 2425 23042 2459
rect 23008 2357 23042 2391
rect 23184 2425 23218 2459
rect 23184 2357 23218 2391
rect 3816 2151 3850 2185
rect 3884 2151 3918 2185
rect 3952 2151 3986 2185
rect 3816 1995 3850 2029
rect 3884 1995 3918 2029
rect 3952 1995 3986 2029
rect 3810 1827 3844 1861
rect 3878 1827 3912 1861
rect 3946 1827 3980 1861
rect 3302 1737 3336 1771
rect 3302 1669 3336 1703
rect 3302 1601 3336 1635
rect 3302 1533 3336 1567
rect 3458 1737 3492 1771
rect 3458 1669 3492 1703
rect 3458 1601 3492 1635
rect 3458 1533 3492 1567
rect 3614 1737 3648 1771
rect 3614 1669 3648 1703
rect 3810 1671 3844 1705
rect 3878 1671 3912 1705
rect 3946 1671 3980 1705
rect 3614 1601 3648 1635
rect 3614 1533 3648 1567
rect 3810 1515 3844 1549
rect 3878 1515 3912 1549
rect 3946 1515 3980 1549
rect 22780 1416 22814 1450
rect 22780 1348 22814 1382
rect 22956 1416 22990 1450
rect 22956 1348 22990 1382
rect 23536 1416 23570 1450
rect 23536 1348 23570 1382
rect 23712 1416 23746 1450
rect 23712 1348 23746 1382
rect 3304 1200 3338 1234
rect 3304 1132 3338 1166
rect 3460 1200 3494 1234
rect 3460 1132 3494 1166
rect 3617 1224 3651 1258
rect 3617 1156 3651 1190
rect 3773 1224 3807 1258
rect 3773 1156 3807 1190
rect 3929 1224 3963 1258
rect 3929 1156 3963 1190
rect 3430 917 3464 951
rect 3644 917 3678 951
rect 3430 741 3464 775
rect 3892 803 3926 837
rect 3644 741 3678 775
rect 3892 627 3926 661
rect 3430 565 3464 599
rect 3644 565 3678 599
rect 3892 451 3926 485
rect 3892 275 3926 309
rect 3892 99 3926 133
<< mvpdiffc >>
rect 22656 2107 22690 2141
rect 22656 2039 22690 2073
rect 22656 1971 22690 2005
rect 22832 2107 22866 2141
rect 22832 2039 22866 2073
rect 22832 1971 22866 2005
rect 23008 2107 23042 2141
rect 23008 2039 23042 2073
rect 23008 1971 23042 2005
rect 23184 2107 23218 2141
rect 23184 2039 23218 2073
rect 23184 1971 23218 2005
rect 23360 2107 23394 2141
rect 23360 2039 23394 2073
rect 23360 1971 23394 2005
rect 22780 1795 22814 1829
rect 22780 1727 22814 1761
rect 22780 1659 22814 1693
rect 22968 1795 23002 1829
rect 22968 1727 23002 1761
rect 22968 1659 23002 1693
rect 23156 1795 23190 1829
rect 23360 1795 23394 1829
rect 23156 1727 23190 1761
rect 23360 1727 23394 1761
rect 23156 1659 23190 1693
rect 23360 1659 23394 1693
rect 23536 1795 23570 1829
rect 23536 1727 23570 1761
rect 23536 1659 23570 1693
rect 23712 1795 23746 1829
rect 23712 1727 23746 1761
rect 23712 1659 23746 1693
rect 5270 475 5304 509
rect 5338 475 5372 509
rect 5406 475 5440 509
rect 6229 475 6263 509
rect 6297 475 6331 509
rect 6365 475 6399 509
rect 5270 299 5304 333
rect 5338 299 5372 333
rect 5406 299 5440 333
rect 6229 299 6263 333
rect 6297 299 6331 333
rect 6365 299 6399 333
rect 6638 344 6672 378
rect 6706 344 6740 378
rect 6774 344 6808 378
rect 6842 344 6876 378
rect 6638 188 6672 222
rect 6706 188 6740 222
rect 6774 188 6808 222
rect 6842 188 6876 222
rect 7117 217 7151 251
rect 7185 217 7219 251
rect 7397 217 7431 251
rect 7465 217 7499 251
rect 5270 123 5304 157
rect 5338 123 5372 157
rect 5406 123 5440 157
rect 6229 123 6263 157
rect 6297 123 6331 157
rect 6365 123 6399 157
rect 5270 -53 5304 -19
rect 5338 -53 5372 -19
rect 5406 -53 5440 -19
rect 6638 64 6672 98
rect 6706 64 6740 98
rect 6774 64 6808 98
rect 6842 64 6876 98
rect 6229 -53 6263 -19
rect 6297 -53 6331 -19
rect 6365 -53 6399 -19
rect 6638 -92 6672 -58
rect 6706 -92 6740 -58
rect 6774 -92 6808 -58
rect 6842 -92 6876 -58
rect 5270 -229 5304 -195
rect 5338 -229 5372 -195
rect 5406 -229 5440 -195
rect 6229 -229 6263 -195
rect 6297 -229 6331 -195
rect 6365 -229 6399 -195
rect 6638 -248 6672 -214
rect 6706 -248 6740 -214
rect 6774 -248 6808 -214
rect 6842 -248 6876 -214
rect 7117 -239 7151 -205
rect 7185 -239 7219 -205
rect 7397 -239 7431 -205
rect 7465 -239 7499 -205
<< psubdiff >>
rect 24006 2463 24040 2487
rect 24006 2393 24040 2429
rect 24006 2323 24040 2359
rect 24006 2253 24040 2289
rect 24006 2183 24040 2219
rect 24006 2112 24040 2149
rect 24006 2041 24040 2078
rect 24006 1970 24040 2007
rect 24006 1899 24040 1936
rect 24006 1828 24040 1865
rect 24006 1770 24040 1794
rect 22639 1205 23844 1239
rect 22639 1171 22661 1205
rect 22695 1171 22731 1205
rect 22765 1171 22801 1205
rect 22835 1171 22871 1205
rect 22905 1171 22941 1205
rect 22975 1171 23011 1205
rect 23045 1171 23081 1205
rect 23115 1171 23151 1205
rect 23185 1171 23221 1205
rect 23255 1171 23291 1205
rect 23325 1171 23361 1205
rect 23395 1171 23431 1205
rect 23465 1171 23500 1205
rect 23534 1171 23569 1205
rect 23603 1171 23638 1205
rect 23672 1171 23707 1205
rect 23741 1171 23776 1205
rect 23810 1171 23844 1205
rect 22639 1137 23844 1171
rect 22639 1103 22661 1137
rect 22695 1103 22731 1137
rect 22765 1103 22801 1137
rect 22835 1103 22871 1137
rect 22905 1103 22941 1137
rect 22975 1103 23011 1137
rect 23045 1103 23081 1137
rect 23115 1103 23151 1137
rect 23185 1103 23221 1137
rect 23255 1103 23291 1137
rect 23325 1103 23361 1137
rect 23395 1103 23431 1137
rect 23465 1103 23500 1137
rect 23534 1103 23569 1137
rect 23603 1103 23638 1137
rect 23672 1103 23707 1137
rect 23741 1103 23776 1137
rect 23810 1103 23844 1137
rect 22639 1069 23844 1103
rect 22639 1035 22661 1069
rect 22695 1035 22731 1069
rect 22765 1035 22801 1069
rect 22835 1035 22871 1069
rect 22905 1035 22941 1069
rect 22975 1035 23011 1069
rect 23045 1035 23081 1069
rect 23115 1035 23151 1069
rect 23185 1035 23221 1069
rect 23255 1035 23291 1069
rect 23325 1035 23361 1069
rect 23395 1035 23431 1069
rect 23465 1035 23500 1069
rect 23534 1035 23569 1069
rect 23603 1035 23638 1069
rect 23672 1035 23707 1069
rect 23741 1035 23776 1069
rect 23810 1035 23844 1069
rect 22639 1001 23844 1035
rect 22639 967 22661 1001
rect 22695 967 22731 1001
rect 22765 967 22801 1001
rect 22835 967 22871 1001
rect 22905 967 22941 1001
rect 22975 967 23011 1001
rect 23045 967 23081 1001
rect 23115 967 23151 1001
rect 23185 967 23221 1001
rect 23255 967 23291 1001
rect 23325 967 23361 1001
rect 23395 967 23431 1001
rect 23465 967 23500 1001
rect 23534 967 23569 1001
rect 23603 967 23638 1001
rect 23672 967 23707 1001
rect 23741 967 23776 1001
rect 23810 967 23844 1001
rect 22639 933 23844 967
rect 22639 899 22661 933
rect 22695 899 22731 933
rect 22765 899 22801 933
rect 22835 899 22871 933
rect 22905 899 22941 933
rect 22975 899 23011 933
rect 23045 899 23081 933
rect 23115 899 23151 933
rect 23185 899 23221 933
rect 23255 899 23291 933
rect 23325 899 23361 933
rect 23395 899 23431 933
rect 23465 899 23500 933
rect 23534 899 23569 933
rect 23603 899 23638 933
rect 23672 899 23707 933
rect 23741 899 23776 933
rect 23810 899 23844 933
rect 22639 898 23844 899
rect 21851 865 22455 898
rect 22489 865 22559 898
rect 22593 865 23844 898
rect 21851 831 21853 865
rect 21887 831 21929 865
rect 21963 831 22005 865
rect 22039 831 22081 865
rect 22115 831 22157 865
rect 22191 831 22233 865
rect 22267 831 22309 865
rect 22343 831 22385 865
rect 22419 831 22421 865
rect 21851 792 22421 831
rect 21851 758 21853 792
rect 21887 758 21929 792
rect 21963 758 22005 792
rect 22039 758 22081 792
rect 22115 758 22157 792
rect 22191 758 22233 792
rect 22267 758 22309 792
rect 22343 758 22385 792
rect 22419 758 22421 792
rect 21851 739 22421 758
rect 21725 719 22421 739
rect 21725 685 21853 719
rect 21887 685 21929 719
rect 21963 685 22005 719
rect 22039 685 22081 719
rect 22115 685 22157 719
rect 22191 685 22233 719
rect 22267 685 22309 719
rect 22343 685 22385 719
rect 22419 685 22421 719
rect 21725 646 22421 685
rect 21725 612 21853 646
rect 21887 612 21929 646
rect 21963 612 22005 646
rect 22039 612 22081 646
rect 22115 612 22157 646
rect 22191 612 22233 646
rect 22267 612 22309 646
rect 22343 612 22385 646
rect 22419 612 22421 646
rect 21725 573 22421 612
rect 21725 539 21853 573
rect 21887 539 21929 573
rect 21963 539 22005 573
rect 22039 539 22081 573
rect 22115 539 22157 573
rect 22191 539 22233 573
rect 22267 539 22309 573
rect 22343 539 22385 573
rect 22419 539 22421 573
rect 21725 500 22421 539
rect 21725 466 21853 500
rect 21887 466 21929 500
rect 21963 466 22005 500
rect 22039 466 22081 500
rect 22115 466 22157 500
rect 22191 466 22233 500
rect 22267 466 22309 500
rect 22343 466 22385 500
rect 22419 466 22421 500
rect 21725 427 22421 466
rect 21725 393 21853 427
rect 21887 393 21929 427
rect 21963 393 22005 427
rect 22039 393 22081 427
rect 22115 393 22157 427
rect 22191 393 22233 427
rect 22267 393 22309 427
rect 22343 393 22385 427
rect 22419 393 22421 427
rect 21725 354 22421 393
rect 21725 320 21853 354
rect 21887 320 21929 354
rect 21963 320 22005 354
rect 22039 320 22081 354
rect 22115 320 22157 354
rect 22191 320 22233 354
rect 22267 320 22309 354
rect 22343 320 22385 354
rect 22419 320 22421 354
rect 21725 281 22421 320
rect 21725 247 21853 281
rect 21887 247 21929 281
rect 21963 247 22005 281
rect 22039 247 22081 281
rect 22115 247 22157 281
rect 22191 247 22233 281
rect 22267 247 22309 281
rect 22343 247 22385 281
rect 22419 247 22421 281
rect 21725 213 22421 247
<< mvpsubdiff >>
rect 22627 1151 22639 1239
rect 22421 1117 22455 1151
rect 22489 1117 22559 1151
rect 22593 1117 22639 1151
rect 21851 1083 22639 1117
rect 21851 1049 21853 1083
rect 21887 1049 21929 1083
rect 21963 1049 22005 1083
rect 22039 1049 22081 1083
rect 22115 1049 22157 1083
rect 22191 1049 22233 1083
rect 22267 1049 22309 1083
rect 22343 1049 22385 1083
rect 22419 1067 22639 1083
rect 22419 1049 22455 1067
rect 21851 1033 22455 1049
rect 22489 1033 22559 1067
rect 22593 1033 22639 1067
rect 21851 1011 22639 1033
rect 21851 977 21853 1011
rect 21887 977 21929 1011
rect 21963 977 22005 1011
rect 22039 977 22081 1011
rect 22115 977 22157 1011
rect 22191 977 22233 1011
rect 22267 977 22309 1011
rect 22343 977 22385 1011
rect 22419 983 22639 1011
rect 22419 977 22455 983
rect 21851 949 22455 977
rect 22489 949 22559 983
rect 22593 949 22639 983
rect 21851 938 22639 949
rect 21851 904 21853 938
rect 21887 904 21929 938
rect 21963 904 22005 938
rect 22039 904 22081 938
rect 22115 904 22157 938
rect 22191 904 22233 938
rect 22267 904 22309 938
rect 22343 904 22385 938
rect 22419 904 22639 938
rect 21851 899 22639 904
rect 21851 898 22455 899
rect 22489 898 22559 899
rect 22593 898 22639 899
<< mvnsubdiff >>
rect 5263 1975 5287 2009
rect 5321 1975 5356 2009
rect 5390 1975 5425 2009
rect 5459 1975 5494 2009
rect 5528 1975 5563 2009
rect 5597 1975 5632 2009
rect 5666 1975 5701 2009
rect 5735 1975 5770 2009
rect 5804 1975 5839 2009
rect 5873 1975 5908 2009
rect 5942 1975 5977 2009
rect 6011 1975 6046 2009
rect 6080 1975 6115 2009
rect 6149 1975 6184 2009
rect 6218 1975 6253 2009
rect 6287 1975 6322 2009
rect 6356 1975 6391 2009
rect 6425 1975 6460 2009
rect 6494 1975 6529 2009
rect 6563 1975 6598 2009
rect 6632 1975 6667 2009
rect 6701 1975 6736 2009
rect 6770 1975 6805 2009
rect 6839 1975 6874 2009
rect 6908 1975 6943 2009
rect 6977 1975 7012 2009
rect 7046 1975 7081 2009
rect 7115 1975 7150 2009
rect 7184 1975 7208 2009
rect 5263 1941 7208 1975
rect 23205 1829 23345 1847
rect 23205 1795 23258 1829
rect 23292 1795 23345 1829
rect 23205 1761 23345 1795
rect 23205 1727 23258 1761
rect 23292 1727 23345 1761
rect 23205 1693 23345 1727
rect 23205 1659 23258 1693
rect 23292 1659 23345 1693
rect 23205 1647 23345 1659
rect 6529 478 6553 512
rect 6587 478 6628 512
rect 6662 478 6703 512
rect 6737 478 6778 512
rect 6812 478 6853 512
rect 6887 478 6927 512
rect 6961 478 6985 512
rect 5584 -237 5608 -203
rect 5642 -237 5683 -203
rect 5717 -237 5758 -203
rect 5792 -237 5833 -203
rect 5867 -237 5908 -203
rect 5942 -237 5982 -203
rect 6016 -237 6040 -203
rect 15865 -197 15889 -163
rect 15923 -197 15959 -163
rect 15993 -197 16029 -163
rect 16063 -197 16098 -163
rect 16132 -197 16167 -163
rect 16201 -197 16236 -163
rect 16270 -197 16305 -163
rect 16339 -197 16374 -163
rect 16408 -197 16443 -163
rect 16477 -197 16512 -163
rect 16546 -197 16581 -163
rect 16615 -197 16650 -163
rect 16684 -197 16719 -163
rect 16753 -197 16788 -163
rect 16822 -197 16857 -163
rect 16891 -197 16926 -163
rect 16960 -197 16995 -163
rect 17029 -197 17053 -163
<< psubdiffcont >>
rect 24006 2429 24040 2463
rect 24006 2359 24040 2393
rect 24006 2289 24040 2323
rect 24006 2219 24040 2253
rect 24006 2149 24040 2183
rect 24006 2078 24040 2112
rect 24006 2007 24040 2041
rect 24006 1936 24040 1970
rect 24006 1865 24040 1899
rect 24006 1794 24040 1828
rect 22661 1171 22695 1205
rect 22731 1171 22765 1205
rect 22801 1171 22835 1205
rect 22871 1171 22905 1205
rect 22941 1171 22975 1205
rect 23011 1171 23045 1205
rect 23081 1171 23115 1205
rect 23151 1171 23185 1205
rect 23221 1171 23255 1205
rect 23291 1171 23325 1205
rect 23361 1171 23395 1205
rect 23431 1171 23465 1205
rect 23500 1171 23534 1205
rect 23569 1171 23603 1205
rect 23638 1171 23672 1205
rect 23707 1171 23741 1205
rect 23776 1171 23810 1205
rect 22661 1103 22695 1137
rect 22731 1103 22765 1137
rect 22801 1103 22835 1137
rect 22871 1103 22905 1137
rect 22941 1103 22975 1137
rect 23011 1103 23045 1137
rect 23081 1103 23115 1137
rect 23151 1103 23185 1137
rect 23221 1103 23255 1137
rect 23291 1103 23325 1137
rect 23361 1103 23395 1137
rect 23431 1103 23465 1137
rect 23500 1103 23534 1137
rect 23569 1103 23603 1137
rect 23638 1103 23672 1137
rect 23707 1103 23741 1137
rect 23776 1103 23810 1137
rect 22661 1035 22695 1069
rect 22731 1035 22765 1069
rect 22801 1035 22835 1069
rect 22871 1035 22905 1069
rect 22941 1035 22975 1069
rect 23011 1035 23045 1069
rect 23081 1035 23115 1069
rect 23151 1035 23185 1069
rect 23221 1035 23255 1069
rect 23291 1035 23325 1069
rect 23361 1035 23395 1069
rect 23431 1035 23465 1069
rect 23500 1035 23534 1069
rect 23569 1035 23603 1069
rect 23638 1035 23672 1069
rect 23707 1035 23741 1069
rect 23776 1035 23810 1069
rect 22661 967 22695 1001
rect 22731 967 22765 1001
rect 22801 967 22835 1001
rect 22871 967 22905 1001
rect 22941 967 22975 1001
rect 23011 967 23045 1001
rect 23081 967 23115 1001
rect 23151 967 23185 1001
rect 23221 967 23255 1001
rect 23291 967 23325 1001
rect 23361 967 23395 1001
rect 23431 967 23465 1001
rect 23500 967 23534 1001
rect 23569 967 23603 1001
rect 23638 967 23672 1001
rect 23707 967 23741 1001
rect 23776 967 23810 1001
rect 22661 899 22695 933
rect 22731 899 22765 933
rect 22801 899 22835 933
rect 22871 899 22905 933
rect 22941 899 22975 933
rect 23011 899 23045 933
rect 23081 899 23115 933
rect 23151 899 23185 933
rect 23221 899 23255 933
rect 23291 899 23325 933
rect 23361 899 23395 933
rect 23431 899 23465 933
rect 23500 899 23534 933
rect 23569 899 23603 933
rect 23638 899 23672 933
rect 23707 899 23741 933
rect 23776 899 23810 933
rect 22455 865 22489 898
rect 22559 865 22593 898
rect 21853 831 21887 865
rect 21929 831 21963 865
rect 22005 831 22039 865
rect 22081 831 22115 865
rect 22157 831 22191 865
rect 22233 831 22267 865
rect 22309 831 22343 865
rect 22385 831 22419 865
rect 21853 758 21887 792
rect 21929 758 21963 792
rect 22005 758 22039 792
rect 22081 758 22115 792
rect 22157 758 22191 792
rect 22233 758 22267 792
rect 22309 758 22343 792
rect 22385 758 22419 792
rect 21853 685 21887 719
rect 21929 685 21963 719
rect 22005 685 22039 719
rect 22081 685 22115 719
rect 22157 685 22191 719
rect 22233 685 22267 719
rect 22309 685 22343 719
rect 22385 685 22419 719
rect 21853 612 21887 646
rect 21929 612 21963 646
rect 22005 612 22039 646
rect 22081 612 22115 646
rect 22157 612 22191 646
rect 22233 612 22267 646
rect 22309 612 22343 646
rect 22385 612 22419 646
rect 21853 539 21887 573
rect 21929 539 21963 573
rect 22005 539 22039 573
rect 22081 539 22115 573
rect 22157 539 22191 573
rect 22233 539 22267 573
rect 22309 539 22343 573
rect 22385 539 22419 573
rect 21853 466 21887 500
rect 21929 466 21963 500
rect 22005 466 22039 500
rect 22081 466 22115 500
rect 22157 466 22191 500
rect 22233 466 22267 500
rect 22309 466 22343 500
rect 22385 466 22419 500
rect 21853 393 21887 427
rect 21929 393 21963 427
rect 22005 393 22039 427
rect 22081 393 22115 427
rect 22157 393 22191 427
rect 22233 393 22267 427
rect 22309 393 22343 427
rect 22385 393 22419 427
rect 21853 320 21887 354
rect 21929 320 21963 354
rect 22005 320 22039 354
rect 22081 320 22115 354
rect 22157 320 22191 354
rect 22233 320 22267 354
rect 22309 320 22343 354
rect 22385 320 22419 354
rect 21853 247 21887 281
rect 21929 247 21963 281
rect 22005 247 22039 281
rect 22081 247 22115 281
rect 22157 247 22191 281
rect 22233 247 22267 281
rect 22309 247 22343 281
rect 22385 247 22419 281
<< mvpsubdiffcont >>
rect 22455 1117 22489 1151
rect 22559 1117 22593 1151
rect 21853 1049 21887 1083
rect 21929 1049 21963 1083
rect 22005 1049 22039 1083
rect 22081 1049 22115 1083
rect 22157 1049 22191 1083
rect 22233 1049 22267 1083
rect 22309 1049 22343 1083
rect 22385 1049 22419 1083
rect 22455 1033 22489 1067
rect 22559 1033 22593 1067
rect 21853 977 21887 1011
rect 21929 977 21963 1011
rect 22005 977 22039 1011
rect 22081 977 22115 1011
rect 22157 977 22191 1011
rect 22233 977 22267 1011
rect 22309 977 22343 1011
rect 22385 977 22419 1011
rect 22455 949 22489 983
rect 22559 949 22593 983
rect 21853 904 21887 938
rect 21929 904 21963 938
rect 22005 904 22039 938
rect 22081 904 22115 938
rect 22157 904 22191 938
rect 22233 904 22267 938
rect 22309 904 22343 938
rect 22385 904 22419 938
rect 22455 898 22489 899
rect 22559 898 22593 899
<< mvnsubdiffcont >>
rect 5287 1975 5321 2009
rect 5356 1975 5390 2009
rect 5425 1975 5459 2009
rect 5494 1975 5528 2009
rect 5563 1975 5597 2009
rect 5632 1975 5666 2009
rect 5701 1975 5735 2009
rect 5770 1975 5804 2009
rect 5839 1975 5873 2009
rect 5908 1975 5942 2009
rect 5977 1975 6011 2009
rect 6046 1975 6080 2009
rect 6115 1975 6149 2009
rect 6184 1975 6218 2009
rect 6253 1975 6287 2009
rect 6322 1975 6356 2009
rect 6391 1975 6425 2009
rect 6460 1975 6494 2009
rect 6529 1975 6563 2009
rect 6598 1975 6632 2009
rect 6667 1975 6701 2009
rect 6736 1975 6770 2009
rect 6805 1975 6839 2009
rect 6874 1975 6908 2009
rect 6943 1975 6977 2009
rect 7012 1975 7046 2009
rect 7081 1975 7115 2009
rect 7150 1975 7184 2009
rect 23258 1795 23292 1829
rect 23258 1727 23292 1761
rect 23258 1659 23292 1693
rect 6553 478 6587 512
rect 6628 478 6662 512
rect 6703 478 6737 512
rect 6778 478 6812 512
rect 6853 478 6887 512
rect 6927 478 6961 512
rect 5608 -237 5642 -203
rect 5683 -237 5717 -203
rect 5758 -237 5792 -203
rect 5833 -237 5867 -203
rect 5908 -237 5942 -203
rect 5982 -237 6016 -203
rect 15889 -197 15923 -163
rect 15959 -197 15993 -163
rect 16029 -197 16063 -163
rect 16098 -197 16132 -163
rect 16167 -197 16201 -163
rect 16236 -197 16270 -163
rect 16305 -197 16339 -163
rect 16374 -197 16408 -163
rect 16443 -197 16477 -163
rect 16512 -197 16546 -163
rect 16581 -197 16615 -163
rect 16650 -197 16684 -163
rect 16719 -197 16753 -163
rect 16788 -197 16822 -163
rect 16857 -197 16891 -163
rect 16926 -197 16960 -163
rect 16995 -197 17029 -163
<< poly >>
rect 4030 2593 4096 2609
rect 4030 2575 4046 2593
rect 3766 2475 3798 2575
rect 3998 2559 4046 2575
rect 4080 2559 4096 2593
rect 3998 2525 4096 2559
rect 3998 2491 4046 2525
rect 4080 2491 4096 2525
rect 3998 2475 4096 2491
rect 22877 2471 22997 2503
rect 23053 2471 23173 2503
rect 22877 2299 22997 2331
rect 3766 2196 3798 2296
rect 3998 2255 4096 2296
rect 3998 2221 4046 2255
rect 4080 2221 4096 2255
rect 3998 2196 4096 2221
rect 4030 2173 4096 2196
rect 4030 2140 4046 2173
rect 3766 2040 3798 2140
rect 3998 2139 4046 2140
rect 4080 2139 4096 2173
rect 22701 2267 22997 2299
rect 22701 2233 22721 2267
rect 22755 2233 22795 2267
rect 22829 2233 22869 2267
rect 22903 2233 22943 2267
rect 22977 2233 22997 2267
rect 22701 2202 22997 2233
rect 22701 2159 22821 2202
rect 22877 2159 22997 2202
rect 23053 2299 23173 2331
rect 23053 2267 23349 2299
rect 23053 2233 23073 2267
rect 23107 2233 23147 2267
rect 23181 2233 23221 2267
rect 23255 2233 23295 2267
rect 23329 2233 23349 2267
rect 23053 2202 23349 2233
rect 23053 2159 23173 2202
rect 23229 2159 23349 2202
rect 3998 2090 4096 2139
rect 3998 2056 4046 2090
rect 4080 2056 4096 2090
rect 3998 2040 4096 2056
rect 22701 1933 22821 1959
rect 22877 1933 22997 1959
rect 23053 1933 23173 1959
rect 23229 1933 23349 1959
rect 3347 1821 3447 1853
rect 3503 1821 3603 1853
rect 22825 1847 22945 1873
rect 23025 1847 23145 1873
rect 23405 1847 23525 1873
rect 23581 1847 23701 1873
rect 3766 1716 3798 1816
rect 3998 1800 4096 1816
rect 3998 1766 4046 1800
rect 4080 1766 4096 1800
rect 3998 1716 4096 1766
rect 4030 1705 4096 1716
rect 4030 1671 4046 1705
rect 4080 1671 4096 1705
rect 4030 1660 4096 1671
rect 3766 1560 3798 1660
rect 3998 1610 4096 1660
rect 3998 1576 4046 1610
rect 4080 1576 4096 1610
rect 3998 1560 4096 1576
rect 22825 1605 22945 1647
rect 23025 1605 23145 1647
rect 22825 1576 23145 1605
rect 3347 1489 3447 1521
rect 3313 1473 3447 1489
rect 3313 1439 3329 1473
rect 3363 1439 3397 1473
rect 3431 1439 3447 1473
rect 3313 1423 3447 1439
rect 3503 1489 3603 1521
rect 22825 1542 22845 1576
rect 22879 1542 22927 1576
rect 22961 1542 23009 1576
rect 23043 1542 23091 1576
rect 23125 1542 23145 1576
rect 22825 1508 23145 1542
rect 23405 1605 23525 1647
rect 23581 1605 23701 1647
rect 23405 1576 23701 1605
rect 23405 1542 23425 1576
rect 23459 1542 23499 1576
rect 23533 1542 23573 1576
rect 23607 1542 23647 1576
rect 23681 1542 23701 1576
rect 23405 1508 23701 1542
rect 3503 1473 3637 1489
rect 22825 1476 22945 1508
rect 23581 1476 23701 1508
rect 3503 1439 3519 1473
rect 3553 1439 3587 1473
rect 3621 1439 3637 1473
rect 3503 1423 3637 1439
rect 3334 1357 3468 1373
rect 3334 1323 3350 1357
rect 3384 1323 3418 1357
rect 3452 1323 3468 1357
rect 3334 1307 3468 1323
rect 3349 1270 3449 1307
rect 22825 1304 22945 1336
rect 23581 1304 23701 1336
rect 3662 1270 3762 1302
rect 3818 1270 3918 1302
rect 3349 1088 3449 1120
rect 3662 1088 3762 1120
rect 3573 1072 3762 1088
rect 3573 1038 3589 1072
rect 3623 1038 3657 1072
rect 3691 1038 3762 1072
rect 3573 1022 3762 1038
rect 3818 1088 3918 1120
rect 3818 1072 3952 1088
rect 3818 1038 3834 1072
rect 3868 1038 3902 1072
rect 3936 1038 3952 1072
rect 3818 1022 3952 1038
rect 3386 786 3418 906
rect 3502 890 3632 906
rect 3502 856 3550 890
rect 3584 856 3632 890
rect 3502 792 3632 856
rect 3502 786 3550 792
rect 3534 758 3550 786
rect 3584 786 3632 792
rect 3716 786 3748 906
rect 3584 758 3600 786
rect 3534 730 3600 758
rect 3386 610 3418 730
rect 3502 694 3632 730
rect 3502 660 3550 694
rect 3584 660 3632 694
rect 3502 610 3632 660
rect 3716 610 3748 730
rect 3848 672 3880 792
rect 3964 776 4062 792
rect 3964 742 4012 776
rect 4046 742 4062 776
rect 3964 699 4062 742
rect 3964 672 4012 699
rect 3996 665 4012 672
rect 4046 665 4062 699
rect 3996 622 4062 665
rect 3996 616 4012 622
rect 3848 496 3880 616
rect 3964 588 4012 616
rect 4046 588 4062 622
rect 3964 545 4062 588
rect 3964 511 4012 545
rect 4046 511 4062 545
rect 3964 496 4062 511
rect 3996 468 4062 496
rect 3996 440 4012 468
rect 3848 320 3880 440
rect 3964 434 4012 440
rect 4046 434 4062 468
rect 3964 392 4062 434
rect 3964 358 4012 392
rect 4046 358 4062 392
rect 3964 320 4062 358
rect 5226 344 5258 464
rect 5458 448 5556 464
rect 5458 414 5506 448
rect 5540 414 5556 448
rect 5458 376 5556 414
rect 5458 344 5506 376
rect 3996 316 4062 320
rect 3996 282 4012 316
rect 4046 282 4062 316
rect 5490 342 5506 344
rect 5540 342 5556 376
rect 5490 304 5556 342
rect 5490 288 5506 304
rect 3996 264 4062 282
rect 3848 144 3880 264
rect 3964 240 4062 264
rect 3964 206 4012 240
rect 4046 206 4062 240
rect 3964 144 4062 206
rect 5226 168 5258 288
rect 5458 270 5506 288
rect 5540 270 5556 304
rect 5458 231 5556 270
rect 5458 197 5506 231
rect 5540 197 5556 231
rect 5458 168 5556 197
rect 6113 448 6211 464
rect 6113 414 6129 448
rect 6163 414 6211 448
rect 6113 372 6211 414
rect 6113 338 6129 372
rect 6163 344 6211 372
rect 6411 344 6443 464
rect 6528 351 6594 367
rect 6163 338 6179 344
rect 6113 295 6179 338
rect 6113 261 6129 295
rect 6163 288 6179 295
rect 6528 317 6544 351
rect 6578 333 6594 351
rect 6578 317 6626 333
rect 6163 261 6211 288
rect 6113 218 6211 261
rect 6113 184 6129 218
rect 6163 184 6211 218
rect 6113 168 6211 184
rect 6411 168 6443 288
rect 6528 283 6626 317
rect 6528 249 6544 283
rect 6578 249 6626 283
rect 6528 233 6626 249
rect 6926 233 6958 333
rect 5490 158 5556 168
rect 5490 124 5506 158
rect 5540 124 5556 158
rect 5490 112 5556 124
rect 5226 -8 5258 112
rect 5458 85 5556 112
rect 5458 51 5506 85
rect 5540 51 5556 85
rect 5458 12 5556 51
rect 5458 -8 5506 12
rect 5490 -22 5506 -8
rect 5540 -22 5556 12
rect 5490 -61 5556 -22
rect 5490 -64 5506 -61
rect 5226 -184 5258 -64
rect 5458 -95 5506 -64
rect 5540 -95 5556 -61
rect 5458 -134 5556 -95
rect 5458 -168 5506 -134
rect 5540 -168 5556 -134
rect 5458 -184 5556 -168
rect 6113 96 6211 112
rect 6113 62 6129 96
rect 6163 62 6211 96
rect 6113 20 6211 62
rect 6113 -14 6129 20
rect 6163 -8 6211 20
rect 6411 -8 6443 112
rect 6528 64 6594 80
rect 6528 30 6544 64
rect 6578 53 6594 64
rect 6578 30 6626 53
rect 6528 -4 6626 30
rect 6163 -14 6179 -8
rect 6113 -57 6179 -14
rect 6113 -91 6129 -57
rect 6163 -64 6179 -57
rect 6528 -38 6544 -4
rect 6578 -38 6626 -4
rect 6528 -47 6626 -38
rect 6926 -47 6958 53
rect 6528 -54 6594 -47
rect 6163 -91 6211 -64
rect 6113 -134 6211 -91
rect 6113 -168 6129 -134
rect 6163 -168 6211 -134
rect 6113 -184 6211 -168
rect 6411 -184 6443 -64
rect 6528 -103 6594 -96
rect 6528 -112 6626 -103
rect 6528 -146 6544 -112
rect 6578 -146 6626 -112
rect 6528 -180 6626 -146
rect 6528 -214 6544 -180
rect 6578 -203 6626 -180
rect 6926 -203 6958 -103
rect 7073 -194 7105 206
rect 7255 159 7385 206
rect 7255 125 7303 159
rect 7337 125 7385 159
rect 7255 84 7385 125
rect 7255 50 7303 84
rect 7337 50 7385 84
rect 7255 8 7385 50
rect 7255 -26 7303 8
rect 7337 -26 7385 8
rect 7255 -68 7385 -26
rect 7255 -102 7303 -68
rect 7337 -102 7385 -68
rect 7255 -144 7385 -102
rect 7255 -178 7303 -144
rect 7337 -178 7385 -144
rect 7255 -194 7385 -178
rect 7535 -194 7567 206
rect 6578 -214 6594 -203
rect 6528 -230 6594 -214
<< polycont >>
rect 4046 2559 4080 2593
rect 4046 2491 4080 2525
rect 4046 2221 4080 2255
rect 4046 2139 4080 2173
rect 22721 2233 22755 2267
rect 22795 2233 22829 2267
rect 22869 2233 22903 2267
rect 22943 2233 22977 2267
rect 23073 2233 23107 2267
rect 23147 2233 23181 2267
rect 23221 2233 23255 2267
rect 23295 2233 23329 2267
rect 4046 2056 4080 2090
rect 4046 1766 4080 1800
rect 4046 1671 4080 1705
rect 4046 1576 4080 1610
rect 3329 1439 3363 1473
rect 3397 1439 3431 1473
rect 22845 1542 22879 1576
rect 22927 1542 22961 1576
rect 23009 1542 23043 1576
rect 23091 1542 23125 1576
rect 23425 1542 23459 1576
rect 23499 1542 23533 1576
rect 23573 1542 23607 1576
rect 23647 1542 23681 1576
rect 3519 1439 3553 1473
rect 3587 1439 3621 1473
rect 3350 1323 3384 1357
rect 3418 1323 3452 1357
rect 3589 1038 3623 1072
rect 3657 1038 3691 1072
rect 3834 1038 3868 1072
rect 3902 1038 3936 1072
rect 3550 856 3584 890
rect 3550 758 3584 792
rect 3550 660 3584 694
rect 4012 742 4046 776
rect 4012 665 4046 699
rect 4012 588 4046 622
rect 4012 511 4046 545
rect 4012 434 4046 468
rect 4012 358 4046 392
rect 5506 414 5540 448
rect 4012 282 4046 316
rect 5506 342 5540 376
rect 4012 206 4046 240
rect 5506 270 5540 304
rect 5506 197 5540 231
rect 6129 414 6163 448
rect 6129 338 6163 372
rect 6129 261 6163 295
rect 6544 317 6578 351
rect 6129 184 6163 218
rect 6544 249 6578 283
rect 5506 124 5540 158
rect 5506 51 5540 85
rect 5506 -22 5540 12
rect 5506 -95 5540 -61
rect 5506 -168 5540 -134
rect 6129 62 6163 96
rect 6129 -14 6163 20
rect 6544 30 6578 64
rect 6129 -91 6163 -57
rect 6544 -38 6578 -4
rect 6129 -168 6163 -134
rect 6544 -146 6578 -112
rect 6544 -214 6578 -180
rect 7303 125 7337 159
rect 7303 50 7337 84
rect 7303 -26 7337 8
rect 7303 -102 7337 -68
rect 7303 -178 7337 -144
<< locali >>
rect 18040 2832 23412 2927
rect 17530 2797 17797 2832
rect 17935 2797 20701 2832
rect 20851 2797 23412 2832
rect 2722 2654 2760 2688
rect 3612 2687 4002 2688
rect 3612 2653 3641 2687
rect 3675 2653 4002 2687
rect 3612 2620 4002 2653
rect 3612 2615 3816 2620
rect 3612 2581 3641 2615
rect 3675 2586 3816 2615
rect 3850 2586 3884 2620
rect 3918 2586 3952 2620
rect 3986 2586 4002 2620
rect 21281 2660 23412 2797
rect 21281 2614 24132 2660
rect 3675 2581 4002 2586
rect 4046 2596 4080 2609
rect 4046 2525 4080 2559
rect 22676 2558 24132 2614
rect 3450 2464 4002 2499
rect 4046 2475 4080 2490
rect 3450 2430 3816 2464
rect 3850 2430 3884 2464
rect 3918 2430 3952 2464
rect 3986 2430 4002 2464
rect 3450 2429 4002 2430
rect 22832 2459 22866 2475
rect 2695 1147 2816 2356
rect 3302 1937 3409 1949
rect 3302 1903 3369 1937
rect 3403 1903 3409 1937
rect 3302 1865 3409 1903
rect 3302 1831 3369 1865
rect 3403 1831 3409 1865
rect 3302 1771 3409 1831
rect 3336 1737 3409 1771
rect 3302 1703 3409 1737
rect 3336 1669 3409 1703
rect 3302 1635 3409 1669
rect 3336 1601 3409 1635
rect 3302 1567 3409 1601
rect 3336 1533 3409 1567
rect 3302 1473 3409 1533
rect 3450 1775 3563 2429
rect 22832 2391 22866 2413
rect 3450 1737 3458 1775
rect 3492 1737 3563 1775
rect 3450 1703 3563 1737
rect 3450 1637 3458 1703
rect 3492 1637 3563 1703
rect 3450 1635 3563 1637
rect 3450 1601 3458 1635
rect 3492 1601 3563 1635
rect 3450 1567 3563 1601
rect 3450 1533 3458 1567
rect 3492 1533 3563 1567
rect 3450 1526 3563 1533
rect 3613 2356 3711 2369
rect 3613 2322 3643 2356
rect 3677 2322 3711 2356
rect 3613 2284 3711 2322
rect 3800 2341 4159 2372
rect 23008 2459 23042 2558
rect 23360 2475 23394 2558
rect 23008 2391 23042 2425
rect 23008 2341 23042 2357
rect 23184 2459 23218 2475
rect 23184 2391 23218 2413
rect 23968 2463 24132 2558
rect 23968 2429 24006 2463
rect 24040 2429 24132 2463
rect 23968 2393 24132 2429
rect 23968 2359 24006 2393
rect 24040 2359 24132 2393
rect 3800 2307 3816 2341
rect 3850 2307 3884 2341
rect 3918 2307 3952 2341
rect 3986 2333 4159 2341
rect 3986 2317 4125 2333
rect 3986 2307 4002 2317
rect 3613 2250 3643 2284
rect 3677 2261 3711 2284
rect 3677 2250 4002 2261
rect 3613 2185 4002 2250
rect 3613 2151 3816 2185
rect 3850 2151 3884 2185
rect 3918 2151 3952 2185
rect 3986 2151 4002 2185
rect 3613 2080 4002 2151
rect 4125 2261 4159 2299
rect 23968 2323 24132 2359
rect 23968 2289 24006 2323
rect 24040 2289 24132 2323
rect 22705 2233 22721 2267
rect 22755 2233 22795 2267
rect 22829 2233 22869 2267
rect 22903 2233 22909 2267
rect 22977 2233 22993 2267
rect 23057 2233 23073 2267
rect 23107 2255 23147 2267
rect 23127 2233 23147 2255
rect 23181 2233 23221 2267
rect 23255 2233 23295 2267
rect 23329 2233 23345 2267
rect 23968 2253 24132 2289
rect 4046 2184 4080 2221
rect 20194 2192 20222 2221
rect 20194 2169 20256 2192
rect 22909 2195 22943 2233
rect 4046 2090 4080 2139
rect 3613 1937 3711 2080
rect 4046 2040 4080 2052
rect 3800 1995 3816 2029
rect 3850 1995 3860 2029
rect 3918 1995 3932 2029
rect 3986 1995 4002 2029
rect 5321 2009 5367 2015
rect 5401 2009 5446 2015
rect 5480 2009 5525 2015
rect 5559 2009 5604 2015
rect 5638 2009 5683 2015
rect 5717 2009 5762 2015
rect 5796 2009 5841 2015
rect 5875 2009 5920 2015
rect 5954 2009 5999 2015
rect 6895 2009 6954 2163
rect 20194 2154 20328 2169
rect 20194 2120 20222 2154
rect 20256 2120 20328 2154
rect 20194 2053 20328 2120
rect 22656 2141 22690 2157
rect 22656 2073 22690 2107
rect 5257 1975 5287 2009
rect 5321 1975 5356 2009
rect 5401 1981 5425 2009
rect 5480 1981 5494 2009
rect 5559 1981 5563 2009
rect 5390 1975 5425 1981
rect 5459 1975 5494 1981
rect 5528 1975 5563 1981
rect 5597 1981 5604 2009
rect 5666 1981 5683 2009
rect 5735 1981 5762 2009
rect 5597 1975 5632 1981
rect 5666 1975 5701 1981
rect 5735 1975 5770 1981
rect 5804 1975 5839 2009
rect 5875 1981 5908 2009
rect 5954 1981 5977 2009
rect 6033 1981 6046 2009
rect 5873 1975 5908 1981
rect 5942 1975 5977 1981
rect 6011 1975 6046 1981
rect 6080 1975 6115 2009
rect 6149 1975 6184 2009
rect 6218 1975 6253 2009
rect 6287 1975 6322 2009
rect 6356 1975 6391 2009
rect 6425 1975 6460 2009
rect 6494 1975 6529 2009
rect 6563 1975 6598 2009
rect 6632 1975 6667 2009
rect 6701 1975 6736 2009
rect 6770 1975 6805 2009
rect 6839 1975 6874 2009
rect 6908 1975 6943 2009
rect 6977 1975 7012 2009
rect 7046 1975 7081 2009
rect 7115 1975 7150 2009
rect 7184 1975 7208 2009
rect 5257 1948 7208 1975
rect 22656 2006 22690 2039
rect 3613 1903 3643 1937
rect 3677 1903 3711 1937
rect 3613 1865 3711 1903
rect 22656 1934 22690 1971
rect 23093 2183 23127 2221
rect 22832 2098 22866 2107
rect 22832 2005 22866 2039
rect 22832 1955 22866 1971
rect 23008 2141 23042 2157
rect 23968 2219 24006 2253
rect 24040 2219 24132 2253
rect 23968 2183 24132 2219
rect 23008 2073 23042 2107
rect 23008 2006 23042 2039
rect 23008 1934 23042 1971
rect 23360 2156 23394 2157
rect 23184 2097 23218 2107
rect 23184 2005 23218 2039
rect 23184 1955 23218 1971
rect 23284 2141 23394 2156
rect 23284 2107 23360 2141
rect 23284 2073 23394 2107
rect 23284 2039 23360 2073
rect 23284 2006 23394 2039
rect 23968 2149 24006 2183
rect 24040 2149 24132 2183
rect 23968 2112 24132 2149
rect 23968 2078 24006 2112
rect 24040 2078 24132 2112
rect 23968 2041 24132 2078
rect 23968 2007 24006 2041
rect 24040 2007 24132 2041
rect 23284 1971 23360 2006
rect 23284 1926 23394 1971
rect 23284 1892 23360 1926
rect 3613 1831 3643 1865
rect 3677 1831 3711 1865
rect 3613 1771 3711 1831
rect 3794 1857 3810 1861
rect 3794 1827 3801 1857
rect 3844 1827 3878 1861
rect 3912 1827 3946 1861
rect 3980 1827 3996 1861
rect 22780 1829 22814 1852
rect 23284 1846 23394 1892
rect 3613 1737 3614 1771
rect 3648 1737 3711 1771
rect 3801 1785 3835 1823
rect 4046 1800 4080 1816
rect 3613 1705 3711 1737
rect 4046 1705 4080 1766
rect 3613 1703 3810 1705
rect 3613 1669 3614 1703
rect 3648 1671 3810 1703
rect 3844 1671 3878 1705
rect 3912 1671 3946 1705
rect 3980 1671 3996 1705
rect 3648 1669 3996 1671
rect 3613 1635 3996 1669
rect 3613 1601 3614 1635
rect 3648 1618 3996 1635
rect 3648 1601 3711 1618
rect 3613 1567 3711 1601
rect 3613 1533 3614 1567
rect 3648 1533 3711 1567
rect 4046 1610 4080 1666
rect 22780 1761 22814 1780
rect 22968 1829 23002 1845
rect 22968 1761 23002 1795
rect 22780 1693 22814 1727
rect 22990 1716 23002 1727
rect 22956 1693 23002 1716
rect 18645 1605 19234 1653
rect 22780 1643 22814 1659
rect 22854 1672 22916 1684
rect 22163 1576 22197 1614
rect 22854 1638 22865 1672
rect 22899 1638 22916 1672
rect 22956 1678 22968 1693
rect 22990 1644 23002 1659
rect 22968 1643 23002 1644
rect 23190 1795 23258 1846
rect 23292 1795 23360 1846
rect 23712 1933 23746 1972
rect 23712 1860 23746 1899
rect 23156 1774 23394 1795
rect 23190 1727 23258 1774
rect 23292 1727 23360 1774
rect 23156 1702 23394 1727
rect 23190 1659 23258 1702
rect 23292 1659 23360 1702
rect 23156 1643 23394 1659
rect 23536 1829 23570 1845
rect 23536 1761 23570 1795
rect 23536 1693 23570 1716
rect 23536 1643 23570 1644
rect 23968 1970 24132 2007
rect 23968 1936 24006 1970
rect 24040 1936 24132 1970
rect 23968 1899 24132 1936
rect 23968 1865 24006 1899
rect 24040 1865 24132 1899
rect 23968 1828 24132 1865
rect 23968 1804 24006 1828
rect 23712 1761 23746 1795
rect 23712 1693 23746 1727
rect 23712 1643 23746 1659
rect 23961 1794 24006 1804
rect 24040 1794 24132 1828
rect 22854 1600 22916 1638
rect 22854 1576 22865 1600
rect 22899 1576 22916 1600
rect 4046 1560 4080 1572
rect 3458 1517 3492 1526
rect 3613 1517 3711 1533
rect 3794 1515 3810 1549
rect 3844 1515 3878 1549
rect 3912 1526 3946 1549
rect 3980 1526 3996 1549
rect 21742 1542 21780 1576
rect 22829 1542 22845 1576
rect 22899 1566 22927 1576
rect 22879 1542 22927 1566
rect 22961 1542 23009 1576
rect 23043 1542 23091 1576
rect 23125 1542 23141 1576
rect 23392 1542 23425 1576
rect 23464 1542 23499 1576
rect 23533 1542 23573 1576
rect 23607 1542 23647 1576
rect 23681 1542 23697 1576
rect 3924 1515 3946 1526
rect 3794 1492 3890 1515
rect 3924 1492 3962 1515
rect 3794 1491 3996 1492
rect 3302 1440 3329 1473
rect 3313 1439 3329 1440
rect 3363 1439 3397 1473
rect 3431 1439 3447 1473
rect 3503 1439 3515 1473
rect 3553 1439 3587 1473
rect 3625 1439 3637 1473
rect 22780 1450 22814 1466
rect 3506 1372 3951 1397
rect 3334 1323 3346 1357
rect 3384 1323 3418 1357
rect 3456 1323 3468 1357
rect 3506 1338 3843 1372
rect 3877 1338 3915 1372
rect 3949 1338 3951 1372
rect 3506 1321 3951 1338
rect 22780 1382 22814 1404
rect 22956 1394 22990 1416
rect 22956 1332 22990 1348
rect 23712 1450 23746 1466
rect 23536 1394 23570 1416
rect 23536 1332 23570 1348
rect 23726 1404 23746 1416
rect 23692 1382 23746 1404
rect 23692 1366 23712 1382
rect 23726 1332 23746 1348
rect 3506 1297 3574 1321
rect 3491 1250 3574 1297
rect 3244 1234 3338 1250
rect 3244 1200 3304 1234
rect 3244 1166 3338 1200
rect 3244 1132 3304 1166
rect 3244 1004 3338 1132
rect 3460 1234 3574 1250
rect 3494 1200 3574 1234
rect 3460 1166 3574 1200
rect 3494 1132 3574 1166
rect 3617 1258 3651 1274
rect 3763 1258 3807 1274
rect 3617 1221 3618 1224
rect 3652 1221 3690 1255
rect 3763 1224 3773 1258
rect 3617 1190 3651 1221
rect 3763 1190 3807 1224
rect 3763 1185 3773 1190
rect 3617 1140 3651 1156
rect 3742 1156 3773 1185
rect 3742 1140 3807 1156
rect 3929 1258 3963 1274
rect 22654 1239 23309 1242
rect 3929 1213 3930 1224
rect 3929 1190 3964 1213
rect 3963 1175 3964 1190
rect 3929 1141 3930 1156
rect 22627 1238 23844 1239
rect 23961 1238 24132 1794
rect 22627 1236 24132 1238
rect 22627 1205 22686 1236
rect 22720 1205 22766 1236
rect 22627 1171 22661 1205
rect 22720 1202 22731 1205
rect 22695 1171 22731 1202
rect 22765 1202 22766 1205
rect 22800 1205 22846 1236
rect 22880 1205 22926 1236
rect 22960 1205 23006 1236
rect 23040 1205 23085 1236
rect 23119 1205 23164 1236
rect 23198 1205 23243 1236
rect 23277 1205 23321 1236
rect 23355 1205 23400 1236
rect 23434 1205 23479 1236
rect 23513 1205 23558 1236
rect 23592 1205 23637 1236
rect 23671 1205 23716 1236
rect 23750 1205 23795 1236
rect 22800 1202 22801 1205
rect 22765 1171 22801 1202
rect 22835 1202 22846 1205
rect 22905 1202 22926 1205
rect 22975 1202 23006 1205
rect 22835 1171 22871 1202
rect 22905 1171 22941 1202
rect 22975 1171 23011 1202
rect 23045 1171 23081 1205
rect 23119 1202 23151 1205
rect 23198 1202 23221 1205
rect 23277 1202 23291 1205
rect 23355 1202 23361 1205
rect 23115 1171 23151 1202
rect 23185 1171 23221 1202
rect 23255 1171 23291 1202
rect 23325 1171 23361 1202
rect 23395 1202 23400 1205
rect 23465 1202 23479 1205
rect 23534 1202 23558 1205
rect 23603 1202 23637 1205
rect 23395 1171 23431 1202
rect 23465 1171 23500 1202
rect 23534 1171 23569 1202
rect 23603 1171 23638 1202
rect 23672 1171 23707 1205
rect 23750 1202 23776 1205
rect 23829 1202 24132 1236
rect 23741 1171 23776 1202
rect 23810 1171 24132 1202
rect 22627 1164 24132 1171
rect 22627 1151 22686 1164
rect 3929 1140 3963 1141
rect 3460 1116 3574 1132
rect 3623 1038 3645 1072
rect 3691 1038 3707 1072
rect 2816 1002 3480 1004
rect 3742 1002 3783 1140
rect 22421 1117 22455 1151
rect 22489 1117 22559 1151
rect 22593 1137 22686 1151
rect 22720 1137 22766 1164
rect 22593 1117 22661 1137
rect 22720 1130 22731 1137
rect 4125 1084 4159 1116
rect 3818 1078 4159 1084
rect 3818 1072 4125 1078
rect 3818 1038 3834 1072
rect 3868 1038 3902 1072
rect 3936 1044 4125 1072
rect 3936 1038 4159 1044
rect 21851 1103 22661 1117
rect 22695 1103 22731 1130
rect 22765 1130 22766 1137
rect 22800 1137 22846 1164
rect 22880 1137 22926 1164
rect 22960 1137 23006 1164
rect 23040 1137 23085 1164
rect 23119 1137 23164 1164
rect 23198 1137 23243 1164
rect 23277 1137 24132 1164
rect 22800 1130 22801 1137
rect 22765 1103 22801 1130
rect 22835 1130 22846 1137
rect 22905 1130 22926 1137
rect 22975 1130 23006 1137
rect 22835 1103 22871 1130
rect 22905 1103 22941 1130
rect 22975 1103 23011 1130
rect 23045 1103 23081 1137
rect 23119 1130 23151 1137
rect 23198 1130 23221 1137
rect 23277 1130 23291 1137
rect 23115 1103 23151 1130
rect 23185 1103 23221 1130
rect 23255 1103 23291 1130
rect 23325 1124 23361 1137
rect 23355 1103 23361 1124
rect 23395 1124 23431 1137
rect 23465 1124 23500 1137
rect 23534 1124 23569 1137
rect 23603 1124 23638 1137
rect 23395 1103 23400 1124
rect 23465 1103 23479 1124
rect 23534 1103 23558 1124
rect 23603 1103 23637 1124
rect 23672 1103 23707 1137
rect 23741 1124 23776 1137
rect 23810 1124 24132 1137
rect 23750 1103 23776 1124
rect 21851 1092 23321 1103
rect 21851 1083 22686 1092
rect 21851 1049 21853 1083
rect 21887 1049 21929 1083
rect 21963 1049 22005 1083
rect 22039 1049 22081 1083
rect 22115 1049 22157 1083
rect 22191 1049 22233 1083
rect 22267 1049 22309 1083
rect 22343 1049 22385 1083
rect 22419 1069 22686 1083
rect 22720 1069 22766 1092
rect 22419 1067 22661 1069
rect 22419 1049 22455 1067
rect 2816 951 3783 1002
rect 2816 917 3430 951
rect 3464 942 3644 951
rect 3464 917 3480 942
rect 3628 917 3644 942
rect 3678 942 3783 951
rect 3678 917 3694 942
rect 3742 941 3783 942
rect 21851 1033 22455 1049
rect 22489 1033 22559 1067
rect 22593 1035 22661 1067
rect 22720 1058 22731 1069
rect 22695 1035 22731 1058
rect 22765 1058 22766 1069
rect 22800 1069 22846 1092
rect 22880 1069 22926 1092
rect 22960 1069 23006 1092
rect 23040 1069 23085 1092
rect 23119 1069 23164 1092
rect 23198 1069 23243 1092
rect 23277 1090 23321 1092
rect 23355 1090 23400 1103
rect 23434 1090 23479 1103
rect 23513 1090 23558 1103
rect 23592 1090 23637 1103
rect 23671 1090 23716 1103
rect 23750 1090 23795 1103
rect 23829 1090 24132 1124
rect 23277 1069 24132 1090
rect 22800 1058 22801 1069
rect 22765 1035 22801 1058
rect 22835 1058 22846 1069
rect 22905 1058 22926 1069
rect 22975 1058 23006 1069
rect 22835 1035 22871 1058
rect 22905 1035 22941 1058
rect 22975 1035 23011 1058
rect 23045 1035 23081 1069
rect 23119 1058 23151 1069
rect 23198 1058 23221 1069
rect 23277 1058 23291 1069
rect 23115 1035 23151 1058
rect 23185 1035 23221 1058
rect 23255 1035 23291 1058
rect 23325 1035 23361 1069
rect 23395 1035 23431 1069
rect 23465 1035 23500 1069
rect 23534 1035 23569 1069
rect 23603 1035 23638 1069
rect 23672 1035 23707 1069
rect 23741 1035 23776 1069
rect 23810 1035 24132 1069
rect 22593 1033 24132 1035
rect 21851 1020 24132 1033
rect 21851 1011 22686 1020
rect 21851 977 21853 1011
rect 21887 977 21929 1011
rect 21963 977 22005 1011
rect 22039 977 22081 1011
rect 22115 977 22157 1011
rect 22191 977 22233 1011
rect 22267 977 22309 1011
rect 22343 977 22385 1011
rect 22419 1001 22686 1011
rect 22720 1001 22766 1020
rect 22419 983 22661 1001
rect 22720 986 22731 1001
rect 22419 977 22455 983
rect 21851 949 22455 977
rect 22489 949 22559 983
rect 22593 967 22661 983
rect 22695 967 22731 986
rect 22765 986 22766 1001
rect 22800 1001 22846 1020
rect 22880 1001 22926 1020
rect 22960 1001 23006 1020
rect 23040 1001 23085 1020
rect 23119 1001 23164 1020
rect 23198 1001 23243 1020
rect 23277 1001 24132 1020
rect 22800 986 22801 1001
rect 22765 967 22801 986
rect 22835 986 22846 1001
rect 22905 986 22926 1001
rect 22975 986 23006 1001
rect 22835 967 22871 986
rect 22905 967 22941 986
rect 22975 967 23011 986
rect 23045 967 23081 1001
rect 23119 986 23151 1001
rect 23198 986 23221 1001
rect 23277 986 23291 1001
rect 23115 967 23151 986
rect 23185 967 23221 986
rect 23255 967 23291 986
rect 23325 967 23361 1001
rect 23395 967 23431 1001
rect 23465 967 23500 1001
rect 23534 967 23569 1001
rect 23603 967 23638 1001
rect 23672 967 23707 1001
rect 23741 967 23776 1001
rect 23810 967 24132 1001
rect 22593 949 24132 967
rect 21851 938 24132 949
rect 2816 914 3480 917
rect 3550 894 3584 906
rect 3461 775 3495 793
rect 3414 741 3430 775
rect 3464 755 3495 775
rect 3550 792 3584 856
rect 21851 904 21853 938
rect 21887 904 21929 938
rect 21963 904 22005 938
rect 22039 904 22081 938
rect 22115 904 22157 938
rect 22191 904 22233 938
rect 22267 904 22309 938
rect 22343 904 22385 938
rect 22419 933 24132 938
rect 22419 904 22661 933
rect 21851 899 22661 904
rect 22695 899 22731 933
rect 22765 899 22801 933
rect 22835 899 22871 933
rect 22905 899 22941 933
rect 22975 899 23011 933
rect 23045 899 23081 933
rect 23115 899 23151 933
rect 23185 899 23221 933
rect 23255 899 23291 933
rect 23325 899 23361 933
rect 23395 899 23431 933
rect 23465 899 23500 933
rect 23534 899 23569 933
rect 23603 899 23638 933
rect 23672 899 23707 933
rect 23741 899 23776 933
rect 23810 899 24132 933
rect 21851 865 22455 899
rect 22489 865 22559 899
rect 22593 869 24132 899
rect 22593 865 23844 869
rect 3780 803 3892 837
rect 3926 803 3943 837
rect 3550 694 3584 758
rect 3628 748 3644 775
rect 3678 748 3694 775
rect 3780 764 3943 803
rect 4012 776 4046 792
rect 3628 741 3640 748
rect 3678 741 3712 748
rect 3674 714 3712 741
rect 3550 644 3584 656
rect 3780 599 3824 764
rect 4045 711 4046 742
rect 4011 699 4046 711
rect 4011 665 4012 699
rect 3926 627 3930 661
rect 4011 659 4046 665
rect 3411 565 3430 599
rect 3464 565 3644 599
rect 3678 565 3824 599
rect 3411 521 3824 565
rect 3459 508 3824 521
rect 4045 625 4046 659
rect 4011 622 4046 625
rect 4011 588 4012 622
rect 4011 573 4046 588
rect 4045 545 4046 573
rect 4011 511 4012 539
rect 3459 485 3943 508
rect 3459 451 3892 485
rect 3926 451 3943 485
rect 3459 435 3943 451
rect 4011 486 4046 511
rect 4045 468 4046 486
rect 3459 407 3815 435
rect 3763 145 3815 407
rect 4011 434 4012 452
rect 4011 399 4046 434
rect 4045 392 4046 399
rect 4012 316 4046 358
rect 3926 275 3930 309
rect 4012 240 4046 282
rect 4012 190 4046 206
rect 3457 135 3815 145
rect 4106 135 4174 837
rect 21851 831 21853 865
rect 21887 831 21929 865
rect 21963 831 22005 865
rect 22039 831 22081 865
rect 22115 831 22157 865
rect 22191 831 22233 865
rect 22267 831 22309 865
rect 22343 831 22385 865
rect 22419 831 22421 865
rect 21851 792 22421 831
rect 21851 758 21853 792
rect 21887 758 21929 792
rect 21963 758 22005 792
rect 22039 758 22081 792
rect 22115 758 22157 792
rect 22191 758 22233 792
rect 22267 758 22309 792
rect 22343 758 22385 792
rect 22419 758 22421 792
rect 21851 739 22421 758
rect 21615 719 22421 739
rect 21615 685 21853 719
rect 21887 685 21929 719
rect 21963 685 22005 719
rect 22039 685 22081 719
rect 22115 685 22157 719
rect 22191 685 22233 719
rect 22267 685 22309 719
rect 22343 685 22385 719
rect 22419 685 22421 719
rect 21615 646 22421 685
rect 21615 612 21853 646
rect 21887 612 21929 646
rect 21963 612 22005 646
rect 22039 612 22081 646
rect 22115 612 22157 646
rect 22191 612 22233 646
rect 22267 612 22309 646
rect 22343 612 22385 646
rect 22419 612 22421 646
rect 7542 570 8014 582
rect 5145 526 5456 539
rect 5145 492 5151 526
rect 5185 509 5456 526
rect 7542 536 7547 570
rect 7581 536 8014 570
rect 5185 492 5270 509
rect 5145 475 5270 492
rect 5304 475 5338 509
rect 5372 475 5406 509
rect 5440 475 5456 509
rect 6213 475 6229 509
rect 6263 475 6297 509
rect 6331 475 6365 509
rect 6420 478 6458 512
rect 6529 478 6553 512
rect 6587 478 6628 512
rect 6662 478 6703 512
rect 6737 478 6772 512
rect 6812 478 6853 512
rect 6890 478 6927 512
rect 6973 478 6985 512
rect 7542 499 8014 536
rect 7542 498 7712 499
rect 6399 475 6415 478
rect 5145 454 5456 475
rect 7542 473 7547 498
rect 7581 473 7712 498
rect 7940 473 8014 499
rect 15914 508 15948 546
rect 21615 573 22421 612
rect 5145 446 5151 454
rect 5185 446 5456 454
rect 5506 452 5540 464
rect 6129 452 6163 464
rect 6153 448 6163 452
rect 5506 376 5540 414
rect 5254 333 5456 369
rect 5254 299 5270 333
rect 5304 299 5338 333
rect 5372 309 5406 333
rect 5440 309 5456 333
rect 5373 299 5406 309
rect 5254 275 5339 299
rect 5373 275 5411 299
rect 5445 275 5456 309
rect 5254 263 5456 275
rect 5506 304 5540 341
rect 5506 231 5540 263
rect 3457 133 4174 135
rect 3457 99 3892 133
rect 3926 99 4174 133
rect 3457 33 4174 99
rect 5145 163 5151 188
rect 5185 163 5456 188
rect 5145 157 5456 163
rect 5145 125 5270 157
rect 5145 95 5151 125
rect 5185 123 5270 125
rect 5304 123 5338 157
rect 5372 123 5406 157
rect 5440 123 5456 157
rect 5185 95 5456 123
rect 5506 158 5540 185
rect 5764 283 5823 431
rect 16001 439 16035 477
rect 6119 414 6129 418
rect 6119 379 6163 414
rect 16171 409 16205 447
rect 6153 372 6163 379
rect 6119 338 6129 345
rect 6119 306 6163 338
rect 6153 295 6163 306
rect 5764 249 5792 283
rect 5764 211 5826 249
rect 5764 177 5792 211
rect 6119 261 6129 272
rect 6213 347 6293 369
rect 6327 347 6415 369
rect 6213 333 6415 347
rect 6213 299 6229 333
rect 6263 309 6297 333
rect 6263 299 6293 309
rect 6331 299 6365 333
rect 6399 299 6415 333
rect 6213 275 6293 299
rect 6327 275 6415 299
rect 6213 263 6415 275
rect 6544 355 6578 367
rect 6622 344 6634 378
rect 6672 344 6706 378
rect 6740 344 6774 378
rect 6808 344 6842 378
rect 6876 344 6892 378
rect 7294 367 7328 405
rect 16970 508 17004 546
rect 16266 439 16300 477
rect 16525 409 16559 447
rect 16618 409 16652 447
rect 17479 497 17513 535
rect 21615 539 21853 573
rect 21887 539 21929 573
rect 21963 539 22005 573
rect 22039 539 22081 573
rect 22115 539 22157 573
rect 22191 539 22233 573
rect 22267 539 22309 573
rect 22343 539 22385 573
rect 22419 539 22421 573
rect 21615 500 22421 539
rect 21615 466 21853 500
rect 21887 466 21929 500
rect 21963 466 22005 500
rect 22039 466 22081 500
rect 22115 466 22157 500
rect 22191 466 22233 500
rect 22267 466 22309 500
rect 22343 466 22385 500
rect 22419 466 22421 500
rect 16883 409 16917 447
rect 21615 427 22421 466
rect 21615 393 21853 427
rect 21887 393 21929 427
rect 21963 393 22005 427
rect 22039 393 22081 427
rect 22115 393 22157 427
rect 22191 393 22233 427
rect 22267 393 22309 427
rect 22343 393 22385 427
rect 22419 393 22421 427
rect 6544 283 6578 317
rect 6119 232 6163 261
rect 6544 233 6578 249
rect 7101 251 7515 294
rect 6153 218 6163 232
rect 6119 184 6129 198
rect 6622 188 6638 222
rect 6672 188 6706 222
rect 6740 188 6774 222
rect 6808 188 6842 222
rect 6891 188 6929 222
rect 7101 217 7117 251
rect 7151 217 7185 251
rect 7219 217 7397 251
rect 7431 217 7465 251
rect 7499 217 7515 251
rect 18541 247 19184 392
rect 21615 354 22421 393
rect 21615 320 21853 354
rect 21887 320 21929 354
rect 21963 320 22005 354
rect 22039 320 22081 354
rect 22115 320 22157 354
rect 22191 320 22233 354
rect 22267 320 22309 354
rect 22343 320 22385 354
rect 22419 320 22421 354
rect 21615 281 22421 320
rect 21615 247 21853 281
rect 21887 247 21929 281
rect 21963 247 22005 281
rect 22039 247 22081 281
rect 22115 247 22157 281
rect 22191 247 22233 281
rect 22267 247 22309 281
rect 22343 247 22385 281
rect 22419 247 22421 281
rect 7101 216 7515 217
rect 3457 -1 3773 33
rect 3807 -1 4174 33
rect 3457 -39 4174 -1
rect 5506 85 5540 107
rect 6119 168 6163 184
rect 6119 158 6153 168
rect 6119 112 6153 124
rect 6213 123 6229 157
rect 6263 123 6297 157
rect 6331 123 6365 157
rect 6420 123 6458 157
rect 7101 135 7269 216
rect 18583 189 18628 223
rect 18662 189 18707 223
rect 18741 189 18786 223
rect 18820 189 18865 223
rect 18899 189 18944 223
rect 18978 189 19023 223
rect 19057 189 19101 223
rect 21615 213 22421 247
rect 6119 96 6163 112
rect 7101 101 7113 135
rect 7147 101 7185 135
rect 7219 101 7269 135
rect 6119 84 6129 96
rect 6153 50 6163 62
rect 5506 12 5540 29
rect 3457 -73 3773 -39
rect 3807 -73 4174 -39
rect 5254 -53 5265 -19
rect 5304 -53 5337 -19
rect 5372 -53 5406 -19
rect 5440 -53 5456 -19
rect 3457 -86 4174 -73
rect 5506 -61 5540 -49
rect 5506 -134 5540 -127
rect 5506 -184 5540 -168
rect 5254 -229 5266 -195
rect 5304 -229 5338 -195
rect 5372 -229 5406 -195
rect 5444 -229 5456 -195
rect 5805 -203 5851 37
rect 6119 20 6163 50
rect 6119 10 6129 20
rect 6288 72 6578 80
rect 6288 38 6299 72
rect 6333 38 6371 72
rect 6405 64 6578 72
rect 6622 64 6634 98
rect 6672 64 6706 98
rect 6740 64 6774 98
rect 6808 64 6842 98
rect 6876 64 6892 98
rect 6405 38 6544 64
rect 6288 30 6544 38
rect 6288 17 6578 30
rect 6977 21 7011 47
rect 6153 -24 6163 -14
rect 6544 -4 6578 17
rect 6119 -57 6163 -24
rect 6213 -53 6225 -19
rect 6263 -53 6297 -19
rect 6331 -53 6365 -19
rect 6399 -53 6415 -19
rect 6544 -54 6578 -38
rect 6622 9 7040 21
rect 6622 -25 6977 9
rect 7011 -25 7040 9
rect 6622 -37 7040 -25
rect 6119 -64 6129 -57
rect 6153 -98 6163 -91
rect 6622 -58 6936 -37
rect 6622 -92 6638 -58
rect 6672 -92 6706 -58
rect 6740 -92 6774 -58
rect 6808 -92 6842 -58
rect 6876 -92 6936 -58
rect 7101 -90 7269 101
rect 6119 -134 6163 -98
rect 6119 -138 6129 -134
rect 6153 -172 6163 -168
rect 6129 -184 6163 -172
rect 6544 -112 6578 -96
rect 6987 -126 7269 -90
rect 6578 -146 7269 -126
rect 6544 -159 7269 -146
rect 7303 163 7337 175
rect 7303 86 7337 125
rect 18549 115 19135 189
rect 18583 81 18628 115
rect 18662 81 18707 115
rect 18741 81 18786 115
rect 18820 81 18865 115
rect 18899 81 18944 115
rect 18978 81 19023 115
rect 19057 81 19101 115
rect 7303 8 7337 50
rect 7303 -68 7337 -26
rect 7303 -144 7337 -104
rect 7381 -57 7911 -26
rect 7381 -91 7393 -57
rect 7427 -91 7472 -57
rect 7506 -91 7911 -57
rect 7381 -122 7911 -91
rect 6544 -180 7068 -159
rect 5584 -237 5601 -203
rect 5642 -237 5680 -203
rect 5717 -237 5758 -203
rect 5793 -237 5833 -203
rect 5872 -237 5908 -203
rect 5950 -237 5982 -203
rect 6028 -237 6040 -203
rect 6213 -229 6225 -195
rect 6263 -229 6297 -195
rect 6331 -229 6365 -195
rect 6403 -229 6415 -195
rect 7303 -194 7337 -182
rect 15865 -197 15877 -163
rect 15923 -197 15953 -163
rect 15993 -197 16029 -163
rect 16063 -197 16098 -163
rect 16139 -197 16167 -163
rect 16215 -197 16236 -163
rect 16291 -197 16305 -163
rect 16366 -197 16374 -163
rect 16441 -197 16443 -163
rect 16477 -197 16482 -163
rect 16546 -197 16557 -163
rect 16615 -197 16632 -163
rect 16684 -197 16707 -163
rect 16753 -197 16782 -163
rect 16822 -197 16857 -163
rect 16891 -197 16926 -163
rect 16966 -197 16995 -163
rect 17041 -197 17053 -163
rect 7101 -214 7117 -205
rect 6544 -230 6578 -214
rect 6622 -248 6638 -214
rect 6672 -248 6706 -214
rect 6740 -248 6774 -214
rect 6834 -248 6842 -214
rect 7101 -239 7113 -214
rect 7151 -239 7185 -205
rect 7219 -239 7235 -205
rect 7381 -214 7397 -205
rect 7381 -239 7393 -214
rect 7431 -239 7465 -205
rect 7499 -239 7515 -205
rect 7147 -248 7185 -239
rect 7427 -248 7465 -239
<< viali >>
rect 2688 2654 2722 2688
rect 2760 2654 2794 2688
rect 3641 2653 3675 2687
rect 3641 2581 3675 2615
rect 4046 2593 4080 2596
rect 4046 2562 4080 2593
rect 4046 2491 4080 2524
rect 4046 2490 4080 2491
rect 3369 1903 3403 1937
rect 3369 1831 3403 1865
rect 22832 2425 22866 2447
rect 22832 2413 22866 2425
rect 3458 1771 3492 1775
rect 3458 1741 3492 1771
rect 3458 1669 3492 1671
rect 3458 1637 3492 1669
rect 3458 1533 3492 1567
rect 3643 2322 3677 2356
rect 22832 2357 22866 2375
rect 22832 2341 22866 2357
rect 23184 2425 23218 2447
rect 23184 2413 23218 2425
rect 23184 2357 23218 2375
rect 23184 2341 23218 2357
rect 3643 2250 3677 2284
rect 4125 2299 4159 2333
rect 4046 2255 4080 2281
rect 4046 2247 4080 2255
rect 4125 2227 4159 2261
rect 22909 2233 22943 2267
rect 23093 2233 23107 2255
rect 23107 2233 23127 2255
rect 4046 2173 4080 2184
rect 4046 2150 4080 2173
rect 20222 2192 20256 2226
rect 4046 2056 4080 2086
rect 4046 2052 4080 2056
rect 3860 1995 3884 2029
rect 3884 1995 3894 2029
rect 3932 1995 3952 2029
rect 3952 1995 3966 2029
rect 5287 2009 5321 2015
rect 5367 2009 5401 2015
rect 5446 2009 5480 2015
rect 5525 2009 5559 2015
rect 5604 2009 5638 2015
rect 5683 2009 5717 2015
rect 5762 2009 5796 2015
rect 5841 2009 5875 2015
rect 5920 2009 5954 2015
rect 5999 2009 6033 2015
rect 20222 2120 20256 2154
rect 5287 1981 5321 2009
rect 5367 1981 5390 2009
rect 5390 1981 5401 2009
rect 5446 1981 5459 2009
rect 5459 1981 5480 2009
rect 5525 1981 5528 2009
rect 5528 1981 5559 2009
rect 5604 1981 5632 2009
rect 5632 1981 5638 2009
rect 5683 1981 5701 2009
rect 5701 1981 5717 2009
rect 5762 1981 5770 2009
rect 5770 1981 5796 2009
rect 5841 1981 5873 2009
rect 5873 1981 5875 2009
rect 5920 1981 5942 2009
rect 5942 1981 5954 2009
rect 5999 1981 6011 2009
rect 6011 1981 6033 2009
rect 22656 2005 22690 2006
rect 22656 1972 22690 2005
rect 3643 1903 3677 1937
rect 22832 2141 22866 2170
rect 22909 2161 22943 2195
rect 23093 2221 23127 2233
rect 22832 2136 22866 2141
rect 22832 2073 22866 2098
rect 22832 2064 22866 2073
rect 23093 2149 23127 2183
rect 23008 2005 23042 2006
rect 23008 1972 23042 2005
rect 22656 1900 22690 1934
rect 23184 2141 23218 2169
rect 23184 2135 23218 2141
rect 23184 2073 23218 2097
rect 23184 2063 23218 2073
rect 23360 2005 23394 2006
rect 23360 1972 23394 2005
rect 23008 1900 23042 1934
rect 23360 1892 23394 1926
rect 3643 1831 3677 1865
rect 3801 1827 3810 1857
rect 3810 1827 3835 1857
rect 22780 1852 22814 1886
rect 3801 1823 3835 1827
rect 3801 1751 3835 1785
rect 4046 1671 4080 1700
rect 4046 1666 4080 1671
rect 22780 1795 22814 1814
rect 22780 1780 22814 1795
rect 22956 1727 22968 1750
rect 22968 1727 22990 1750
rect 22956 1716 22990 1727
rect 4046 1576 4080 1606
rect 22163 1614 22197 1648
rect 22865 1638 22899 1672
rect 22956 1659 22968 1678
rect 22968 1659 22990 1678
rect 22956 1644 22990 1659
rect 23156 1829 23190 1846
rect 23156 1812 23190 1829
rect 23258 1829 23292 1846
rect 23258 1812 23292 1829
rect 23360 1829 23394 1846
rect 23712 1972 23746 2006
rect 23712 1899 23746 1933
rect 23360 1812 23394 1829
rect 23156 1761 23190 1774
rect 23156 1740 23190 1761
rect 23258 1761 23292 1774
rect 23258 1740 23292 1761
rect 23360 1761 23394 1774
rect 23360 1740 23394 1761
rect 23156 1693 23190 1702
rect 23156 1668 23190 1693
rect 23258 1693 23292 1702
rect 23258 1668 23292 1693
rect 23360 1693 23394 1702
rect 23360 1668 23394 1693
rect 23536 1727 23570 1750
rect 23536 1716 23570 1727
rect 23536 1659 23570 1678
rect 23536 1644 23570 1659
rect 23712 1829 23746 1860
rect 23712 1826 23746 1829
rect 22865 1576 22899 1600
rect 4046 1572 4080 1576
rect 21708 1542 21742 1576
rect 21780 1542 21814 1576
rect 22163 1542 22197 1576
rect 22865 1566 22879 1576
rect 22879 1566 22899 1576
rect 23358 1542 23392 1576
rect 23430 1542 23459 1576
rect 23459 1542 23464 1576
rect 3890 1515 3912 1526
rect 3912 1515 3924 1526
rect 3962 1515 3980 1526
rect 3980 1515 3996 1526
rect 3890 1492 3924 1515
rect 3962 1492 3996 1515
rect 3515 1439 3519 1473
rect 3519 1439 3549 1473
rect 3591 1439 3621 1473
rect 3621 1439 3625 1473
rect 22780 1416 22814 1438
rect 22780 1404 22814 1416
rect 3346 1323 3350 1357
rect 3350 1323 3380 1357
rect 3422 1323 3452 1357
rect 3452 1323 3456 1357
rect 3843 1338 3877 1372
rect 3915 1338 3949 1372
rect 22780 1348 22814 1366
rect 22780 1332 22814 1348
rect 22956 1450 22990 1466
rect 22956 1432 22990 1450
rect 22956 1382 22990 1394
rect 22956 1360 22990 1382
rect 23536 1450 23570 1466
rect 23536 1432 23570 1450
rect 23536 1382 23570 1394
rect 23536 1360 23570 1382
rect 23692 1416 23712 1438
rect 23712 1416 23726 1438
rect 23692 1404 23726 1416
rect 23692 1348 23712 1366
rect 23712 1348 23726 1366
rect 23692 1332 23726 1348
rect 3618 1224 3651 1255
rect 3651 1224 3652 1255
rect 3618 1221 3652 1224
rect 3690 1221 3724 1255
rect 3930 1224 3963 1247
rect 3963 1224 3964 1247
rect 3930 1213 3964 1224
rect 3930 1156 3963 1175
rect 3963 1156 3964 1175
rect 3930 1141 3964 1156
rect 22686 1205 22720 1236
rect 22686 1202 22695 1205
rect 22695 1202 22720 1205
rect 22766 1202 22800 1236
rect 22846 1205 22880 1236
rect 22926 1205 22960 1236
rect 23006 1205 23040 1236
rect 23085 1205 23119 1236
rect 23164 1205 23198 1236
rect 23243 1205 23277 1236
rect 23321 1205 23355 1236
rect 23400 1205 23434 1236
rect 23479 1205 23513 1236
rect 23558 1205 23592 1236
rect 23637 1205 23671 1236
rect 23716 1205 23750 1236
rect 23795 1205 23829 1236
rect 22846 1202 22871 1205
rect 22871 1202 22880 1205
rect 22926 1202 22941 1205
rect 22941 1202 22960 1205
rect 23006 1202 23011 1205
rect 23011 1202 23040 1205
rect 23085 1202 23115 1205
rect 23115 1202 23119 1205
rect 23164 1202 23185 1205
rect 23185 1202 23198 1205
rect 23243 1202 23255 1205
rect 23255 1202 23277 1205
rect 23321 1202 23325 1205
rect 23325 1202 23355 1205
rect 23400 1202 23431 1205
rect 23431 1202 23434 1205
rect 23479 1202 23500 1205
rect 23500 1202 23513 1205
rect 23558 1202 23569 1205
rect 23569 1202 23592 1205
rect 23637 1202 23638 1205
rect 23638 1202 23671 1205
rect 23716 1202 23741 1205
rect 23741 1202 23750 1205
rect 23795 1202 23810 1205
rect 23810 1202 23829 1205
rect 3573 1038 3589 1072
rect 3589 1038 3607 1072
rect 3645 1038 3657 1072
rect 3657 1038 3679 1072
rect 4125 1116 4159 1150
rect 22686 1137 22720 1164
rect 22686 1130 22695 1137
rect 22695 1130 22720 1137
rect 4125 1044 4159 1078
rect 22766 1130 22800 1164
rect 22846 1137 22880 1164
rect 22926 1137 22960 1164
rect 23006 1137 23040 1164
rect 23085 1137 23119 1164
rect 23164 1137 23198 1164
rect 23243 1137 23277 1164
rect 22846 1130 22871 1137
rect 22871 1130 22880 1137
rect 22926 1130 22941 1137
rect 22941 1130 22960 1137
rect 23006 1130 23011 1137
rect 23011 1130 23040 1137
rect 23085 1130 23115 1137
rect 23115 1130 23119 1137
rect 23164 1130 23185 1137
rect 23185 1130 23198 1137
rect 23243 1130 23255 1137
rect 23255 1130 23277 1137
rect 23321 1103 23325 1124
rect 23325 1103 23355 1124
rect 23400 1103 23431 1124
rect 23431 1103 23434 1124
rect 23479 1103 23500 1124
rect 23500 1103 23513 1124
rect 23558 1103 23569 1124
rect 23569 1103 23592 1124
rect 23637 1103 23638 1124
rect 23638 1103 23671 1124
rect 23716 1103 23741 1124
rect 23741 1103 23750 1124
rect 23795 1103 23810 1124
rect 23810 1103 23829 1124
rect 22686 1069 22720 1092
rect 22686 1058 22695 1069
rect 22695 1058 22720 1069
rect 22766 1058 22800 1092
rect 22846 1069 22880 1092
rect 22926 1069 22960 1092
rect 23006 1069 23040 1092
rect 23085 1069 23119 1092
rect 23164 1069 23198 1092
rect 23243 1069 23277 1092
rect 23321 1090 23355 1103
rect 23400 1090 23434 1103
rect 23479 1090 23513 1103
rect 23558 1090 23592 1103
rect 23637 1090 23671 1103
rect 23716 1090 23750 1103
rect 23795 1090 23829 1103
rect 22846 1058 22871 1069
rect 22871 1058 22880 1069
rect 22926 1058 22941 1069
rect 22941 1058 22960 1069
rect 23006 1058 23011 1069
rect 23011 1058 23040 1069
rect 23085 1058 23115 1069
rect 23115 1058 23119 1069
rect 23164 1058 23185 1069
rect 23185 1058 23198 1069
rect 23243 1058 23255 1069
rect 23255 1058 23277 1069
rect 22686 1001 22720 1020
rect 22686 986 22695 1001
rect 22695 986 22720 1001
rect 22766 986 22800 1020
rect 22846 1001 22880 1020
rect 22926 1001 22960 1020
rect 23006 1001 23040 1020
rect 23085 1001 23119 1020
rect 23164 1001 23198 1020
rect 23243 1001 23277 1020
rect 22846 986 22871 1001
rect 22871 986 22880 1001
rect 22926 986 22941 1001
rect 22941 986 22960 1001
rect 23006 986 23011 1001
rect 23011 986 23040 1001
rect 23085 986 23115 1001
rect 23115 986 23119 1001
rect 23164 986 23185 1001
rect 23185 986 23198 1001
rect 23243 986 23255 1001
rect 23255 986 23277 1001
rect 3550 890 3584 894
rect 3550 860 3584 890
rect 3461 793 3495 827
rect 3461 741 3464 755
rect 3464 741 3495 755
rect 3461 721 3495 741
rect 3550 758 3584 792
rect 3640 741 3644 748
rect 3644 741 3674 748
rect 3640 714 3674 741
rect 3712 714 3746 748
rect 3550 660 3584 690
rect 3550 656 3584 660
rect 4011 742 4012 745
rect 4012 742 4045 745
rect 4011 711 4045 742
rect 3858 627 3892 661
rect 3930 627 3964 661
rect 4011 625 4045 659
rect 4011 545 4045 573
rect 4011 539 4012 545
rect 4012 539 4045 545
rect 4011 468 4045 486
rect 4011 452 4012 468
rect 4012 452 4045 468
rect 4011 392 4045 399
rect 4011 365 4012 392
rect 4012 365 4045 392
rect 3858 275 3892 309
rect 3930 275 3964 309
rect 5151 492 5185 526
rect 7547 536 7581 570
rect 6386 509 6420 512
rect 6386 478 6399 509
rect 6399 478 6420 509
rect 6458 478 6492 512
rect 6772 478 6778 512
rect 6778 478 6806 512
rect 6856 478 6887 512
rect 6887 478 6890 512
rect 6939 478 6961 512
rect 6961 478 6973 512
rect 7547 464 7581 498
rect 15914 546 15948 580
rect 16970 546 17004 580
rect 15914 474 15948 508
rect 16001 477 16035 511
rect 5151 420 5185 454
rect 5506 448 5540 452
rect 5506 418 5540 448
rect 6119 448 6153 452
rect 5339 299 5372 309
rect 5372 299 5373 309
rect 5411 299 5440 309
rect 5440 299 5445 309
rect 5339 275 5373 299
rect 5411 275 5445 299
rect 5506 342 5540 375
rect 5506 341 5540 342
rect 5506 270 5540 297
rect 5506 263 5540 270
rect 5506 197 5540 219
rect 5151 163 5185 197
rect 5151 91 5185 125
rect 5506 185 5540 197
rect 6119 418 6129 448
rect 6129 418 6153 448
rect 7294 405 7328 439
rect 16001 405 16035 439
rect 16171 447 16205 481
rect 6119 372 6153 379
rect 6119 345 6129 372
rect 6129 345 6153 372
rect 6119 295 6153 306
rect 5792 249 5826 283
rect 5792 177 5826 211
rect 6119 272 6129 295
rect 6129 272 6153 295
rect 6293 347 6327 381
rect 6293 299 6297 309
rect 6297 299 6327 309
rect 6293 275 6327 299
rect 6544 351 6578 355
rect 6544 321 6578 351
rect 6634 344 6638 378
rect 6638 344 6668 378
rect 6706 344 6740 378
rect 16171 375 16205 409
rect 16266 477 16300 511
rect 16266 405 16300 439
rect 16525 447 16559 481
rect 16525 375 16559 409
rect 16618 447 16652 481
rect 16618 375 16652 409
rect 16883 447 16917 481
rect 16970 474 17004 508
rect 17479 535 17513 569
rect 17479 463 17513 497
rect 16883 375 16917 409
rect 7294 333 7328 367
rect 6544 249 6578 283
rect 6119 218 6153 232
rect 6119 198 6129 218
rect 6129 198 6153 218
rect 6857 188 6876 222
rect 6876 188 6891 222
rect 6929 188 6963 222
rect 5506 124 5540 141
rect 5506 107 5540 124
rect 3773 -1 3807 33
rect 5506 51 5540 63
rect 5506 29 5540 51
rect 6119 124 6153 158
rect 6386 123 6399 157
rect 6399 123 6420 157
rect 6458 123 6492 157
rect 18549 189 18583 223
rect 18628 189 18662 223
rect 18707 189 18741 223
rect 18786 189 18820 223
rect 18865 189 18899 223
rect 18944 189 18978 223
rect 19023 189 19057 223
rect 19101 189 19135 223
rect 7113 101 7147 135
rect 7185 101 7219 135
rect 6119 62 6129 84
rect 6129 62 6153 84
rect 6119 50 6153 62
rect 3773 -73 3807 -39
rect 5265 -53 5270 -19
rect 5270 -53 5299 -19
rect 5337 -53 5338 -19
rect 5338 -53 5371 -19
rect 5506 -22 5540 -15
rect 5506 -49 5540 -22
rect 5506 -95 5540 -93
rect 5506 -127 5540 -95
rect 5266 -229 5270 -195
rect 5270 -229 5300 -195
rect 5338 -229 5372 -195
rect 5410 -229 5440 -195
rect 5440 -229 5444 -195
rect 6299 38 6333 72
rect 6371 38 6405 72
rect 6634 64 6638 98
rect 6638 64 6668 98
rect 6706 64 6740 98
rect 6977 47 7011 81
rect 6119 -14 6129 10
rect 6129 -14 6153 10
rect 6119 -24 6153 -14
rect 6225 -53 6229 -19
rect 6229 -53 6259 -19
rect 6297 -53 6331 -19
rect 6977 -25 7011 9
rect 6119 -91 6129 -64
rect 6129 -91 6153 -64
rect 6119 -98 6153 -91
rect 6119 -168 6129 -138
rect 6129 -168 6153 -138
rect 6119 -172 6153 -168
rect 7303 159 7337 163
rect 7303 129 7337 159
rect 7303 84 7337 86
rect 7303 52 7337 84
rect 18549 81 18583 115
rect 18628 81 18662 115
rect 18707 81 18741 115
rect 18786 81 18820 115
rect 18865 81 18899 115
rect 18944 81 18978 115
rect 19023 81 19057 115
rect 19101 81 19135 115
rect 7303 -26 7337 8
rect 7303 -102 7337 -70
rect 7303 -104 7337 -102
rect 7393 -91 7427 -57
rect 7472 -91 7506 -57
rect 7303 -178 7337 -148
rect 5601 -237 5608 -203
rect 5608 -237 5635 -203
rect 5680 -237 5683 -203
rect 5683 -237 5714 -203
rect 5759 -237 5792 -203
rect 5792 -237 5793 -203
rect 5838 -237 5867 -203
rect 5867 -237 5872 -203
rect 5916 -237 5942 -203
rect 5942 -237 5950 -203
rect 5994 -237 6016 -203
rect 6016 -237 6028 -203
rect 6225 -229 6229 -195
rect 6229 -229 6259 -195
rect 6297 -229 6331 -195
rect 6369 -229 6399 -195
rect 6399 -229 6403 -195
rect 7303 -182 7337 -178
rect 15877 -197 15889 -163
rect 15889 -197 15911 -163
rect 15953 -197 15959 -163
rect 15959 -197 15987 -163
rect 16029 -197 16063 -163
rect 16105 -197 16132 -163
rect 16132 -197 16139 -163
rect 16181 -197 16201 -163
rect 16201 -197 16215 -163
rect 16257 -197 16270 -163
rect 16270 -197 16291 -163
rect 16332 -197 16339 -163
rect 16339 -197 16366 -163
rect 16407 -197 16408 -163
rect 16408 -197 16441 -163
rect 16482 -197 16512 -163
rect 16512 -197 16516 -163
rect 16557 -197 16581 -163
rect 16581 -197 16591 -163
rect 16632 -197 16650 -163
rect 16650 -197 16666 -163
rect 16707 -197 16719 -163
rect 16719 -197 16741 -163
rect 16782 -197 16788 -163
rect 16788 -197 16816 -163
rect 16857 -197 16891 -163
rect 16932 -197 16960 -163
rect 16960 -197 16966 -163
rect 17007 -197 17029 -163
rect 17029 -197 17041 -163
rect 6800 -248 6808 -214
rect 6808 -248 6834 -214
rect 6872 -248 6876 -214
rect 6876 -248 6906 -214
rect 7113 -239 7117 -214
rect 7117 -239 7147 -214
rect 7185 -239 7219 -214
rect 7393 -239 7397 -214
rect 7397 -239 7427 -214
rect 7465 -239 7499 -214
rect 7113 -248 7147 -239
rect 7185 -248 7219 -239
rect 7393 -248 7427 -239
rect 7465 -248 7499 -239
<< metal1 >>
rect 52 3070 58 3122
rect 110 3070 122 3122
rect 174 3070 180 3122
rect 18489 3065 21683 3114
tri 16991 3038 17013 3060 se
rect 17013 3038 18383 3060
tri 18383 3038 18405 3060 sw
rect 108 2986 114 3038
rect 166 2986 178 3038
rect 230 2986 236 3038
tri 16982 3029 16991 3038 se
rect 16991 3029 18405 3038
tri 18405 3029 18414 3038 sw
tri 16969 3016 16982 3029 se
rect 16982 3028 18414 3029
rect 16982 3016 17020 3028
rect 164 2898 170 2950
rect 222 2898 234 2950
rect 286 2898 292 2950
rect 784 2914 3704 3016
tri 16939 2986 16969 3016 se
rect 16969 2989 17020 3016
tri 17020 2989 17059 3028 nw
tri 18369 2998 18399 3028 ne
rect 18399 3013 18414 3028
tri 18414 3013 18430 3029 sw
rect 18489 3013 18495 3065
rect 18547 3013 18567 3065
rect 18619 3062 21683 3065
rect 21735 3062 21755 3114
rect 21807 3062 21813 3114
rect 18619 3013 18625 3062
tri 18685 3013 18701 3029 se
rect 18701 3013 21590 3029
rect 18399 2998 18430 3013
rect 17091 2989 18358 2998
rect 16969 2986 17014 2989
tri 16936 2983 16939 2986 se
rect 16939 2983 17014 2986
tri 17014 2983 17020 2989 nw
tri 17079 2983 17085 2989 se
rect 17085 2983 18358 2989
tri 18358 2983 18373 2998 sw
tri 18399 2983 18414 2998 ne
rect 18414 2986 18430 2998
tri 18430 2986 18457 3013 sw
tri 18658 2986 18685 3013 se
rect 18685 2997 21590 3013
rect 18685 2986 18701 2997
rect 18414 2983 18457 2986
tri 18457 2983 18460 2986 sw
tri 18655 2983 18658 2986 se
rect 18658 2983 18701 2986
tri 18701 2983 18715 2997 nw
tri 21205 2983 21219 2997 ne
rect 21219 2983 21590 2997
tri 16935 2982 16936 2983 se
rect 16936 2982 17013 2983
tri 17013 2982 17014 2983 nw
tri 17078 2982 17079 2983 se
rect 17079 2982 18373 2983
tri 18373 2982 18374 2983 sw
tri 18414 2982 18415 2983 ne
rect 18415 2982 18695 2983
tri 16930 2977 16935 2982 se
rect 16935 2977 17008 2982
tri 17008 2977 17013 2982 nw
tri 17073 2977 17078 2982 se
rect 17078 2977 18374 2982
tri 18374 2977 18379 2982 sw
tri 18415 2977 18420 2982 ne
rect 18420 2977 18695 2982
tri 18695 2977 18701 2983 nw
tri 21219 2977 21225 2983 ne
rect 21225 2977 21590 2983
rect 21642 2977 21662 3029
rect 21714 2977 21720 3029
tri 16920 2967 16930 2977 se
rect 16930 2967 16998 2977
tri 16998 2967 17008 2977 nw
tri 17063 2967 17073 2977 se
rect 17073 2967 18379 2977
tri 18379 2967 18389 2977 sw
tri 18420 2967 18430 2977 ne
rect 18430 2967 18685 2977
tri 18685 2967 18695 2977 nw
tri 16903 2950 16920 2967 se
rect 16920 2950 16974 2967
tri 16899 2946 16903 2950 se
rect 16903 2946 16974 2950
rect 224 2862 276 2868
rect 224 2798 276 2810
rect 224 2740 276 2746
rect 784 2700 839 2914
rect 1226 2806 1442 2914
rect 1226 2754 1232 2806
rect 1284 2754 1308 2806
rect 1360 2754 1383 2806
rect 1435 2754 1442 2806
rect 1226 2714 1442 2754
rect 2110 2736 2116 2788
rect 2168 2736 2180 2788
rect 2232 2736 2238 2788
rect -31 249 2 2654
rect 978 2629 1024 2684
rect 1226 2662 1232 2714
rect 1284 2662 1308 2714
rect 1360 2662 1383 2714
rect 1435 2662 1442 2714
rect 1226 2661 1442 2662
rect 2071 2700 2123 2706
rect 2159 2649 2205 2736
rect 2071 2636 2123 2648
rect 2071 2578 2123 2584
rect 2077 2490 2123 2578
rect 2289 2637 2341 2770
rect 2289 2573 2341 2585
rect 2289 2515 2341 2521
rect 2377 2512 2423 2768
rect 2676 2688 2806 2914
rect 2676 2654 2688 2688
rect 2722 2654 2760 2688
rect 2794 2654 2806 2688
rect 2676 2648 2806 2654
rect 3614 2687 3704 2914
rect 16789 2894 16795 2946
rect 16847 2894 16867 2946
rect 16919 2943 16974 2946
tri 16974 2943 16998 2967 nw
tri 17047 2951 17063 2967 se
rect 17063 2966 18389 2967
tri 18389 2966 18390 2967 sw
tri 18430 2966 18431 2967 ne
rect 18431 2966 18669 2967
rect 17063 2951 17093 2966
tri 17093 2951 17108 2966 nw
tri 18344 2951 18359 2966 ne
rect 18359 2962 18390 2966
tri 18390 2962 18394 2966 sw
tri 18431 2962 18435 2966 ne
rect 18435 2962 18669 2966
rect 18359 2951 18394 2962
tri 18394 2951 18405 2962 sw
tri 18435 2951 18446 2962 ne
rect 18446 2951 18669 2962
tri 18669 2951 18685 2967 nw
tri 18717 2951 18733 2967 se
rect 18733 2951 19548 2967
tri 17039 2943 17047 2951 se
rect 17047 2943 17085 2951
tri 17085 2943 17093 2951 nw
tri 18359 2943 18367 2951 ne
rect 18367 2943 18405 2951
rect 16919 2935 16966 2943
tri 16966 2935 16974 2943 nw
tri 17031 2935 17039 2943 se
rect 17039 2935 17077 2943
tri 17077 2935 17085 2943 nw
tri 18367 2936 18374 2943 ne
rect 18374 2936 18405 2943
tri 17128 2935 17129 2936 se
rect 17129 2935 18332 2936
tri 18332 2935 18333 2936 sw
tri 18374 2935 18375 2936 ne
rect 18375 2935 18405 2936
tri 18405 2935 18421 2951 sw
tri 18701 2935 18717 2951 se
rect 18717 2935 19548 2951
rect 16919 2932 16963 2935
tri 16963 2932 16966 2935 nw
tri 17028 2932 17031 2935 se
rect 17031 2932 17057 2935
rect 16919 2915 16946 2932
tri 16946 2915 16963 2932 nw
tri 17011 2915 17028 2932 se
rect 17028 2915 17057 2932
tri 17057 2915 17077 2935 nw
tri 17108 2915 17128 2935 se
rect 17128 2920 18333 2935
tri 18333 2920 18348 2935 sw
tri 18375 2920 18390 2935 ne
rect 18390 2921 18421 2935
tri 18421 2921 18435 2935 sw
tri 18687 2921 18701 2935 se
rect 18701 2921 18732 2935
rect 18390 2920 18732 2921
tri 18732 2920 18747 2935 nw
tri 19522 2920 19537 2935 ne
rect 19537 2920 19548 2935
rect 17128 2915 18348 2920
tri 18348 2915 18353 2920 sw
tri 18390 2915 18395 2920 ne
rect 18395 2915 18727 2920
tri 18727 2915 18732 2920 nw
tri 19537 2915 19542 2920 ne
rect 19542 2915 19548 2920
rect 19600 2915 19620 2967
rect 19672 2915 19678 2967
tri 19783 2950 19800 2967 se
rect 19800 2950 19874 2967
tri 19768 2935 19783 2950 se
rect 19783 2935 19874 2950
tri 19748 2915 19768 2935 se
rect 19768 2915 19874 2935
rect 19926 2915 19946 2967
rect 19998 2915 20004 2967
tri 20276 2927 20308 2959 se
rect 20308 2927 21171 2959
tri 21171 2927 21203 2959 sw
tri 20264 2915 20276 2927 se
rect 20276 2915 20310 2927
tri 20310 2915 20322 2927 nw
tri 21157 2915 21169 2927 ne
rect 21169 2915 21203 2927
rect 16919 2905 16936 2915
tri 16936 2905 16946 2915 nw
tri 17001 2905 17011 2915 se
rect 17011 2905 17047 2915
tri 17047 2905 17057 2915 nw
rect 17108 2905 18353 2915
tri 18353 2905 18363 2915 sw
tri 18395 2905 18405 2915 ne
rect 18405 2905 18717 2915
tri 18717 2905 18727 2915 nw
tri 19738 2905 19748 2915 se
rect 19748 2905 19766 2915
rect 16919 2894 16925 2905
tri 16925 2894 16936 2905 nw
tri 16993 2897 17001 2905 se
rect 17001 2897 17039 2905
tri 17039 2897 17047 2905 nw
rect 17108 2904 18363 2905
tri 18363 2904 18364 2905 sw
tri 18405 2904 18406 2905 ne
rect 18406 2904 18701 2905
rect 17108 2897 17162 2904
tri 17162 2897 17169 2904 nw
tri 18318 2897 18325 2904 ne
rect 18325 2901 18364 2904
tri 18364 2901 18367 2904 sw
tri 18406 2901 18409 2904 ne
rect 18409 2901 18701 2904
rect 18325 2897 18367 2901
tri 18367 2897 18371 2901 sw
tri 18409 2897 18413 2901 ne
rect 18413 2897 18701 2901
tri 16990 2894 16993 2897 se
rect 16993 2894 17015 2897
tri 16969 2873 16990 2894 se
rect 16990 2873 17015 2894
tri 17015 2873 17039 2897 nw
rect 17108 2889 17154 2897
tri 17154 2889 17162 2897 nw
tri 18325 2889 18333 2897 ne
rect 18333 2889 18371 2897
tri 18371 2889 18379 2897 sw
tri 18413 2889 18421 2897 ne
rect 18421 2889 18701 2897
tri 18701 2889 18717 2905 nw
tri 18743 2889 18759 2905 se
rect 18759 2898 19494 2905
tri 19494 2898 19501 2905 sw
tri 19731 2898 19738 2905 se
rect 19738 2898 19766 2905
rect 18759 2889 19501 2898
tri 16964 2868 16969 2873 se
rect 16969 2868 17010 2873
tri 17010 2868 17015 2873 nw
tri 16960 2864 16964 2868 se
rect 16964 2864 17006 2868
tri 17006 2864 17010 2868 nw
rect 16800 2812 16806 2864
rect 16858 2812 16878 2864
rect 16930 2855 16997 2864
tri 16997 2855 17006 2864 nw
rect 16930 2816 16958 2855
tri 16958 2816 16997 2855 nw
rect 16930 2812 16954 2816
tri 16954 2812 16958 2816 nw
rect 17108 2800 17147 2889
tri 17147 2882 17154 2889 nw
tri 18333 2882 18340 2889 ne
rect 18340 2882 18379 2889
tri 18340 2875 18347 2882 ne
rect 18347 2875 18379 2882
rect 17011 2748 17017 2800
rect 17069 2748 17089 2800
rect 17141 2748 17147 2800
tri 17189 2843 17221 2875 se
rect 17221 2873 18302 2875
tri 18302 2873 18304 2875 sw
tri 18347 2873 18349 2875 ne
rect 18349 2873 18379 2875
tri 18379 2873 18395 2889 sw
tri 18727 2873 18743 2889 se
rect 18743 2887 19501 2889
tri 19501 2887 19512 2898 sw
tri 19720 2887 19731 2898 se
rect 19731 2887 19766 2898
tri 19766 2887 19794 2915 nw
tri 20249 2900 20264 2915 se
rect 20264 2900 20295 2915
tri 20295 2900 20310 2915 nw
tri 21169 2900 21184 2915 ne
rect 21184 2900 21203 2915
tri 20236 2887 20249 2900 se
rect 20249 2887 20282 2900
tri 20282 2887 20295 2900 nw
tri 21184 2887 21197 2900 ne
rect 21197 2887 21203 2900
rect 18743 2873 19752 2887
tri 19752 2873 19766 2887 nw
tri 20235 2886 20236 2887 se
rect 20236 2886 20281 2887
tri 20281 2886 20282 2887 nw
tri 21197 2886 21198 2887 ne
rect 21198 2886 21203 2887
tri 21203 2886 21244 2927 sw
tri 19829 2873 19842 2886 se
rect 19842 2873 20249 2886
rect 17221 2868 18304 2873
tri 18304 2868 18309 2873 sw
tri 18349 2868 18354 2873 ne
rect 18354 2868 18395 2873
rect 17221 2864 18309 2868
tri 18309 2864 18313 2868 sw
tri 18354 2864 18358 2868 ne
rect 18358 2864 18395 2868
rect 17221 2858 18313 2864
tri 18313 2858 18319 2864 sw
tri 18358 2858 18364 2864 ne
rect 18364 2859 18395 2864
tri 18395 2859 18409 2873 sw
tri 18713 2859 18727 2873 se
rect 18727 2868 18768 2873
tri 18768 2868 18773 2873 nw
tri 19480 2868 19485 2873 ne
rect 19485 2868 19734 2873
rect 18727 2859 18758 2868
rect 18364 2858 18758 2859
tri 18758 2858 18768 2868 nw
tri 19485 2858 19495 2868 ne
rect 19495 2858 19734 2868
rect 17221 2855 18319 2858
tri 18319 2855 18322 2858 sw
tri 18364 2855 18367 2858 ne
rect 18367 2855 18755 2858
tri 18755 2855 18758 2858 nw
tri 19495 2855 19498 2858 ne
rect 19498 2855 19734 2858
tri 19734 2855 19752 2873 nw
tri 19811 2855 19829 2873 se
rect 19829 2855 20249 2873
rect 17221 2843 18322 2855
tri 18322 2843 18334 2855 sw
tri 18367 2843 18379 2855 ne
rect 18379 2843 18727 2855
rect 17189 2827 17249 2843
tri 17249 2827 17265 2843 nw
tri 18288 2827 18304 2843 ne
rect 18304 2827 18334 2843
tri 18334 2827 18350 2843 sw
tri 18379 2827 18395 2843 ne
rect 18395 2827 18727 2843
tri 18727 2827 18755 2855 nw
tri 19798 2842 19811 2855 se
rect 19811 2854 20249 2855
tri 20249 2854 20281 2886 nw
tri 21198 2881 21203 2886 ne
rect 21203 2881 21287 2886
tri 21203 2854 21230 2881 ne
rect 21230 2854 21287 2881
rect 19811 2842 19842 2854
tri 18775 2827 18790 2842 se
rect 18790 2840 19455 2842
tri 19455 2840 19457 2842 sw
tri 19796 2840 19798 2842 se
rect 19798 2840 19842 2842
tri 19842 2840 19856 2854 nw
rect 18790 2827 19457 2840
rect 17189 2735 17241 2827
tri 17241 2819 17249 2827 nw
tri 18304 2819 18312 2827 ne
rect 18312 2819 18350 2827
tri 18312 2815 18316 2819 ne
rect 18316 2815 18350 2819
rect 17309 2763 17315 2815
rect 17367 2763 17387 2815
rect 17439 2763 17459 2815
rect 17511 2763 17531 2815
rect 17583 2763 17602 2815
rect 17654 2763 17673 2815
rect 17725 2763 17744 2815
rect 17796 2763 17802 2815
tri 18316 2810 18321 2815 ne
rect 18321 2810 18350 2815
tri 18350 2810 18367 2827 sw
tri 18758 2810 18775 2827 se
rect 18775 2826 19457 2827
tri 19457 2826 19471 2840 sw
tri 19782 2826 19796 2840 se
rect 19796 2826 19828 2840
tri 19828 2826 19842 2840 nw
rect 18775 2816 19818 2826
tri 19818 2816 19828 2826 nw
rect 20845 2821 21159 2827
rect 18775 2810 19812 2816
tri 19812 2810 19818 2816 nw
tri 18321 2808 18323 2810 ne
rect 18323 2808 18367 2810
tri 18323 2797 18334 2808 ne
rect 18334 2797 18367 2808
tri 18367 2797 18380 2810 sw
tri 18745 2797 18758 2810 se
rect 18758 2808 18802 2810
tri 18802 2808 18804 2810 nw
tri 19441 2808 19443 2810 ne
rect 19443 2808 19810 2810
tri 19810 2808 19812 2810 nw
rect 18758 2797 18791 2808
tri 18791 2797 18802 2808 nw
tri 19443 2797 19454 2808 ne
rect 19454 2797 19796 2808
tri 18334 2764 18367 2797 ne
rect 18367 2796 18380 2797
tri 18380 2796 18381 2797 sw
tri 18744 2796 18745 2797 se
rect 18745 2796 18758 2797
rect 18367 2764 18758 2796
tri 18758 2764 18791 2797 nw
tri 19454 2794 19457 2797 ne
rect 19457 2794 19796 2797
tri 19796 2794 19810 2808 nw
rect 17309 2751 17802 2763
rect 17309 2699 17315 2751
rect 17367 2699 17387 2751
rect 17439 2699 17459 2751
rect 17511 2699 17531 2751
rect 17583 2699 17602 2751
rect 17654 2699 17673 2751
rect 17725 2699 17744 2751
rect 17796 2699 17802 2751
rect 20845 2705 20848 2821
rect 21156 2800 21159 2821
tri 21159 2800 21166 2807 sw
rect 21156 2764 21166 2800
tri 21166 2764 21202 2800 sw
rect 21379 2764 21385 2816
rect 21437 2764 21449 2816
rect 21501 2794 21806 2816
tri 21806 2794 21828 2816 sw
rect 21501 2784 22989 2794
rect 21501 2770 21513 2784
tri 21513 2770 21527 2784 nw
tri 21773 2770 21787 2784 ne
rect 21787 2770 22989 2784
rect 21501 2768 21511 2770
tri 21511 2768 21513 2770 nw
tri 21787 2768 21789 2770 ne
rect 21789 2768 22989 2770
rect 21501 2764 21507 2768
tri 21507 2764 21511 2768 nw
tri 21789 2764 21793 2768 ne
rect 21793 2764 22989 2768
rect 21156 2762 21202 2764
tri 21202 2762 21204 2764 sw
tri 21793 2762 21795 2764 ne
rect 21795 2762 22989 2764
rect 21156 2748 21204 2762
tri 21204 2748 21218 2762 sw
tri 22963 2752 22973 2762 ne
rect 22973 2752 22989 2762
rect 21156 2732 21218 2748
tri 21218 2732 21234 2748 sw
rect 21156 2705 21234 2732
rect 20845 2700 21234 2705
tri 21234 2700 21266 2732 sw
rect 21592 2700 21598 2752
rect 21650 2700 21662 2752
rect 21714 2748 21720 2752
tri 21720 2748 21724 2752 sw
tri 22973 2748 22977 2752 ne
rect 22977 2748 22989 2752
rect 21714 2732 21724 2748
tri 21724 2732 21740 2748 sw
tri 22977 2742 22983 2748 ne
rect 22983 2742 22989 2748
rect 23041 2742 23053 2794
rect 23105 2742 23111 2794
rect 21714 2700 22737 2732
rect 20845 2699 21266 2700
rect 21063 2689 21266 2699
rect 3614 2653 3641 2687
rect 3675 2653 3704 2687
tri 21125 2664 21150 2689 ne
rect 21150 2664 21266 2689
tri 21266 2664 21302 2700 sw
tri 22711 2680 22731 2700 ne
rect 22731 2680 22737 2700
rect 22789 2680 22801 2732
rect 22853 2680 22859 2732
tri 21150 2656 21158 2664 ne
rect 21158 2656 21295 2664
rect 3614 2615 3704 2653
rect 3614 2581 3641 2615
rect 3675 2581 3704 2615
tri 21158 2608 21206 2656 ne
rect 21206 2608 21295 2656
rect 3148 2524 3243 2557
tri 3243 2524 3276 2557 sw
rect 3148 2512 3276 2524
tri 3276 2512 3288 2524 sw
tri 2123 2490 2141 2508 sw
tri 2359 2490 2377 2508 se
rect 2377 2490 2383 2512
rect 2077 2486 2141 2490
tri 2141 2486 2145 2490 sw
tri 2355 2486 2359 2490 se
rect 2359 2486 2383 2490
rect 2077 2459 2178 2486
tri 2178 2459 2205 2486 sw
tri 2295 2459 2322 2486 se
rect 2322 2460 2383 2486
rect 2435 2460 2447 2512
rect 2499 2460 2505 2512
rect 3148 2511 3288 2512
tri 3212 2490 3233 2511 ne
rect 3233 2490 3288 2511
tri 3288 2490 3310 2512 sw
tri 3233 2488 3235 2490 ne
rect 3235 2488 3310 2490
tri 3310 2488 3312 2490 sw
tri 3235 2480 3243 2488 ne
rect 3243 2480 3312 2488
tri 3243 2477 3246 2480 ne
rect 3246 2477 3312 2480
rect 3154 2471 3206 2477
tri 3246 2474 3249 2477 ne
rect 2322 2459 2423 2460
rect 2077 2457 2160 2459
tri 2143 2447 2153 2457 ne
rect 2153 2447 2160 2457
tri 2153 2440 2160 2447 ne
rect 2340 2457 2423 2459
rect 2340 2447 2347 2457
tri 2347 2447 2357 2457 nw
tri 2340 2440 2347 2447 nw
rect 1143 2427 1189 2433
tri 1189 2427 1195 2433 sw
rect 1143 2421 1195 2427
rect 1143 2357 1195 2369
rect 1340 2421 1392 2427
rect 1143 2297 1195 2305
rect 1143 2240 1189 2297
tri 1189 2291 1195 2297 nw
rect 890 1978 942 2040
tri 1260 1775 1262 1777 se
rect 1262 1775 1308 2368
tri 1226 1741 1260 1775 se
rect 1260 1741 1308 1775
tri 1201 1716 1226 1741 se
rect 1226 1716 1308 1741
tri 1192 1707 1201 1716 se
rect 1201 1707 1299 1716
tri 1299 1707 1308 1716 nw
rect 1340 2357 1392 2369
rect 3154 2407 3206 2419
rect 3249 2467 3312 2477
rect 3249 2415 3255 2467
rect 3307 2415 3319 2467
rect 3371 2415 3377 2467
rect 3154 2349 3206 2355
rect 3614 2356 3704 2581
rect 1340 1724 1392 2305
rect 3614 2322 3643 2356
rect 3677 2322 3704 2356
rect 3614 2284 3704 2322
rect 3614 2250 3643 2284
rect 3677 2250 3704 2284
rect 793 1546 845 1552
rect 793 1482 845 1494
rect 793 1424 845 1430
rect 1192 1505 1299 1707
rect 1340 1660 1392 1672
rect 1340 1602 1392 1608
rect 2159 1752 2341 2092
rect 3614 1949 3704 2250
rect 4040 2596 4086 2608
rect 4040 2562 4046 2596
rect 4080 2562 4086 2596
tri 21206 2572 21242 2608 ne
rect 21242 2572 21295 2608
rect 4040 2524 4086 2562
rect 4040 2490 4046 2524
rect 4080 2490 4086 2524
rect 4040 2281 4086 2490
rect 17627 2453 17633 2505
rect 17685 2453 17699 2505
rect 17751 2453 17757 2505
rect 17808 2430 17814 2482
rect 17866 2430 17880 2482
rect 17932 2430 17938 2482
rect 18798 2470 18804 2522
rect 18856 2470 18868 2522
rect 18920 2470 18926 2522
rect 19159 2476 19484 2522
rect 20710 2459 20716 2511
rect 20768 2459 20780 2511
rect 20832 2459 20838 2511
rect 20891 2459 20897 2511
rect 20949 2459 20961 2511
rect 21013 2459 21019 2511
rect 22820 2453 22872 2459
rect 22407 2367 22413 2419
rect 22465 2367 22477 2419
rect 22529 2367 22535 2419
rect 22820 2389 22872 2401
rect 4040 2247 4046 2281
rect 4080 2247 4086 2281
rect 4040 2184 4086 2247
rect 4040 2150 4046 2184
rect 4080 2150 4086 2184
rect 4040 2086 4086 2150
rect 4040 2052 4046 2086
rect 4080 2052 4086 2086
rect 3848 2029 3978 2035
rect 3848 1995 3860 2029
rect 3894 1995 3932 2029
rect 3966 1995 3978 2029
rect 3848 1989 3978 1995
tri 3848 1981 3856 1989 ne
rect 3856 1981 3950 1989
tri 3950 1981 3958 1989 nw
tri 3856 1972 3865 1981 ne
rect 3865 1972 3941 1981
tri 3941 1972 3950 1981 nw
tri 3865 1957 3880 1972 ne
rect 3363 1937 3704 1949
rect 3363 1903 3369 1937
rect 3403 1903 3643 1937
rect 3677 1903 3704 1937
rect 3363 1865 3704 1903
rect 3363 1831 3369 1865
rect 3403 1831 3643 1865
rect 3677 1831 3704 1865
rect 3363 1819 3704 1831
rect 3789 1863 3841 1869
rect 3880 1825 3926 1972
tri 3926 1957 3941 1972 nw
rect 4040 1924 4086 2052
rect 3958 1872 3964 1924
rect 4016 1872 4028 1924
rect 4080 1872 4086 1924
rect 4119 2333 4165 2345
rect 4119 2299 4125 2333
rect 4159 2299 4165 2333
rect 4119 2261 4165 2299
rect 18575 2290 18581 2342
rect 18633 2290 18645 2342
rect 18697 2290 18703 2342
rect 19964 2290 19970 2342
rect 20022 2290 20034 2342
rect 20086 2290 20092 2342
rect 22820 2331 22872 2337
rect 23072 2407 23078 2459
rect 23130 2407 23142 2459
rect 23194 2447 23224 2459
rect 23218 2413 23224 2447
rect 23194 2407 23224 2413
rect 23072 2375 23224 2407
rect 23072 2341 23184 2375
rect 23218 2341 23224 2375
rect 23072 2334 23224 2341
tri 22820 2325 22826 2331 ne
rect 4119 2227 4125 2261
rect 4159 2227 4165 2261
rect 21359 2245 21365 2297
rect 21417 2245 21429 2297
rect 21481 2245 21487 2297
rect 3789 1799 3841 1811
rect 3452 1775 3498 1787
rect 2159 1700 2197 1752
rect 2249 1700 2261 1752
rect 2313 1700 2341 1752
rect 3091 1700 3097 1752
rect 3149 1700 3161 1752
rect 3213 1700 3219 1752
rect 3452 1741 3458 1775
rect 3492 1741 3498 1775
rect 3872 1773 3878 1825
rect 3930 1773 3942 1825
rect 3994 1773 4000 1825
rect 3789 1741 3841 1747
rect 1735 1546 1787 1552
rect 1192 1492 1253 1505
tri 1253 1492 1266 1505 nw
rect 793 1291 839 1424
rect 1192 1323 1240 1492
tri 1240 1479 1253 1492 nw
rect 1735 1482 1787 1494
rect 1735 1424 1787 1430
tri 1240 1323 1253 1336 sw
rect 1192 1314 1253 1323
tri 1253 1314 1262 1323 sw
rect 1192 1303 1262 1314
tri 1192 1291 1204 1303 ne
rect 1204 1291 1262 1303
tri 1204 1282 1213 1291 ne
rect 1213 1282 1262 1291
rect 793 1276 845 1282
tri 1213 1255 1240 1282 ne
rect 1240 1255 1262 1282
tri 1262 1255 1321 1314 sw
rect 1735 1276 1787 1282
tri 1240 1233 1262 1255 ne
rect 1262 1233 1321 1255
tri 1321 1233 1343 1255 sw
rect 793 1212 845 1224
tri 1262 1221 1274 1233 ne
rect 1274 1221 1343 1233
tri 1274 1213 1282 1221 ne
rect 1282 1213 1343 1221
tri 1282 1202 1293 1213 ne
rect 1293 1202 1343 1213
tri 1293 1200 1295 1202 ne
rect 793 1154 845 1160
rect 1295 352 1343 1202
rect 1735 1212 1787 1224
rect 1735 1154 1787 1160
rect 2159 1083 2341 1700
rect 3452 1671 3498 1741
rect 3795 1739 3841 1741
rect 3452 1637 3458 1671
rect 3492 1637 3498 1671
rect 3452 1572 3498 1637
rect 4040 1700 4086 1712
rect 4040 1666 4046 1700
rect 4080 1666 4086 1700
rect 4040 1619 4086 1666
tri 3498 1572 3512 1586 sw
rect 3452 1567 3512 1572
tri 3512 1567 3517 1572 sw
rect 3958 1567 3964 1619
rect 4016 1567 4028 1619
rect 4080 1567 4086 1619
rect 2770 1546 2822 1552
rect 3452 1533 3458 1567
rect 3492 1553 3706 1567
tri 3706 1553 3720 1567 sw
rect 4040 1560 4086 1567
rect 3492 1533 3720 1553
rect 3452 1521 3720 1533
rect 3880 1532 3886 1538
tri 3666 1507 3680 1521 ne
rect 2770 1482 2822 1494
tri 3272 1473 3278 1479 se
rect 3278 1473 3637 1479
rect 2770 1424 2822 1430
tri 3264 1465 3272 1473 se
rect 3272 1465 3515 1473
rect 3264 1439 3515 1465
rect 3549 1439 3591 1473
rect 3625 1439 3637 1473
rect 3264 1433 3637 1439
rect 2770 1276 2822 1282
rect 2770 1212 2822 1224
rect 2770 1154 2822 1160
rect 3264 1078 3304 1433
tri 3304 1419 3318 1433 nw
tri 3675 1372 3680 1377 se
rect 3680 1372 3720 1521
rect 3878 1486 3886 1532
rect 3938 1486 3950 1538
rect 4002 1486 4008 1538
rect 3831 1398 3838 1450
rect 3890 1398 3902 1450
rect 3954 1398 3961 1450
tri 3720 1372 3729 1381 sw
rect 3831 1372 3961 1398
tri 3669 1366 3675 1372 se
rect 3675 1366 3729 1372
tri 3729 1366 3735 1372 sw
rect 3334 1314 3340 1366
rect 3392 1314 3406 1366
rect 3458 1363 3464 1366
rect 3458 1317 3468 1363
rect 3458 1314 3464 1317
rect 3669 1314 3675 1366
rect 3727 1314 3739 1366
rect 3791 1314 3797 1366
rect 3831 1338 3843 1372
rect 3877 1338 3915 1372
rect 3949 1338 3961 1372
rect 3831 1332 3961 1338
rect 3606 1212 3612 1264
rect 3664 1212 3678 1264
rect 3730 1212 3736 1264
rect 3924 1247 3970 1259
rect 3924 1213 3930 1247
rect 3964 1213 3970 1247
rect 3924 1175 3970 1213
rect 3924 1141 3930 1175
rect 3964 1141 3970 1175
tri 3304 1078 3308 1082 sw
rect 3264 1072 3308 1078
tri 3308 1072 3314 1078 sw
rect 3455 1072 3691 1078
rect 3264 1063 3314 1072
tri 3314 1063 3323 1072 sw
rect 3264 1011 3304 1063
rect 3356 1011 3368 1063
rect 3420 1011 3426 1063
rect 3455 1038 3573 1072
rect 3607 1038 3645 1072
rect 3679 1038 3691 1072
rect 3455 1032 3691 1038
rect 3455 1020 3522 1032
tri 3522 1020 3534 1032 nw
rect 3455 839 3506 1020
tri 3506 1004 3522 1020 nw
tri 3909 1004 3924 1019 se
rect 3924 1004 3970 1141
rect 4119 1150 4165 2227
rect 20213 2232 20265 2238
tri 18282 2192 18283 2193 sw
rect 18282 2170 18283 2192
tri 18283 2170 18305 2192 sw
rect 18282 2154 18305 2170
tri 18305 2154 18321 2170 sw
rect 20213 2168 20265 2180
rect 18282 2153 18321 2154
tri 18321 2153 18322 2154 sw
rect 17662 2061 17668 2113
rect 17720 2061 17738 2113
rect 17790 2061 17796 2113
rect 18019 2061 18025 2113
rect 18077 2061 18095 2113
rect 18147 2061 18153 2113
rect 18282 2101 18424 2153
rect 18476 2101 18488 2153
rect 18540 2101 18546 2153
rect 18282 2100 18311 2101
tri 18311 2100 18312 2101 nw
rect 18878 2100 18884 2152
rect 18936 2100 18948 2152
rect 19000 2100 19006 2152
rect 19634 2100 19640 2152
rect 19692 2100 19704 2152
rect 19756 2100 19762 2152
rect 22360 2135 22413 2196
rect 22826 2170 22872 2331
tri 23144 2300 23178 2334 ne
rect 22826 2136 22832 2170
rect 22866 2136 22872 2170
rect 22903 2273 22955 2279
rect 22903 2207 22955 2221
rect 22903 2149 22955 2155
rect 23084 2261 23136 2267
rect 23084 2195 23136 2209
rect 23084 2137 23136 2143
rect 23178 2169 23224 2334
rect 20213 2110 20265 2116
rect 20216 2108 20262 2110
rect 18282 2098 18309 2100
tri 18309 2098 18311 2100 nw
tri 18282 2071 18309 2098 nw
rect 18715 2053 18767 2059
rect 20501 2058 20507 2110
rect 20559 2058 20571 2110
rect 20623 2058 20629 2110
rect 20969 2058 20975 2110
rect 21027 2058 21039 2110
rect 21091 2058 21097 2110
rect 22826 2098 22872 2136
rect 22826 2064 22832 2098
rect 22866 2064 22872 2098
rect 5275 2015 6045 2021
rect 5275 1981 5287 2015
rect 5321 1981 5367 2015
rect 5401 1981 5446 2015
rect 5480 1981 5525 2015
rect 5559 1981 5604 2015
rect 5638 1981 5683 2015
rect 5717 1981 5762 2015
rect 5796 1981 5841 2015
rect 5875 1981 5920 2015
rect 5954 1981 5999 2015
rect 6033 1981 6045 2015
rect 5275 1975 6045 1981
rect 22826 2052 22872 2064
rect 23178 2135 23184 2169
rect 23218 2135 23224 2169
tri 23576 2166 23610 2200 sw
rect 23178 2097 23224 2135
rect 23178 2063 23184 2097
rect 23218 2063 23224 2097
rect 23178 2051 23224 2063
tri 21341 2006 21362 2027 se
rect 21362 2018 22612 2027
tri 22612 2018 22621 2027 sw
rect 21362 2008 23461 2018
tri 23461 2008 23471 2018 sw
tri 23696 2008 23706 2018 se
rect 23706 2008 23849 2018
rect 21362 2006 23849 2008
rect 18715 1989 18767 2001
rect 5278 1973 5313 1975
tri 21307 1972 21341 2006 se
rect 21341 1972 22656 2006
rect 22690 1972 23008 2006
rect 23042 1972 23360 2006
rect 23394 1972 23712 2006
rect 23746 1972 23849 2006
rect 8202 1928 8254 1934
rect 18715 1931 18767 1937
tri 21292 1957 21307 1972 se
rect 21307 1957 23849 1972
rect 21292 1934 23849 1957
rect 4522 1872 4528 1924
rect 4580 1872 4592 1924
rect 4644 1904 4650 1924
rect 4644 1872 4853 1904
rect 4727 1832 4779 1838
rect 4727 1768 4779 1780
rect 4554 1700 4560 1752
rect 4612 1700 4624 1752
rect 4676 1700 4694 1752
rect 4488 1490 4494 1542
rect 4546 1490 4558 1542
rect 4610 1490 4616 1542
rect 4485 1444 4537 1450
rect 4485 1380 4537 1392
rect 4321 1314 4327 1366
rect 4379 1314 4391 1366
rect 4443 1314 4449 1366
tri 4367 1286 4395 1314 ne
rect 4119 1116 4125 1150
rect 4159 1116 4165 1150
rect 4119 1078 4165 1116
rect 4119 1044 4125 1078
rect 4159 1044 4165 1078
tri 3970 1004 3985 1019 sw
tri 3908 1003 3909 1004 se
rect 3909 1003 3985 1004
tri 3985 1003 3986 1004 sw
rect 3866 951 3872 1003
rect 3924 951 3938 1003
rect 3990 951 3996 1003
rect 3454 833 3506 839
tri 1343 352 1347 356 sw
rect 1295 345 1347 352
rect 1295 281 1347 293
tri 2 249 11 258 sw
rect -31 240 11 249
tri 11 240 20 249 sw
rect -31 106 20 240
rect 1295 223 1347 229
rect 1295 219 1343 223
tri 1343 219 1347 223 nw
rect 1295 218 1342 219
tri 1342 218 1343 219 nw
tri 1781 125 1785 129 sw
rect 1781 121 1785 125
tri 1785 121 1789 125 sw
rect 1781 106 1789 121
tri 1789 106 1804 121 sw
rect 1781 99 1804 106
tri 1804 99 1811 106 sw
rect 2206 99 2335 831
rect 3454 767 3506 781
rect 3454 709 3506 715
rect 3455 703 3506 709
rect 3544 894 3590 906
rect 3544 860 3550 894
rect 3584 860 3590 894
rect 3864 871 3870 923
rect 3922 871 3934 923
rect 3986 871 3992 923
rect 3544 792 3590 860
tri 3880 845 3906 871 ne
rect 3544 758 3550 792
rect 3584 758 3590 792
rect 3544 690 3590 758
rect 3906 757 3952 871
tri 3952 845 3978 871 nw
rect 4119 839 4165 1044
rect 4304 1278 4357 1284
rect 4304 1226 4305 1278
rect 4304 1214 4357 1226
rect 4304 1162 4305 1214
tri 3952 757 3987 792 sw
rect 4035 787 4041 839
rect 4093 787 4107 839
rect 4159 787 4166 839
tri 4098 769 4116 787 ne
rect 4116 769 4166 787
tri 4116 759 4126 769 ne
rect 3754 754 3802 755
rect 3628 748 3802 754
rect 3628 714 3640 748
rect 3674 714 3712 748
rect 3746 714 3802 748
rect 3906 745 4051 757
rect 3906 741 4011 745
tri 3906 718 3929 741 ne
rect 3929 718 4011 741
rect 3628 708 3802 714
tri 3981 711 3988 718 ne
rect 3988 711 4011 718
rect 4045 711 4051 745
rect 3544 656 3550 690
rect 3584 656 3590 690
tri 3513 495 3544 526 se
rect 3544 495 3590 656
tri 3590 495 3621 526 sw
rect 3506 443 3512 495
rect 3564 443 3576 495
rect 3628 443 3634 495
rect 3370 313 3422 319
rect 3754 316 3802 708
tri 3988 694 4005 711 ne
rect 3846 616 3852 668
rect 3904 616 3918 668
rect 3970 616 3976 668
rect 4005 659 4051 711
rect 4005 625 4011 659
rect 4045 625 4051 659
rect 4005 573 4051 625
rect 4005 539 4011 573
rect 4045 539 4051 573
rect 4005 486 4051 539
rect 4005 452 4011 486
rect 4045 452 4051 486
rect 4005 399 4051 452
rect 4005 365 4011 399
rect 4045 365 4051 399
rect 4005 353 4051 365
tri 4125 353 4126 354 se
rect 4126 353 4166 769
tri 4113 341 4125 353 se
rect 4125 341 4166 353
tri 4093 321 4113 341 se
rect 4113 321 4166 341
tri 4088 316 4093 321 se
rect 4093 316 4166 321
rect 3686 264 3692 316
rect 3744 264 3756 316
rect 3808 264 3814 316
tri 4087 315 4088 316 se
rect 4088 315 4166 316
rect 3846 309 4166 315
rect 3846 275 3858 309
rect 3892 275 3930 309
rect 3964 275 4166 309
rect 3846 269 4166 275
rect 3370 249 3422 261
rect 3370 191 3422 197
rect 4304 226 4357 1162
rect 4304 174 4305 226
rect 4304 162 4357 174
rect 3265 138 3312 150
rect 3259 132 3312 138
rect 1781 94 1811 99
rect 1735 93 1811 94
tri 1735 91 1737 93 ne
rect 1737 91 1811 93
tri 1811 91 1819 99 sw
tri 2197 91 2205 99 se
rect 2205 91 2335 99
tri 2335 91 2343 99 sw
tri 1737 84 1744 91 ne
rect 1744 84 1819 91
tri 1819 84 1826 91 sw
tri 2191 85 2197 91 se
rect 2197 85 2343 91
tri 2343 85 2349 91 sw
tri 1744 63 1765 84 ne
rect 1765 63 1826 84
tri 1826 63 1847 84 sw
tri 1765 39 1789 63 ne
rect 1789 33 1847 63
tri 1847 33 1877 63 sw
rect 2191 33 2197 85
rect 2249 33 2299 85
rect 2351 33 2357 85
rect 3311 80 3312 132
rect 4304 110 4305 162
rect 4304 104 4357 110
rect 4395 145 4449 1314
rect 1789 23 1877 33
tri 1877 23 1887 33 sw
rect 1789 21 1887 23
tri 1887 21 1889 23 sw
tri 2774 21 2776 23 se
rect 2776 21 2822 77
rect 3259 68 3312 80
rect 1789 5 1889 21
tri 1889 5 1905 21 sw
tri 2758 5 2774 21 se
rect 2774 10 2822 21
tri 2822 10 2833 21 sw
rect 3311 16 3312 68
rect 4395 93 4396 145
rect 4448 93 4449 145
rect 4395 81 4449 93
rect 3259 12 3312 16
rect 3767 33 3813 45
rect 3259 10 3311 12
rect 2774 5 2833 10
rect 1789 -1 2833 5
tri 2833 -1 2844 10 sw
rect 3767 -1 3773 33
rect 3807 -1 3813 33
rect 4395 29 4396 81
rect 4448 29 4449 81
rect 4395 23 4449 29
rect 4485 62 4537 1328
rect 4569 316 4616 1490
rect 4652 668 4694 1700
rect 4727 1710 4779 1716
rect 4727 755 4769 1710
rect 4821 824 4853 1872
rect 8202 1864 8254 1876
rect 21292 1900 22656 1934
rect 22690 1900 23008 1934
rect 23042 1933 23849 1934
rect 23042 1926 23712 1933
rect 23042 1900 23360 1926
rect 21292 1892 23360 1900
rect 23394 1899 23712 1926
rect 23746 1899 23849 1933
rect 23394 1892 23849 1899
rect 21292 1886 23849 1892
tri 14219 1852 14226 1859 se
rect 14226 1852 14581 1859
tri 14581 1852 14588 1859 sw
tri 14213 1846 14219 1852 se
rect 14219 1846 14588 1852
tri 14588 1846 14594 1852 sw
tri 14206 1839 14213 1846 se
rect 14213 1839 14594 1846
tri 14594 1839 14601 1846 sw
rect 8202 1799 8254 1812
rect 14200 1820 14761 1839
rect 14200 1814 14242 1820
tri 14242 1814 14248 1820 nw
tri 14531 1814 14537 1820 ne
rect 14537 1814 14761 1820
rect 14200 1793 14221 1814
tri 14221 1793 14242 1814 nw
tri 14537 1801 14550 1814 ne
rect 14550 1792 14761 1814
rect 8202 1734 8254 1747
rect 8202 1676 8254 1682
rect 14441 1785 14493 1791
rect 14441 1721 14493 1733
rect 14441 1663 14493 1669
rect 14441 1583 14447 1635
rect 14499 1583 14511 1635
rect 14563 1583 14569 1635
rect 17500 1502 18137 1838
rect 18562 1649 19386 1860
rect 21292 1852 22780 1886
rect 22814 1860 23849 1886
rect 22814 1852 23712 1860
rect 21292 1846 23712 1852
rect 21292 1830 23156 1846
rect 20740 1791 20868 1818
rect 20740 1739 20746 1791
rect 20798 1739 20810 1791
rect 20862 1739 20868 1791
rect 20740 1712 20868 1739
rect 21292 1715 21721 1830
tri 22559 1814 22575 1830 ne
rect 22575 1814 23156 1830
tri 22728 1800 22742 1814 ne
rect 22742 1800 22780 1814
tri 22742 1780 22762 1800 ne
rect 22762 1780 22780 1800
rect 22814 1812 22864 1814
tri 22864 1812 22866 1814 nw
tri 23080 1812 23082 1814 ne
rect 23082 1812 23156 1814
rect 23190 1812 23258 1846
rect 23292 1812 23360 1846
rect 23394 1826 23712 1846
rect 23746 1826 23849 1860
rect 23394 1814 23849 1826
rect 23394 1812 23456 1814
rect 22814 1800 22852 1812
tri 22852 1800 22864 1812 nw
tri 23082 1800 23094 1812 ne
rect 23094 1800 23456 1812
tri 23456 1800 23470 1814 nw
rect 22814 1780 22826 1800
tri 22762 1774 22768 1780 ne
rect 22768 1774 22826 1780
tri 22826 1774 22852 1800 nw
tri 23094 1774 23120 1800 ne
rect 23120 1774 23418 1800
tri 22768 1768 22774 1774 ne
rect 22774 1768 22820 1774
tri 22820 1768 22826 1774 nw
tri 23120 1768 23126 1774 ne
rect 23126 1768 23156 1774
tri 23126 1762 23132 1768 ne
rect 23132 1762 23156 1768
rect 22950 1750 22996 1762
rect 22950 1716 22956 1750
rect 22990 1716 22996 1750
tri 23132 1744 23150 1762 ne
rect 22853 1678 22905 1684
rect 21771 1666 21823 1672
rect 18562 1648 19298 1649
tri 19298 1648 19299 1649 nw
rect 18562 1550 19264 1648
tri 19264 1614 19298 1648 nw
tri 21769 1614 21771 1616 se
tri 21755 1600 21769 1614 se
rect 21769 1600 21823 1614
tri 21737 1582 21755 1600 se
rect 21755 1594 21823 1600
rect 21755 1582 21771 1594
rect 21696 1576 21771 1582
rect 22154 1655 22206 1661
rect 22154 1583 22206 1603
rect 21696 1542 21708 1576
rect 21742 1542 21771 1576
rect 21823 1542 21826 1582
rect 21696 1536 21826 1542
rect 22853 1612 22905 1626
rect 22853 1554 22905 1560
rect 22950 1678 22996 1716
rect 22950 1644 22956 1678
rect 22990 1644 22996 1678
rect 23150 1740 23156 1762
rect 23190 1740 23258 1774
rect 23292 1740 23360 1774
rect 23394 1762 23418 1774
tri 23418 1762 23456 1800 nw
rect 23394 1750 23406 1762
tri 23406 1750 23418 1762 nw
rect 23530 1750 23576 1762
rect 23394 1740 23400 1750
tri 23400 1744 23406 1750 nw
rect 23150 1702 23400 1740
rect 23150 1668 23156 1702
rect 23190 1668 23258 1702
rect 23292 1668 23360 1702
rect 23394 1668 23400 1702
rect 23150 1656 23400 1668
rect 23530 1716 23536 1750
rect 23570 1716 23576 1750
rect 23530 1678 23576 1716
rect 22154 1525 22206 1531
rect 21890 1452 21944 1515
rect 22246 1435 22290 1496
rect 22950 1479 22996 1644
rect 23530 1644 23536 1678
rect 23570 1644 23576 1678
rect 23224 1533 23230 1585
rect 23282 1533 23294 1585
rect 23346 1576 23476 1585
rect 23346 1542 23358 1576
rect 23392 1542 23430 1576
rect 23464 1542 23476 1576
rect 23346 1533 23476 1542
tri 23499 1482 23530 1513 se
rect 23530 1482 23576 1644
tri 22996 1479 22999 1482 sw
tri 23496 1479 23499 1482 se
rect 23499 1479 23576 1482
rect 22950 1476 22999 1479
tri 22999 1476 23002 1479 sw
rect 22950 1470 23002 1476
rect 22774 1438 22820 1450
rect 22774 1404 22780 1438
rect 22814 1404 22820 1438
rect 18230 1369 18282 1375
rect 22774 1366 22820 1404
rect 22774 1332 22780 1366
rect 22814 1332 22820 1366
rect 22950 1406 23002 1418
rect 22950 1348 23002 1354
rect 23327 1473 23576 1479
rect 23379 1466 23576 1473
rect 23379 1433 23536 1466
rect 23379 1432 23412 1433
tri 23412 1432 23413 1433 nw
tri 23496 1432 23497 1433 ne
rect 23497 1432 23536 1433
rect 23570 1432 23576 1466
rect 23379 1421 23384 1432
rect 23327 1409 23384 1421
rect 23379 1404 23384 1409
tri 23384 1404 23412 1432 nw
tri 23497 1404 23525 1432 ne
rect 23525 1404 23576 1432
tri 23379 1399 23384 1404 nw
tri 23525 1399 23530 1404 ne
rect 23327 1351 23379 1357
rect 23530 1394 23576 1404
rect 23530 1360 23536 1394
rect 23570 1360 23576 1394
rect 23530 1348 23576 1360
rect 23686 1438 23732 1450
rect 23686 1404 23692 1438
rect 23726 1404 23732 1438
rect 23686 1366 23732 1404
rect 18230 1305 18282 1317
rect 18230 1247 18282 1253
rect 18326 1322 18378 1328
rect 18326 1258 18378 1270
tri 22740 1242 22774 1276 se
rect 22774 1242 22820 1332
rect 23686 1332 23692 1366
rect 23726 1332 23732 1366
tri 22820 1242 22854 1276 sw
tri 23652 1242 23686 1276 se
rect 23686 1242 23732 1332
tri 23732 1242 23766 1276 sw
rect 18326 1200 18378 1206
rect 22654 1236 23841 1242
rect 22654 1202 22686 1236
rect 22720 1202 22766 1236
rect 22800 1202 22846 1236
rect 22880 1202 22926 1236
rect 22960 1202 23006 1236
rect 23040 1202 23085 1236
rect 23119 1202 23164 1236
rect 23198 1202 23243 1236
rect 23277 1202 23321 1236
rect 23355 1202 23400 1236
rect 23434 1202 23479 1236
rect 23513 1202 23558 1236
rect 23592 1202 23637 1236
rect 23671 1202 23716 1236
rect 23750 1202 23795 1236
rect 23829 1202 23841 1236
rect 17662 1146 17668 1198
rect 17720 1146 17738 1198
rect 17790 1146 17796 1198
rect 18019 1145 18025 1197
rect 18077 1145 18095 1197
rect 18147 1145 18153 1197
tri 21764 1164 21791 1191 sw
tri 22043 1164 22070 1191 se
rect 21764 1157 21791 1164
tri 21791 1157 21798 1164 sw
tri 22036 1157 22043 1164 se
rect 22043 1157 22070 1164
tri 22116 1164 22143 1191 sw
tri 22395 1164 22422 1191 se
rect 22116 1157 22143 1164
tri 22143 1157 22150 1164 sw
tri 22388 1157 22395 1164 se
rect 22395 1157 22422 1164
rect 22654 1164 23841 1202
rect 18846 1105 18852 1157
rect 18904 1105 18916 1157
rect 18968 1105 18974 1157
rect 21718 1094 22468 1157
rect 22654 1130 22686 1164
rect 22720 1130 22766 1164
rect 22800 1130 22846 1164
rect 22880 1130 22926 1164
rect 22960 1130 23006 1164
rect 23040 1130 23085 1164
rect 23119 1130 23164 1164
rect 23198 1130 23243 1164
rect 23277 1130 23841 1164
rect 22654 1124 23841 1130
rect 21718 1092 22042 1094
tri 22042 1092 22044 1094 nw
rect 22654 1092 23321 1124
rect 21718 1077 22008 1092
rect 21718 1025 21726 1077
rect 21778 1025 21804 1077
rect 21856 1058 22008 1077
tri 22008 1058 22042 1092 nw
rect 22654 1058 22686 1092
rect 22720 1058 22766 1092
rect 22800 1058 22846 1092
rect 22880 1058 22926 1092
rect 22960 1058 23006 1092
rect 23040 1058 23085 1092
rect 23119 1058 23164 1092
rect 23198 1058 23243 1092
rect 23277 1090 23321 1092
rect 23355 1090 23400 1124
rect 23434 1090 23479 1124
rect 23513 1090 23558 1124
rect 23592 1090 23637 1124
rect 23671 1090 23716 1124
rect 23750 1090 23795 1124
rect 23829 1090 23841 1124
rect 23277 1084 23841 1090
rect 23277 1058 23309 1084
rect 21856 1025 21970 1058
rect 21718 1020 21970 1025
tri 21970 1020 22008 1058 nw
rect 22654 1020 23309 1058
rect 21718 1007 21957 1020
tri 21957 1007 21970 1020 nw
rect 22543 1006 22595 1012
tri 14068 986 14088 1006 se
rect 14088 986 15777 1006
tri 15777 986 15797 1006 sw
tri 14048 966 14068 986 se
rect 14068 968 15797 986
tri 15797 968 15815 986 sw
rect 14068 966 15815 968
tri 15815 966 15817 968 sw
tri 14005 923 14048 966 se
rect 14048 923 15817 966
rect 5460 871 5466 923
rect 5518 871 5530 923
rect 5582 871 5588 923
rect 6631 871 6637 923
rect 6689 871 6703 923
rect 6755 871 6761 923
tri 13998 916 14005 923 se
rect 14005 916 15817 923
rect 18547 916 18553 968
rect 18605 916 18617 968
rect 18669 916 18675 968
rect 22654 986 22686 1020
rect 22720 986 22766 1020
rect 22800 986 22846 1020
rect 22880 986 22926 1020
rect 22960 986 23006 1020
rect 23040 986 23085 1020
rect 23119 986 23164 1020
rect 23198 986 23243 1020
rect 23277 986 23309 1020
rect 22654 980 23309 986
rect 22543 942 22595 954
tri 22519 916 22543 940 se
tri 13953 871 13998 916 se
rect 13998 871 14094 916
tri 5474 845 5500 871 ne
rect 4821 792 4932 824
rect 4727 703 4733 755
rect 4785 703 4797 755
rect 4849 703 4855 755
rect 4652 616 4658 668
rect 4710 616 4722 668
rect 4774 616 4780 668
rect 4569 264 4575 316
rect 4627 264 4639 316
rect 4691 264 4697 316
rect 4485 10 4491 62
rect 4543 10 4555 62
rect 4607 10 4613 62
rect 1789 -15 2844 -1
tri 2844 -15 2858 -1 sw
rect 1789 -19 2858 -15
tri 2858 -19 2862 -15 sw
rect 1789 -20 2862 -19
tri 2862 -20 2863 -19 sw
rect 3767 -20 3813 -1
rect 1789 -39 3813 -20
rect 1789 -73 3773 -39
rect 3807 -73 3813 -39
rect 1789 -87 3813 -73
rect 4900 -362 4932 792
rect 5327 787 5333 839
rect 5385 787 5399 839
rect 5451 787 5457 839
tri 5375 769 5393 787 ne
rect 5210 616 5216 668
rect 5268 616 5282 668
rect 5334 616 5340 668
tri 5223 590 5249 616 ne
rect 5145 526 5213 539
rect 5145 492 5151 526
rect 5185 492 5213 526
rect 5145 454 5213 492
rect 5145 420 5151 454
rect 5185 420 5213 454
rect 5145 197 5213 420
rect 5145 163 5151 197
rect 5185 163 5213 197
rect 5145 125 5213 163
rect 5145 91 5151 125
rect 5185 91 5213 125
rect 5145 -172 5213 91
rect 5249 10 5295 616
tri 5295 590 5321 616 nw
tri 5380 321 5393 334 se
rect 5393 321 5439 787
tri 5439 769 5457 787 nw
rect 5500 536 5546 871
tri 5546 845 5572 871 nw
tri 6643 847 6667 871 ne
rect 6492 787 6498 839
rect 6550 787 6564 839
rect 6616 787 6622 839
tri 6520 769 6538 787 ne
rect 6240 703 6246 755
rect 6298 703 6312 755
rect 6364 703 6370 755
tri 6269 685 6287 703 ne
tri 5546 536 5564 554 sw
rect 5500 535 5564 536
tri 5564 535 5565 536 sw
rect 5500 530 5565 535
tri 5565 530 5570 535 sw
rect 5500 484 5639 530
rect 5500 478 5565 484
tri 5565 478 5571 484 nw
rect 5500 464 5551 478
tri 5551 464 5565 478 nw
rect 5500 452 5546 464
tri 5546 459 5551 464 nw
rect 5500 418 5506 452
rect 5540 418 5546 452
rect 5500 375 5546 418
rect 5500 341 5506 375
rect 5540 341 5546 375
tri 5439 321 5452 334 sw
tri 5374 315 5380 321 se
rect 5380 315 5452 321
tri 5452 315 5458 321 sw
rect 5327 309 5458 315
rect 5327 275 5339 309
rect 5373 275 5411 309
rect 5445 275 5458 309
rect 5327 269 5458 275
rect 5500 297 5546 341
rect 5500 263 5506 297
rect 5540 263 5546 297
rect 6113 452 6159 464
rect 6113 418 6119 452
rect 6153 418 6159 452
rect 6113 379 6159 418
rect 6113 345 6119 379
rect 6153 345 6159 379
rect 6113 306 6159 345
rect 5500 219 5546 263
rect 5786 283 5832 295
rect 5786 249 5792 283
rect 5826 249 5832 283
rect 5786 241 5832 249
rect 5500 185 5506 219
rect 5540 185 5546 219
rect 5500 141 5546 185
rect 5500 107 5506 141
rect 5540 107 5546 141
rect 5500 63 5546 107
rect 5500 29 5506 63
rect 5540 29 5546 63
tri 5295 10 5309 24 sw
rect 5249 -13 5309 10
tri 5309 -13 5332 10 sw
rect 5249 -19 5383 -13
rect 5249 -53 5265 -19
rect 5299 -53 5337 -19
rect 5371 -53 5383 -19
rect 5249 -59 5383 -53
rect 5500 -15 5546 29
rect 5500 -49 5506 -15
rect 5540 -49 5546 -15
rect 5500 -93 5546 -49
rect 5500 -127 5506 -93
rect 5540 -127 5546 -93
rect 5500 -139 5546 -127
rect 5574 211 5832 241
rect 5574 187 5792 211
tri 5213 -172 5219 -166 sw
rect 5574 -170 5609 187
rect 5786 177 5792 187
rect 5826 177 5832 211
rect 5786 165 5832 177
rect 6113 272 6119 306
rect 6153 272 6159 306
rect 6113 232 6159 272
rect 6113 198 6119 232
rect 6153 198 6159 232
rect 6113 158 6159 198
rect 6113 124 6119 158
rect 6153 124 6159 158
rect 6113 84 6159 124
rect 6113 50 6119 84
rect 6153 50 6159 84
rect 6113 10 6159 50
rect 6113 -24 6119 10
rect 6153 -24 6159 10
rect 6113 -64 6159 -24
rect 6199 395 6251 401
rect 6199 322 6251 343
rect 6199 9 6251 270
rect 6287 381 6333 703
tri 6333 685 6351 703 nw
rect 6287 347 6293 381
rect 6327 347 6333 381
rect 6287 309 6333 347
rect 6287 275 6293 309
rect 6327 275 6333 309
rect 6287 78 6333 275
rect 6374 469 6380 521
rect 6432 469 6446 521
rect 6498 469 6504 521
rect 6374 188 6504 469
rect 6538 355 6584 787
tri 6584 769 6602 787 nw
tri 6661 405 6667 411 se
rect 6667 405 6725 871
tri 6725 847 6749 871 nw
tri 13945 863 13953 871 se
rect 13953 863 14094 871
tri 11396 859 11400 863 se
rect 11400 859 11829 863
tri 11829 859 11833 863 sw
tri 13941 859 13945 863 se
rect 13945 859 14094 863
tri 14094 859 14151 916 nw
tri 15636 859 15693 916 ne
rect 15693 859 15817 916
tri 22509 906 22519 916 se
rect 22519 906 22543 916
tri 22062 883 22085 906 se
rect 22085 890 22543 906
tri 23468 941 23502 975 sw
rect 22085 883 22595 890
tri 11384 847 11396 859 se
rect 11396 847 14045 859
tri 11347 810 11384 847 se
rect 11384 810 14045 847
tri 14045 810 14094 859 nw
tri 15693 858 15694 859 ne
rect 15694 828 15817 859
rect 21570 877 21622 883
tri 11345 808 11347 810 se
rect 11347 808 14043 810
tri 14043 808 14045 810 nw
rect 11276 807 14007 808
rect 8502 772 14007 807
tri 14007 772 14043 808 nw
rect 8502 765 13947 772
tri 13947 765 13954 772 nw
rect 8502 758 11463 765
tri 11463 758 11470 765 nw
tri 13671 758 13678 765 ne
rect 13678 758 13940 765
tri 13940 758 13947 765 nw
rect 8502 750 11455 758
tri 11455 750 11463 758 nw
tri 13678 750 13686 758 ne
rect 13686 750 13932 758
tri 13932 750 13940 758 nw
rect 8502 738 11443 750
tri 11443 738 11455 750 nw
tri 13686 738 13698 750 ne
rect 13698 739 13921 750
tri 13921 739 13932 750 nw
rect 13698 738 13714 739
rect 8502 606 11419 738
tri 11419 714 11443 738 nw
tri 13698 722 13714 738 ne
rect 11276 605 11419 606
rect 7541 570 7587 582
rect 7541 536 7547 570
rect 7581 536 7587 570
rect 6760 469 6766 521
rect 6818 469 6832 521
rect 6884 512 7017 521
rect 6890 478 6939 512
rect 6973 478 7017 512
rect 6884 469 7017 478
tri 6922 464 6927 469 ne
rect 6927 464 7017 469
tri 6927 447 6944 464 ne
rect 6944 447 7017 464
rect 7541 498 7587 536
rect 7541 464 7547 498
rect 7581 464 7587 498
tri 6944 441 6950 447 ne
tri 6725 405 6731 411 sw
tri 6640 384 6661 405 se
rect 6661 384 6731 405
tri 6731 384 6752 405 sw
rect 6538 321 6544 355
rect 6578 321 6584 355
rect 6622 378 6752 384
rect 6622 344 6634 378
rect 6668 344 6706 378
rect 6740 344 6752 378
rect 6622 338 6752 344
rect 6538 283 6584 321
rect 6538 249 6544 283
rect 6578 249 6584 283
rect 6538 237 6584 249
tri 6923 237 6950 264 se
rect 6950 237 7017 447
rect 7288 439 7334 451
rect 7288 405 7294 439
rect 7328 405 7334 439
rect 7288 388 7334 405
tri 7334 388 7346 400 sw
tri 6918 232 6923 237 se
rect 6923 232 7017 237
tri 6504 188 6520 204 sw
rect 6374 163 6520 188
tri 6520 163 6545 188 sw
rect 6624 180 6630 232
rect 6682 180 6694 232
rect 6746 180 6752 232
tri 6914 228 6918 232 se
rect 6918 228 7017 232
rect 6845 222 7017 228
rect 6845 188 6857 222
rect 6891 188 6929 222
rect 6963 188 7017 222
rect 6845 182 7017 188
rect 7053 271 7158 388
rect 7288 377 7346 388
tri 7346 377 7357 388 sw
rect 7288 375 7357 377
tri 7357 375 7359 377 sw
tri 7539 375 7541 377 se
rect 7541 375 7587 464
rect 7288 367 7359 375
rect 7288 333 7294 367
rect 7328 353 7359 367
tri 7359 353 7381 375 sw
tri 7517 353 7539 375 se
rect 7539 353 7587 375
rect 7328 333 7587 353
rect 7288 330 7587 333
rect 7288 321 7578 330
tri 7578 321 7587 330 nw
tri 7288 308 7301 321 ne
rect 7301 308 7556 321
tri 7158 271 7195 308 sw
tri 7301 299 7310 308 ne
rect 7310 299 7556 308
tri 7556 299 7578 321 nw
tri 7353 271 7381 299 ne
rect 7381 271 7528 299
tri 7528 271 7556 299 nw
rect 7053 251 7323 271
tri 7323 251 7343 271 sw
rect 7053 183 7343 251
rect 6374 157 6545 163
rect 6374 123 6386 157
rect 6420 123 6458 157
rect 6492 135 6545 157
tri 6545 135 6573 163 sw
rect 6492 123 6573 135
tri 6573 123 6585 135 sw
rect 6374 117 6585 123
tri 6419 104 6432 117 ne
rect 6432 104 6585 117
rect 6624 104 6752 180
tri 6904 175 6911 182 ne
rect 6911 175 7017 182
tri 7267 175 7275 183 ne
rect 7275 175 7343 183
tri 6911 163 6923 175 ne
rect 6923 163 7017 175
tri 7275 163 7287 175 ne
rect 7287 163 7343 175
tri 6923 153 6933 163 ne
rect 6933 153 7017 163
tri 7287 153 7297 163 ne
tri 6933 144 6942 153 ne
rect 6942 144 7017 153
tri 6942 136 6950 144 ne
tri 6432 101 6435 104 ne
rect 6435 101 6585 104
tri 6435 98 6438 101 ne
rect 6438 98 6585 101
tri 6438 82 6454 98 ne
rect 6287 72 6417 78
rect 6287 38 6299 72
rect 6333 38 6371 72
rect 6405 38 6417 72
rect 6287 32 6417 38
tri 6251 9 6270 28 sw
rect 6199 -13 6270 9
tri 6270 -13 6292 9 sw
rect 6199 -19 6343 -13
rect 6199 -53 6225 -19
rect 6259 -53 6297 -19
rect 6331 -53 6343 -19
rect 6199 -59 6343 -53
rect 6113 -98 6119 -64
rect 6153 -98 6159 -64
rect 6113 -138 6159 -98
rect 5145 -182 5219 -172
tri 5219 -182 5229 -172 sw
rect 5145 -184 5229 -182
tri 5229 -184 5231 -182 sw
rect 5145 -189 5231 -184
tri 5231 -189 5236 -184 sw
rect 5574 -189 6079 -170
rect 6113 -172 6119 -138
rect 6153 -172 6159 -138
rect 6113 -184 6159 -172
rect 5145 -195 6079 -189
rect 5145 -229 5266 -195
rect 5300 -229 5338 -195
rect 5372 -229 5410 -195
rect 5444 -203 6079 -195
rect 5444 -229 5601 -203
rect 5145 -237 5601 -229
rect 5635 -237 5680 -203
rect 5714 -237 5759 -203
rect 5793 -237 5838 -203
rect 5872 -237 5916 -203
rect 5950 -237 5994 -203
rect 6028 -214 6079 -203
rect 6213 -195 6415 -189
rect 6213 -214 6225 -195
rect 6028 -229 6225 -214
rect 6259 -229 6297 -195
rect 6331 -229 6369 -195
rect 6403 -214 6415 -195
rect 6454 -214 6585 98
rect 6622 98 6752 104
rect 6622 64 6634 98
rect 6668 64 6706 98
rect 6740 64 6752 98
rect 6622 58 6752 64
rect 6950 81 7017 144
rect 7101 92 7107 144
rect 7159 92 7171 144
rect 7223 141 7229 144
rect 7223 95 7231 141
rect 7297 129 7303 163
rect 7337 129 7343 163
rect 7223 92 7229 95
rect 6403 -229 6585 -214
rect 6028 -237 6585 -229
rect 5145 -257 6585 -237
rect 6788 10 6794 62
rect 6846 10 6860 62
rect 6912 10 6918 62
rect 6788 -214 6918 10
rect 6788 -248 6800 -214
rect 6834 -248 6872 -214
rect 6906 -248 6918 -214
rect 6788 -254 6918 -248
rect 6950 47 6977 81
rect 7011 47 7017 81
rect 6950 9 7017 47
rect 6950 -25 6977 9
rect 7011 -25 7017 9
rect 6950 -182 7017 -25
rect 7297 86 7343 129
rect 7297 52 7303 86
rect 7337 52 7343 86
rect 7297 8 7343 52
rect 7297 -26 7303 8
rect 7337 -26 7343 8
rect 7297 -70 7343 -26
rect 7297 -104 7303 -70
rect 7337 -104 7343 -70
rect 7297 -148 7343 -104
tri 7017 -182 7034 -165 sw
rect 7297 -182 7303 -148
rect 7337 -182 7343 -148
rect 6950 -194 7034 -182
tri 7034 -194 7046 -182 sw
rect 7297 -194 7343 -182
rect 7381 -57 7518 271
tri 7518 261 7528 271 nw
rect 7381 -91 7393 -57
rect 7427 -91 7472 -57
rect 7506 -91 7518 -57
rect 6950 -197 7046 -194
tri 7046 -197 7049 -194 sw
rect 6950 -203 7049 -197
tri 7049 -203 7055 -197 sw
rect 6950 -208 7055 -203
tri 7055 -208 7060 -203 sw
rect 6950 -214 7231 -208
tri 7231 -214 7237 -208 sw
tri 7375 -214 7381 -208 se
rect 7381 -214 7518 -91
rect 15694 24 15818 828
rect 21570 813 21622 825
rect 17629 758 17635 810
rect 17687 758 17699 810
rect 17751 758 17757 810
rect 17950 750 17956 802
rect 18008 750 18020 802
rect 18072 750 18078 802
rect 18735 738 18741 790
rect 18793 738 18805 790
rect 18857 738 18863 790
rect 21570 738 21622 761
rect 21652 877 22595 883
rect 21704 867 22595 877
rect 22693 921 22745 927
tri 22689 867 22693 871 se
rect 22693 867 22745 869
rect 21704 844 22077 867
tri 22077 844 22100 867 nw
tri 22666 844 22689 867 se
rect 22689 857 22745 867
rect 22689 844 22693 857
rect 21704 837 21731 844
tri 21731 837 21738 844 nw
tri 22659 837 22666 844 se
rect 22666 837 22693 844
rect 21652 813 21704 825
tri 21704 810 21731 837 nw
tri 22084 810 22111 837 se
rect 22111 810 22693 837
tri 22073 799 22084 810 se
rect 22084 805 22693 810
rect 22084 799 22745 805
tri 22057 783 22073 799 se
rect 22073 783 22111 799
tri 22111 783 22127 799 nw
tri 22039 765 22057 783 se
rect 22057 765 22093 783
tri 22093 765 22111 783 nw
rect 21652 755 21704 761
tri 21815 755 21825 765 se
rect 21825 755 22055 765
tri 21802 742 21815 755 se
rect 21815 742 22055 755
tri 21622 738 21626 742 sw
tri 21798 738 21802 742 se
rect 21802 738 22055 742
rect 21570 711 21626 738
tri 21626 711 21653 738 sw
tri 21771 711 21798 738 se
rect 21798 727 22055 738
tri 22055 727 22093 765 nw
rect 21798 711 21825 727
tri 21825 711 21841 727 nw
rect 21570 708 21653 711
tri 21653 708 21656 711 sw
tri 21768 708 21771 711 se
rect 21771 708 21822 711
tri 21822 708 21825 711 nw
rect 21570 673 21787 708
tri 21787 673 21822 708 nw
tri 19067 597 19099 629 se
rect 19099 597 19254 629
tri 19063 593 19067 597 se
rect 19067 593 19109 597
tri 19109 593 19113 597 nw
tri 19228 593 19232 597 ne
rect 19232 593 19254 597
rect 15905 587 15957 593
rect 15905 520 15957 535
rect 16961 587 17013 593
tri 19060 590 19063 593 se
rect 19063 590 19098 593
tri 17577 582 17585 590 se
tri 19052 582 19060 590 se
rect 19060 582 19098 590
tri 19098 582 19109 593 nw
tri 19232 582 19243 593 ne
rect 19243 582 19254 593
tri 17576 581 17577 582 se
rect 17577 581 17585 582
tri 17461 569 17473 581 se
rect 17473 569 17519 581
tri 17519 569 17531 581 sw
tri 17564 569 17576 581 se
rect 17576 569 17585 581
tri 19039 569 19052 582 se
rect 15905 462 15957 468
rect 15992 517 16044 523
rect 16257 517 16309 523
rect 15992 451 16044 465
rect 15992 393 16044 399
rect 16162 481 16214 493
rect 16162 447 16171 481
rect 16205 447 16214 481
rect 16162 431 16214 447
rect 16961 520 17013 535
rect 16257 451 16309 465
rect 16257 393 16309 399
rect 16516 481 16568 493
rect 16516 447 16525 481
rect 16559 447 16568 481
rect 16516 409 16568 447
rect 16162 375 16171 379
rect 16205 375 16214 379
rect 16162 367 16214 375
rect 16162 309 16214 315
rect 16516 375 16525 409
rect 16559 375 16568 409
rect 16516 280 16568 375
rect 16609 487 16661 493
rect 16609 421 16661 435
rect 16609 363 16661 369
rect 16874 487 16926 493
rect 16961 462 17013 468
rect 17473 535 17479 569
rect 17513 535 17519 569
tri 19038 568 19039 569 se
rect 19039 568 19052 569
rect 17473 497 17519 535
rect 18126 516 18132 568
rect 18184 516 18196 568
rect 18248 536 19052 568
tri 19052 536 19098 582 nw
tri 19243 577 19248 582 ne
rect 19248 577 19254 582
rect 19306 577 19318 629
rect 19370 577 19376 629
tri 21702 601 21718 617 se
rect 21718 612 21862 618
tri 21461 577 21485 601 se
tri 21451 567 21461 577 se
rect 21461 567 21485 577
tri 21537 577 21561 601 sw
tri 21678 577 21702 601 se
rect 21702 577 21718 601
rect 21537 567 21561 577
tri 21561 567 21571 577 sw
tri 21668 567 21678 577 se
rect 21678 567 21718 577
tri 21637 536 21668 567 se
rect 21668 560 21718 567
rect 21770 560 21810 612
rect 21668 536 21862 560
rect 18248 526 18264 536
tri 18264 526 18274 536 nw
tri 21627 526 21637 536 se
rect 21637 526 21862 536
rect 18248 516 18254 526
tri 18254 516 18264 526 nw
tri 19097 516 19107 526 se
rect 19107 516 19254 526
tri 19087 506 19097 516 se
rect 19097 506 19254 516
rect 17473 463 17479 497
rect 17513 463 17519 497
rect 17473 451 17519 463
tri 18287 462 18290 465 se
rect 18290 462 18296 506
tri 18279 454 18287 462 se
rect 18287 454 18296 462
rect 18348 454 18360 506
rect 18412 474 19254 506
rect 19306 474 19318 526
rect 19370 474 19376 526
tri 21594 493 21627 526 se
rect 21627 523 21862 526
rect 21627 493 21718 523
rect 19561 488 21718 493
rect 18412 454 18418 474
tri 18276 451 18279 454 se
rect 18279 451 18322 454
rect 16874 421 16926 435
tri 18236 411 18276 451 se
rect 18276 411 18282 451
tri 18282 411 18322 451 nw
rect 16874 363 16926 369
tri 18190 365 18236 411 se
tri 18236 365 18282 411 nw
tri 18188 363 18190 365 se
rect 18190 363 18234 365
tri 18234 363 18236 365 nw
tri 18175 350 18188 363 se
rect 18188 350 18201 363
tri 17998 330 18018 350 se
rect 18018 330 18201 350
tri 18201 330 18234 363 nw
rect 17386 278 17392 330
rect 17444 278 17456 330
rect 17508 319 18190 330
tri 18190 319 18201 330 nw
rect 17508 298 18012 319
tri 18012 298 18033 319 nw
rect 19561 308 20746 488
rect 20862 471 21718 488
rect 21770 471 21810 523
rect 20862 465 21862 471
rect 22087 479 22139 485
rect 20862 462 21858 465
tri 21858 462 21861 465 nw
rect 20862 363 21759 462
tri 21759 363 21858 462 nw
rect 22087 415 22139 427
tri 21932 363 21958 389 se
rect 21958 363 22087 389
rect 20862 308 21693 363
rect 17508 297 17647 298
rect 19561 297 21693 308
tri 21693 297 21759 363 nw
tri 21926 357 21932 363 se
rect 21932 357 22139 363
tri 21912 343 21926 357 se
rect 21926 343 21968 357
tri 21968 343 21982 357 nw
tri 21866 297 21912 343 se
rect 21912 333 21958 343
tri 21958 333 21968 343 nw
rect 17508 278 17514 297
tri 21856 287 21866 297 se
rect 21866 287 21912 297
tri 21912 287 21958 333 nw
tri 21847 278 21856 287 se
tri 21828 259 21847 278 se
rect 21847 259 21856 278
tri 19356 229 19386 259 se
rect 19386 229 20135 259
rect 16516 216 16568 228
rect 18537 223 19147 229
rect 18537 189 18549 223
rect 18583 189 18628 223
rect 18662 189 18707 223
rect 18741 189 18786 223
rect 18820 189 18865 223
rect 18899 189 18944 223
rect 18978 189 19023 223
rect 19057 189 19101 223
rect 19135 189 19147 223
tri 19334 207 19356 229 se
rect 19356 207 20135 229
rect 20187 207 20199 259
rect 20251 207 20257 259
tri 21800 231 21828 259 se
rect 21828 231 21856 259
tri 21856 231 21912 287 nw
tri 21776 207 21800 231 se
rect 16516 158 16568 164
rect 17477 173 17529 179
rect 17477 109 17529 121
rect 18537 115 19147 189
tri 19312 185 19334 207 se
rect 19334 185 19386 207
tri 19386 185 19408 207 nw
tri 21754 185 21776 207 se
rect 21776 185 21800 207
tri 19306 179 19312 185 se
rect 19312 179 19380 185
tri 19380 179 19386 185 nw
tri 21748 179 21754 185 se
rect 21754 179 21800 185
tri 19302 175 19306 179 se
rect 19306 175 19376 179
tri 19376 175 19380 179 nw
tri 21744 175 21748 179 se
rect 21748 175 21800 179
tri 21800 175 21856 231 nw
tri 19250 123 19302 175 se
rect 19302 123 19324 175
tri 19324 123 19376 175 nw
rect 19481 123 19973 175
rect 20025 123 20037 175
rect 20089 141 21766 175
tri 21766 141 21800 175 nw
rect 20089 123 21418 141
rect 17529 98 17725 103
tri 17725 98 17730 103 sw
rect 17529 81 17730 98
tri 17730 81 17747 98 sw
rect 18537 81 18549 115
rect 18583 81 18628 115
rect 18662 81 18707 115
rect 18741 81 18786 115
rect 18820 81 18865 115
rect 18899 81 18944 115
rect 18978 81 19023 115
rect 19057 81 19101 115
rect 19135 81 19147 115
tri 19238 111 19250 123 se
rect 19250 111 19312 123
tri 19312 111 19324 123 nw
tri 19230 103 19238 111 se
tri 19225 98 19230 103 se
rect 19230 98 19238 103
rect 17529 57 17747 81
rect 17477 51 17747 57
tri 17703 47 17707 51 ne
rect 17707 47 17747 51
tri 15818 24 15841 47 sw
tri 17707 24 17730 47 ne
rect 17730 24 17747 47
tri 17747 24 17804 81 sw
rect 18537 75 19147 81
tri 19202 75 19225 98 se
rect 19225 75 19238 98
tri 19164 37 19202 75 se
rect 19202 37 19238 75
tri 19238 37 19312 111 nw
tri 19156 29 19164 37 se
rect 19164 29 19230 37
tri 19230 29 19238 37 nw
rect 15694 6 15841 24
tri 15841 6 15859 24 sw
tri 17730 6 17748 24 ne
rect 17748 6 17804 24
tri 17804 6 17822 24 sw
rect 15694 -50 17692 6
tri 17692 -50 17748 6 sw
tri 17748 -50 17804 6 ne
rect 17804 -18 17822 6
tri 17822 -18 17846 6 sw
rect 17804 -50 17846 -18
tri 17846 -50 17878 -18 sw
rect 18699 -23 19178 29
tri 19178 -23 19230 29 nw
rect 15694 -62 17748 -50
tri 17748 -62 17760 -50 sw
tri 17804 -62 17816 -50 ne
rect 17816 -62 18461 -50
rect 15694 -92 17760 -62
tri 17760 -92 17790 -62 sw
tri 17816 -92 17846 -62 ne
rect 17846 -92 18461 -62
rect 15694 -102 17790 -92
tri 17790 -102 17800 -92 sw
tri 17846 -102 17856 -92 ne
rect 17856 -102 18461 -92
rect 18513 -102 18525 -50
rect 18577 -102 18583 -50
rect 15694 -114 17800 -102
tri 17800 -114 17812 -102 sw
rect 18751 -114 18757 -62
rect 18809 -114 18821 -62
rect 18873 -114 18879 -62
rect 15694 -148 17812 -114
tri 17812 -148 17846 -114 sw
rect 15694 -149 18873 -148
rect 15694 -163 18586 -149
rect 15694 -197 15877 -163
rect 15911 -197 15953 -163
rect 15987 -197 16029 -163
rect 16063 -197 16105 -163
rect 16139 -197 16181 -163
rect 16215 -197 16257 -163
rect 16291 -197 16332 -163
rect 16366 -197 16407 -163
rect 16441 -197 16482 -163
rect 16516 -197 16557 -163
rect 16591 -197 16632 -163
rect 16666 -197 16707 -163
rect 16741 -197 16782 -163
rect 16816 -197 16857 -163
rect 16891 -197 16932 -163
rect 16966 -197 17007 -163
rect 17041 -197 18586 -163
rect 15694 -201 18586 -197
rect 18638 -201 18650 -149
rect 18702 -201 18987 -149
rect 15694 -203 18987 -201
rect 6950 -248 7113 -214
rect 7147 -248 7185 -214
rect 7219 -224 7237 -214
tri 7237 -224 7247 -214 sw
tri 7365 -224 7375 -214 se
rect 7375 -224 7393 -214
rect 7219 -248 7393 -224
rect 7427 -248 7465 -214
rect 7499 -224 7518 -214
tri 7518 -224 7534 -208 sw
rect 7499 -248 7534 -224
rect 5145 -263 6670 -257
tri 6670 -263 6676 -257 sw
rect 5145 -284 6676 -263
tri 6676 -284 6697 -263 sw
tri 6929 -284 6950 -263 se
rect 6950 -284 7534 -248
rect 5145 -322 7534 -284
tri 6618 -346 6642 -322 ne
rect 6642 -346 7534 -322
rect 4816 -414 4822 -362
rect 4874 -414 4886 -362
rect 4938 -414 4944 -362
<< via1 >>
rect 58 3070 110 3122
rect 122 3070 174 3122
rect 114 2986 166 3038
rect 178 2986 230 3038
rect 170 2898 222 2950
rect 234 2898 286 2950
rect 18495 3013 18547 3065
rect 18567 3013 18619 3065
rect 21683 3062 21735 3114
rect 21755 3062 21807 3114
rect 21590 2977 21642 3029
rect 21662 2977 21714 3029
rect 224 2810 276 2862
rect 224 2746 276 2798
rect 1232 2754 1284 2806
rect 1308 2754 1360 2806
rect 1383 2754 1435 2806
rect 2116 2736 2168 2788
rect 2180 2736 2232 2788
rect 1232 2662 1284 2714
rect 1308 2662 1360 2714
rect 1383 2662 1435 2714
rect 2071 2648 2123 2700
rect 2071 2584 2123 2636
rect 2289 2585 2341 2637
rect 2289 2521 2341 2573
rect 16795 2894 16847 2946
rect 16867 2894 16919 2946
rect 19548 2915 19600 2967
rect 19620 2915 19672 2967
rect 19874 2915 19926 2967
rect 19946 2915 19998 2967
rect 16806 2812 16858 2864
rect 16878 2812 16930 2864
rect 17017 2748 17069 2800
rect 17089 2748 17141 2800
rect 17315 2763 17367 2815
rect 17387 2763 17439 2815
rect 17459 2763 17511 2815
rect 17531 2763 17583 2815
rect 17602 2763 17654 2815
rect 17673 2763 17725 2815
rect 17744 2763 17796 2815
rect 17315 2699 17367 2751
rect 17387 2699 17439 2751
rect 17459 2699 17511 2751
rect 17531 2699 17583 2751
rect 17602 2699 17654 2751
rect 17673 2699 17725 2751
rect 17744 2699 17796 2751
rect 20848 2705 21156 2821
rect 21385 2764 21437 2816
rect 21449 2764 21501 2816
rect 21598 2700 21650 2752
rect 21662 2700 21714 2752
rect 22989 2742 23041 2794
rect 23053 2742 23105 2794
rect 22737 2680 22789 2732
rect 22801 2680 22853 2732
rect 2383 2460 2435 2512
rect 2447 2460 2499 2512
rect 1143 2369 1195 2421
rect 1340 2369 1392 2421
rect 1143 2305 1195 2357
rect 1340 2305 1392 2357
rect 3154 2419 3206 2471
rect 3255 2415 3307 2467
rect 3319 2415 3371 2467
rect 3154 2355 3206 2407
rect 793 1494 845 1546
rect 793 1430 845 1482
rect 1340 1672 1392 1724
rect 1340 1608 1392 1660
rect 17633 2453 17685 2505
rect 17699 2453 17751 2505
rect 17814 2430 17866 2482
rect 17880 2430 17932 2482
rect 18804 2470 18856 2522
rect 18868 2470 18920 2522
rect 20716 2459 20768 2511
rect 20780 2459 20832 2511
rect 20897 2459 20949 2511
rect 20961 2459 21013 2511
rect 22820 2447 22872 2453
rect 22413 2367 22465 2419
rect 22477 2367 22529 2419
rect 22820 2413 22832 2447
rect 22832 2413 22866 2447
rect 22866 2413 22872 2447
rect 22820 2401 22872 2413
rect 22820 2375 22872 2389
rect 3789 1857 3841 1863
rect 3789 1823 3801 1857
rect 3801 1823 3835 1857
rect 3835 1823 3841 1857
rect 3964 1872 4016 1924
rect 4028 1872 4080 1924
rect 18581 2290 18633 2342
rect 18645 2290 18697 2342
rect 19970 2290 20022 2342
rect 20034 2290 20086 2342
rect 22820 2341 22832 2375
rect 22832 2341 22866 2375
rect 22866 2341 22872 2375
rect 22820 2337 22872 2341
rect 23078 2407 23130 2459
rect 23142 2447 23194 2459
rect 23142 2413 23184 2447
rect 23184 2413 23194 2447
rect 23142 2407 23194 2413
rect 21365 2245 21417 2297
rect 21429 2245 21481 2297
rect 3789 1811 3841 1823
rect 2197 1700 2249 1752
rect 2261 1700 2313 1752
rect 3097 1700 3149 1752
rect 3161 1700 3213 1752
rect 3789 1785 3841 1799
rect 3789 1751 3801 1785
rect 3801 1751 3835 1785
rect 3835 1751 3841 1785
rect 3878 1773 3930 1825
rect 3942 1773 3994 1825
rect 3789 1747 3841 1751
rect 1735 1494 1787 1546
rect 1735 1430 1787 1482
rect 793 1224 845 1276
rect 793 1160 845 1212
rect 1735 1224 1787 1276
rect 1735 1160 1787 1212
rect 3964 1567 4016 1619
rect 4028 1606 4080 1619
rect 4028 1572 4046 1606
rect 4046 1572 4080 1606
rect 4028 1567 4080 1572
rect 2770 1494 2822 1546
rect 2770 1430 2822 1482
rect 2770 1224 2822 1276
rect 2770 1160 2822 1212
rect 3886 1526 3938 1538
rect 3886 1492 3890 1526
rect 3890 1492 3924 1526
rect 3924 1492 3938 1526
rect 3886 1486 3938 1492
rect 3950 1526 4002 1538
rect 3950 1492 3962 1526
rect 3962 1492 3996 1526
rect 3996 1492 4002 1526
rect 3950 1486 4002 1492
rect 3838 1398 3890 1450
rect 3902 1398 3954 1450
rect 3340 1357 3392 1366
rect 3340 1323 3346 1357
rect 3346 1323 3380 1357
rect 3380 1323 3392 1357
rect 3340 1314 3392 1323
rect 3406 1357 3458 1366
rect 3406 1323 3422 1357
rect 3422 1323 3456 1357
rect 3456 1323 3458 1357
rect 3406 1314 3458 1323
rect 3675 1314 3727 1366
rect 3739 1314 3791 1366
rect 3612 1255 3664 1264
rect 3612 1221 3618 1255
rect 3618 1221 3652 1255
rect 3652 1221 3664 1255
rect 3612 1212 3664 1221
rect 3678 1255 3730 1264
rect 3678 1221 3690 1255
rect 3690 1221 3724 1255
rect 3724 1221 3730 1255
rect 3678 1212 3730 1221
rect 3304 1011 3356 1063
rect 3368 1011 3420 1063
rect 20213 2226 20265 2232
rect 20213 2192 20222 2226
rect 20222 2192 20256 2226
rect 20256 2192 20265 2226
rect 20213 2180 20265 2192
rect 20213 2154 20265 2168
rect 17668 2061 17720 2113
rect 17738 2061 17790 2113
rect 18025 2061 18077 2113
rect 18095 2061 18147 2113
rect 18424 2101 18476 2153
rect 18488 2101 18540 2153
rect 18884 2100 18936 2152
rect 18948 2100 19000 2152
rect 19640 2100 19692 2152
rect 19704 2100 19756 2152
rect 20213 2120 20222 2154
rect 20222 2120 20256 2154
rect 20256 2120 20265 2154
rect 22903 2267 22955 2273
rect 22903 2233 22909 2267
rect 22909 2233 22943 2267
rect 22943 2233 22955 2267
rect 22903 2221 22955 2233
rect 22903 2195 22955 2207
rect 22903 2161 22909 2195
rect 22909 2161 22943 2195
rect 22943 2161 22955 2195
rect 22903 2155 22955 2161
rect 23084 2255 23136 2261
rect 23084 2221 23093 2255
rect 23093 2221 23127 2255
rect 23127 2221 23136 2255
rect 23084 2209 23136 2221
rect 23084 2183 23136 2195
rect 23084 2149 23093 2183
rect 23093 2149 23127 2183
rect 23127 2149 23136 2183
rect 23084 2143 23136 2149
rect 20213 2116 20265 2120
rect 20507 2058 20559 2110
rect 20571 2058 20623 2110
rect 20975 2058 21027 2110
rect 21039 2058 21091 2110
rect 18715 2001 18767 2053
rect 18715 1937 18767 1989
rect 4528 1872 4580 1924
rect 4592 1872 4644 1924
rect 4727 1780 4779 1832
rect 4560 1700 4612 1752
rect 4624 1700 4676 1752
rect 4494 1490 4546 1542
rect 4558 1490 4610 1542
rect 4485 1392 4537 1444
rect 4327 1314 4379 1366
rect 4391 1314 4443 1366
rect 3872 951 3924 1003
rect 3938 951 3990 1003
rect 1295 293 1347 345
rect 1295 229 1347 281
rect 3454 827 3506 833
rect 3454 793 3461 827
rect 3461 793 3495 827
rect 3495 793 3506 827
rect 3454 781 3506 793
rect 3454 755 3506 767
rect 3454 721 3461 755
rect 3461 721 3495 755
rect 3495 721 3506 755
rect 3454 715 3506 721
rect 3870 871 3922 923
rect 3934 871 3986 923
rect 4305 1226 4357 1278
rect 4305 1162 4357 1214
rect 4041 787 4093 839
rect 4107 787 4159 839
rect 3512 443 3564 495
rect 3576 443 3628 495
rect 3852 661 3904 668
rect 3852 627 3858 661
rect 3858 627 3892 661
rect 3892 627 3904 661
rect 3852 616 3904 627
rect 3918 661 3970 668
rect 3918 627 3930 661
rect 3930 627 3964 661
rect 3964 627 3970 661
rect 3918 616 3970 627
rect 3370 261 3422 313
rect 3692 264 3744 316
rect 3756 264 3808 316
rect 3370 197 3422 249
rect 4305 174 4357 226
rect 2197 33 2249 85
rect 2299 33 2351 85
rect 3259 80 3311 132
rect 4305 110 4357 162
rect 3259 16 3311 68
rect 4396 93 4448 145
rect 4396 29 4448 81
rect 4485 1328 4537 1380
rect 4727 1716 4779 1768
rect 8202 1876 8254 1928
rect 8202 1812 8254 1864
rect 8202 1747 8254 1799
rect 8202 1682 8254 1734
rect 14441 1733 14493 1785
rect 14441 1669 14493 1721
rect 14447 1583 14499 1635
rect 14511 1583 14563 1635
rect 20746 1739 20798 1791
rect 20810 1739 20862 1791
rect 22853 1672 22905 1678
rect 21771 1614 21823 1666
rect 21771 1576 21823 1594
rect 22154 1648 22206 1655
rect 22154 1614 22163 1648
rect 22163 1614 22197 1648
rect 22197 1614 22206 1648
rect 22154 1603 22206 1614
rect 21771 1542 21780 1576
rect 21780 1542 21814 1576
rect 21814 1542 21823 1576
rect 22154 1576 22206 1583
rect 22154 1542 22163 1576
rect 22163 1542 22197 1576
rect 22197 1542 22206 1576
rect 22853 1638 22865 1672
rect 22865 1638 22899 1672
rect 22899 1638 22905 1672
rect 22853 1626 22905 1638
rect 22853 1600 22905 1612
rect 22853 1566 22865 1600
rect 22865 1566 22899 1600
rect 22899 1566 22905 1600
rect 22853 1560 22905 1566
rect 22154 1531 22206 1542
rect 23230 1533 23282 1585
rect 23294 1533 23346 1585
rect 22950 1466 23002 1470
rect 18230 1317 18282 1369
rect 22950 1432 22956 1466
rect 22956 1432 22990 1466
rect 22990 1432 23002 1466
rect 22950 1418 23002 1432
rect 22950 1394 23002 1406
rect 22950 1360 22956 1394
rect 22956 1360 22990 1394
rect 22990 1360 23002 1394
rect 22950 1354 23002 1360
rect 23327 1421 23379 1473
rect 23327 1357 23379 1409
rect 18230 1253 18282 1305
rect 18326 1270 18378 1322
rect 18326 1206 18378 1258
rect 17668 1146 17720 1198
rect 17738 1146 17790 1198
rect 18025 1145 18077 1197
rect 18095 1145 18147 1197
rect 18852 1105 18904 1157
rect 18916 1105 18968 1157
rect 21726 1025 21778 1077
rect 21804 1025 21856 1077
rect 5466 871 5518 923
rect 5530 871 5582 923
rect 6637 871 6689 923
rect 6703 871 6755 923
rect 18553 916 18605 968
rect 18617 916 18669 968
rect 22543 954 22595 1006
rect 4733 703 4785 755
rect 4797 703 4849 755
rect 4658 616 4710 668
rect 4722 616 4774 668
rect 4575 264 4627 316
rect 4639 264 4691 316
rect 4491 10 4543 62
rect 4555 10 4607 62
rect 5333 787 5385 839
rect 5399 787 5451 839
rect 5216 616 5268 668
rect 5282 616 5334 668
rect 6498 787 6550 839
rect 6564 787 6616 839
rect 6246 703 6298 755
rect 6312 703 6364 755
rect 6199 343 6251 395
rect 6199 270 6251 322
rect 6380 512 6432 521
rect 6380 478 6386 512
rect 6386 478 6420 512
rect 6420 478 6432 512
rect 6380 469 6432 478
rect 6446 512 6498 521
rect 6446 478 6458 512
rect 6458 478 6492 512
rect 6492 478 6498 512
rect 6446 469 6498 478
rect 22543 890 22595 942
rect 6766 512 6818 521
rect 6766 478 6772 512
rect 6772 478 6806 512
rect 6806 478 6818 512
rect 6766 469 6818 478
rect 6832 512 6884 521
rect 6832 478 6856 512
rect 6856 478 6884 512
rect 6832 469 6884 478
rect 6630 180 6682 232
rect 6694 180 6746 232
rect 7107 135 7159 144
rect 7107 101 7113 135
rect 7113 101 7147 135
rect 7147 101 7159 135
rect 7107 92 7159 101
rect 7171 135 7223 144
rect 7171 101 7185 135
rect 7185 101 7219 135
rect 7219 101 7223 135
rect 7171 92 7223 101
rect 6794 10 6846 62
rect 6860 10 6912 62
rect 21570 825 21622 877
rect 17635 758 17687 810
rect 17699 758 17751 810
rect 17956 750 18008 802
rect 18020 750 18072 802
rect 18741 738 18793 790
rect 18805 738 18857 790
rect 21570 761 21622 813
rect 21652 825 21704 877
rect 22693 869 22745 921
rect 21652 761 21704 813
rect 22693 805 22745 857
rect 15905 580 15957 587
rect 15905 546 15914 580
rect 15914 546 15948 580
rect 15948 546 15957 580
rect 15905 535 15957 546
rect 16961 580 17013 587
rect 16961 546 16970 580
rect 16970 546 17004 580
rect 17004 546 17013 580
rect 16961 535 17013 546
rect 15905 508 15957 520
rect 15905 474 15914 508
rect 15914 474 15948 508
rect 15948 474 15957 508
rect 15905 468 15957 474
rect 15992 511 16044 517
rect 15992 477 16001 511
rect 16001 477 16035 511
rect 16035 477 16044 511
rect 16257 511 16309 517
rect 15992 465 16044 477
rect 15992 439 16044 451
rect 15992 405 16001 439
rect 16001 405 16035 439
rect 16035 405 16044 439
rect 15992 399 16044 405
rect 16162 409 16214 431
rect 16162 379 16171 409
rect 16171 379 16205 409
rect 16205 379 16214 409
rect 16257 477 16266 511
rect 16266 477 16300 511
rect 16300 477 16309 511
rect 16961 508 17013 520
rect 16257 465 16309 477
rect 16257 439 16309 451
rect 16257 405 16266 439
rect 16266 405 16300 439
rect 16300 405 16309 439
rect 16257 399 16309 405
rect 16162 315 16214 367
rect 16609 481 16661 487
rect 16609 447 16618 481
rect 16618 447 16652 481
rect 16652 447 16661 481
rect 16609 435 16661 447
rect 16609 409 16661 421
rect 16609 375 16618 409
rect 16618 375 16652 409
rect 16652 375 16661 409
rect 16609 369 16661 375
rect 16874 481 16926 487
rect 16874 447 16883 481
rect 16883 447 16917 481
rect 16917 447 16926 481
rect 16961 474 16970 508
rect 16970 474 17004 508
rect 17004 474 17013 508
rect 16961 468 17013 474
rect 18132 516 18184 568
rect 18196 516 18248 568
rect 19254 577 19306 629
rect 19318 577 19370 629
rect 21718 560 21770 612
rect 21810 560 21862 612
rect 18296 454 18348 506
rect 18360 454 18412 506
rect 19254 474 19306 526
rect 19318 474 19370 526
rect 16874 435 16926 447
rect 16874 409 16926 421
rect 16874 375 16883 409
rect 16883 375 16917 409
rect 16917 375 16926 409
rect 16874 369 16926 375
rect 16516 228 16568 280
rect 17392 278 17444 330
rect 17456 278 17508 330
rect 20746 308 20862 488
rect 21718 471 21770 523
rect 21810 471 21862 523
rect 22087 427 22139 479
rect 22087 363 22139 415
rect 16516 164 16568 216
rect 20135 207 20187 259
rect 20199 207 20251 259
rect 17477 121 17529 173
rect 17477 57 17529 109
rect 19973 123 20025 175
rect 20037 123 20089 175
rect 18461 -102 18513 -50
rect 18525 -102 18577 -50
rect 18757 -114 18809 -62
rect 18821 -114 18873 -62
rect 18586 -201 18638 -149
rect 18650 -201 18702 -149
rect 4822 -414 4874 -362
rect 4886 -414 4938 -362
<< metal2 >>
tri 16319 3122 16322 3125 se
rect 16322 3122 18684 3125
tri 18684 3122 18687 3125 sw
rect 52 3070 58 3122
rect 110 3070 122 3122
rect 174 3117 180 3122
tri 16314 3117 16319 3122 se
rect 16319 3117 18687 3122
rect 174 3114 18687 3117
tri 18687 3114 18695 3122 sw
rect 174 3093 18695 3114
rect 174 3085 16377 3093
tri 16377 3085 16385 3093 nw
tri 18640 3085 18648 3093 ne
rect 18648 3085 18695 3093
rect 174 3070 180 3085
tri 180 3070 195 3085 nw
tri 18648 3070 18663 3085 ne
rect 18663 3070 18695 3085
tri 18695 3070 18739 3114 sw
tri 18663 3065 18668 3070 ne
rect 18668 3065 18739 3070
tri 18739 3065 18744 3070 sw
tri 16427 3057 16435 3065 se
rect 16435 3057 18495 3065
tri 204 3038 223 3057 se
rect 223 3038 18495 3057
rect 108 2986 114 3038
rect 166 2986 178 3038
rect 230 3035 18495 3038
rect 230 3022 16465 3035
tri 16465 3022 16478 3035 nw
rect 230 3013 262 3022
tri 262 3013 271 3022 nw
rect 18489 3013 18495 3035
rect 18547 3013 18567 3065
rect 18619 3013 18625 3065
tri 18668 3062 18671 3065 ne
rect 18671 3062 18744 3065
tri 18744 3062 18747 3065 sw
rect 21677 3062 21683 3114
rect 21735 3062 21755 3114
rect 21807 3093 22017 3114
tri 22017 3093 22038 3114 sw
rect 21807 3070 22038 3093
tri 22038 3070 22061 3093 sw
rect 21807 3065 22061 3070
tri 22061 3065 22066 3070 sw
rect 21807 3062 22066 3065
tri 18671 3056 18677 3062 ne
rect 18677 3056 18747 3062
tri 18747 3056 18753 3062 sw
tri 18677 3049 18684 3056 ne
rect 18684 3049 18753 3056
tri 18684 3035 18698 3049 ne
rect 18698 3035 18753 3049
tri 18698 3032 18701 3035 ne
rect 230 3005 254 3013
tri 254 3005 262 3013 nw
rect 230 2992 241 3005
tri 241 2992 254 3005 nw
tri 16547 2992 16560 3005 se
rect 16560 2992 18425 3005
rect 230 2986 236 2992
tri 236 2987 241 2992 nw
tri 310 2987 315 2992 se
rect 315 2987 18425 2992
tri 309 2986 310 2987 se
rect 310 2986 18425 2987
tri 18425 2986 18444 3005 sw
tri 304 2981 309 2986 se
rect 309 2981 18444 2986
tri 18444 2981 18449 2986 sw
tri 300 2977 304 2981 se
rect 304 2977 18449 2981
tri 290 2967 300 2977 se
rect 300 2976 18449 2977
rect 300 2975 18102 2976
tri 18102 2975 18103 2976 nw
tri 18364 2975 18365 2976 ne
rect 18365 2975 18449 2976
rect 300 2967 16592 2975
tri 16592 2967 16600 2975 nw
tri 18365 2967 18373 2975 ne
rect 18373 2967 18449 2975
tri 273 2950 290 2967 se
rect 290 2958 16583 2967
tri 16583 2958 16592 2967 nw
tri 18373 2958 18382 2967 ne
rect 18382 2958 18449 2967
rect 290 2950 344 2958
tri 344 2950 352 2958 nw
tri 18382 2950 18390 2958 ne
rect 18390 2950 18449 2958
rect 164 2898 170 2950
rect 222 2898 234 2950
rect 286 2946 340 2950
tri 340 2946 344 2950 nw
tri 18390 2946 18394 2950 ne
rect 18394 2946 18449 2950
rect 286 2928 322 2946
tri 322 2928 340 2946 nw
rect 16789 2928 16795 2946
rect 286 2898 292 2928
tri 292 2898 322 2928 nw
tri 345 2898 375 2928 se
rect 375 2898 16795 2928
tri 341 2894 345 2898 se
rect 345 2894 16795 2898
rect 16847 2894 16867 2946
rect 16919 2928 16925 2946
tri 18394 2943 18397 2946 ne
rect 16919 2915 18276 2928
tri 18276 2915 18289 2928 sw
rect 16919 2907 18289 2915
tri 18289 2907 18297 2915 sw
rect 16919 2894 18297 2907
tri 18297 2894 18310 2907 sw
tri 315 2868 341 2894 se
rect 341 2868 401 2894
tri 401 2868 427 2894 nw
tri 18256 2868 18282 2894 ne
rect 18282 2868 18310 2894
tri 18310 2868 18336 2894 sw
rect 224 2864 397 2868
tri 397 2864 401 2868 nw
tri 18282 2866 18284 2868 ne
rect 18284 2866 18336 2868
rect 224 2862 349 2864
rect 276 2816 349 2862
tri 349 2816 397 2864 nw
rect 4995 2836 5168 2866
tri 18284 2864 18286 2866 ne
rect 18286 2864 18336 2866
tri 4995 2816 5015 2836 ne
rect 5015 2816 5146 2836
tri 5015 2814 5017 2816 ne
rect 5017 2814 5146 2816
tri 5146 2814 5168 2836 nw
rect 14452 2830 16806 2864
rect 14452 2816 14506 2830
tri 14506 2816 14520 2830 nw
tri 16782 2816 16796 2830 ne
rect 16796 2816 16806 2830
rect 224 2798 276 2810
rect 14452 2812 14502 2816
tri 14502 2812 14506 2816 nw
tri 16796 2812 16800 2816 ne
rect 16800 2812 16806 2816
rect 16858 2812 16878 2864
rect 16930 2812 16936 2864
tri 18286 2853 18297 2864 ne
rect 18297 2853 18336 2864
tri 18336 2853 18351 2868 sw
tri 18297 2851 18299 2853 ne
rect 224 2740 276 2746
rect 1226 2754 1232 2806
rect 1284 2754 1308 2806
rect 1360 2754 1383 2806
rect 1435 2754 1441 2806
tri 2503 2788 2513 2798 se
rect 2513 2788 4924 2798
tri 4924 2788 4934 2798 sw
tri 5214 2788 5224 2798 se
rect 5224 2788 7510 2798
tri 7510 2788 7520 2798 sw
tri 8016 2788 8026 2798 se
rect 8026 2788 9917 2798
rect 1226 2714 1441 2754
rect 2110 2736 2116 2788
rect 2168 2736 2180 2788
rect 2232 2786 4934 2788
tri 4934 2786 4936 2788 sw
tri 5212 2786 5214 2788 se
rect 5214 2786 7520 2788
tri 7520 2786 7522 2788 sw
tri 8014 2786 8016 2788 se
rect 8016 2786 9917 2788
rect 2232 2755 9917 2786
rect 2232 2748 2549 2755
tri 2549 2748 2556 2755 nw
rect 2232 2736 2537 2748
tri 2537 2736 2549 2748 nw
rect 1226 2662 1232 2714
rect 1284 2662 1308 2714
rect 1360 2662 1383 2714
rect 1435 2662 1441 2714
tri 2564 2706 2583 2725 se
rect 2583 2706 9839 2725
rect 2071 2700 9839 2706
rect 2123 2673 9839 2700
rect 2071 2636 2123 2648
rect 2071 2578 2123 2584
rect 2289 2637 2341 2643
rect 2341 2585 8589 2634
rect 2289 2582 8589 2585
rect 2289 2573 2341 2582
rect 8580 2578 8589 2582
rect 8645 2578 8669 2634
rect 8725 2578 8734 2634
tri 2602 2522 2630 2550 se
rect 2630 2541 8519 2550
rect 2630 2522 8463 2541
rect 2289 2515 2341 2521
tri 2595 2515 2602 2522 se
rect 2602 2515 8463 2522
tri 2592 2512 2595 2515 se
rect 2595 2512 8463 2515
rect 2377 2460 2383 2512
rect 2435 2460 2447 2512
rect 2499 2507 8463 2512
rect 2499 2505 3081 2507
tri 3081 2505 3083 2507 nw
tri 3539 2505 3541 2507 ne
rect 3541 2505 8463 2507
rect 2499 2498 3074 2505
tri 3074 2498 3081 2505 nw
tri 3541 2498 3548 2505 ne
rect 3548 2498 8463 2505
rect 2499 2471 2632 2498
tri 2632 2471 2659 2498 nw
rect 3154 2471 3206 2477
rect 2499 2460 2621 2471
tri 2621 2460 2632 2471 nw
rect 1143 2421 1392 2427
rect 1195 2369 1340 2421
rect 1143 2357 1392 2369
rect 1195 2305 1340 2357
rect 3154 2407 3206 2419
rect 3249 2415 3255 2467
rect 3307 2415 3319 2467
rect 3371 2458 8393 2467
rect 3371 2415 8337 2458
rect 3206 2378 8267 2387
rect 3206 2355 8211 2378
rect 3154 2349 8211 2355
tri 7739 2342 7746 2349 ne
rect 7746 2342 8211 2349
tri 7746 2335 7753 2342 ne
rect 7753 2335 8211 2342
rect 1143 2299 1392 2305
rect 8211 2298 8267 2322
rect 8337 2378 8393 2402
rect 8463 2461 8519 2485
rect 8463 2396 8519 2405
rect 8337 2313 8393 2322
rect 8211 2233 8267 2242
rect 8202 1928 8254 1934
rect 3958 1872 3964 1924
rect 4016 1872 4028 1924
rect 4080 1872 4528 1924
rect 4580 1872 4592 1924
rect 4644 1872 4650 1924
rect 3789 1863 3841 1869
rect 8202 1864 8254 1876
rect 4727 1832 4779 1838
rect 3789 1799 3841 1811
rect 1340 1724 1392 1730
tri 1322 1672 1340 1690 se
rect 2191 1700 2197 1752
rect 2249 1700 2261 1752
rect 2313 1700 3097 1752
rect 3149 1700 3161 1752
rect 3213 1747 3668 1752
tri 3668 1747 3673 1752 sw
rect 3872 1773 3878 1825
rect 3930 1773 3942 1825
rect 3994 1814 4000 1825
rect 3994 1782 4727 1814
rect 3994 1773 4000 1782
rect 4727 1768 4779 1780
rect 3213 1713 3673 1747
tri 3673 1713 3707 1747 sw
rect 3789 1745 3841 1747
rect 4554 1745 4560 1752
rect 3789 1713 4560 1745
rect 3213 1700 3707 1713
tri 3707 1700 3720 1713 sw
rect 4554 1700 4560 1713
rect 4612 1700 4624 1752
rect 4676 1700 4682 1752
rect 4727 1710 4779 1716
rect 8202 1799 8254 1812
rect 14452 1791 14493 2812
tri 14493 2803 14502 2812 nw
rect 17011 2783 17017 2800
tri 14524 2755 14552 2783 se
rect 14552 2755 17017 2783
rect 8202 1734 8254 1747
tri 3642 1691 3651 1700 ne
rect 3651 1691 3720 1700
tri 3720 1691 3729 1700 sw
tri 1392 1682 1401 1691 sw
tri 3651 1685 3657 1691 ne
rect 3657 1685 3729 1691
tri 3729 1685 3735 1691 sw
tri 3657 1682 3660 1685 ne
rect 3660 1682 4152 1685
tri 4152 1682 4155 1685 sw
rect 1392 1672 1401 1682
tri 1319 1669 1322 1672 se
rect 1322 1669 1401 1672
tri 1401 1669 1414 1682 sw
tri 3660 1678 3664 1682 ne
rect 3664 1678 4155 1682
tri 4155 1678 4159 1682 sw
tri 3664 1674 3668 1678 ne
rect 3668 1674 4159 1678
tri 3668 1669 3673 1674 ne
rect 3673 1669 4159 1674
tri 4159 1669 4168 1678 sw
tri 1316 1666 1319 1669 se
rect 1319 1666 1414 1669
tri 1414 1666 1417 1669 sw
tri 3673 1666 3676 1669 ne
rect 3676 1666 4168 1669
tri 4168 1666 4171 1669 sw
tri 1310 1660 1316 1666 se
rect 1316 1663 1417 1666
tri 1417 1663 1420 1666 sw
tri 3676 1663 3679 1666 ne
rect 3679 1663 4171 1666
tri 4171 1663 4174 1666 sw
rect 1316 1660 1420 1663
tri 1304 1654 1310 1660 se
rect 1310 1654 1340 1660
rect -237 1608 1340 1654
rect 1392 1654 1420 1660
tri 1420 1654 1429 1663 sw
tri 3679 1654 3688 1663 ne
rect 3688 1654 4174 1663
tri 4174 1654 4183 1663 sw
rect 1392 1651 3382 1654
tri 3382 1651 3385 1654 sw
tri 3688 1651 3691 1654 ne
rect 3691 1651 4183 1654
tri 4183 1651 4186 1654 sw
rect 1392 1635 3385 1651
tri 3385 1635 3401 1651 sw
tri 3691 1647 3695 1651 ne
rect 3695 1647 4186 1651
tri 4129 1635 4141 1647 ne
rect 4141 1635 4186 1647
tri 4186 1635 4202 1651 sw
rect 1392 1619 3401 1635
tri 3401 1619 3417 1635 sw
tri 4141 1619 4157 1635 ne
rect 4157 1619 4202 1635
tri 4202 1619 4218 1635 sw
rect 1392 1608 3964 1619
rect -237 1602 3964 1608
tri 3348 1568 3382 1602 ne
rect 3382 1567 3964 1602
rect 4016 1567 4028 1619
rect 4080 1567 4086 1619
tri 4157 1617 4159 1619 ne
rect 4159 1617 4218 1619
tri 4218 1617 4220 1619 sw
tri 4159 1593 4183 1617 ne
rect 4183 1593 5355 1617
tri 5355 1593 5379 1617 sw
rect 8202 1593 8254 1682
rect 14441 1785 14493 1791
rect 14441 1721 14493 1733
rect 14441 1663 14493 1669
tri 14523 2754 14524 2755 se
rect 14524 2754 17017 2755
rect 14523 2749 17017 2754
rect 14523 2748 14591 2749
tri 14591 2748 14592 2749 nw
rect 17011 2748 17017 2749
rect 17069 2748 17089 2800
rect 17141 2748 17147 2800
rect 17309 2763 17315 2815
rect 17367 2763 17387 2815
rect 17439 2763 17459 2815
rect 17511 2763 17531 2815
rect 17583 2763 17602 2815
rect 17654 2763 17673 2815
rect 17725 2763 17744 2815
rect 17796 2763 17802 2815
rect 17309 2751 17802 2763
rect 14523 2736 14579 2748
tri 14579 2736 14591 2748 nw
rect 14523 2725 14568 2736
tri 14568 2725 14579 2736 nw
tri 14507 1635 14523 1651 se
rect 14523 1635 14556 2725
tri 14556 2713 14568 2725 nw
rect 17309 2699 17315 2751
rect 17367 2699 17387 2751
rect 17439 2699 17459 2751
rect 17511 2699 17531 2751
rect 17583 2699 17602 2751
rect 17654 2699 17673 2751
rect 17725 2699 17744 2751
rect 17796 2699 17802 2751
rect 17854 2719 17863 2775
rect 17919 2719 17944 2775
rect 18000 2719 18025 2775
rect 18081 2719 18105 2775
rect 18161 2719 18185 2775
rect 18241 2719 18250 2775
tri 17882 2680 17901 2699 ne
rect 17901 2680 18073 2699
tri 18073 2680 18092 2699 nw
tri 17901 2670 17911 2680 ne
rect 17911 2670 18063 2680
tri 18063 2670 18073 2680 nw
tri 17911 2658 17923 2670 ne
tri 18051 2658 18063 2670 nw
tri 17395 2453 17447 2505 se
rect 17447 2453 17633 2505
rect 17685 2453 17699 2505
rect 17751 2453 17757 2505
tri 17372 2430 17395 2453 se
rect 17395 2430 17420 2453
tri 17420 2430 17443 2453 nw
rect 17808 2430 17814 2482
rect 17866 2430 17880 2482
rect 17932 2430 17938 2482
tri 18276 2430 18299 2453 se
rect 18299 2431 18351 2853
rect 18299 2430 18339 2431
tri 17366 2424 17372 2430 se
rect 17372 2424 17414 2430
tri 17414 2424 17420 2430 nw
tri 17802 2424 17808 2430 se
rect 17808 2424 17880 2430
rect 17366 2419 17409 2424
tri 17409 2419 17414 2424 nw
tri 17797 2419 17802 2424 se
rect 17802 2419 17880 2424
tri 17880 2419 17891 2430 nw
tri 18265 2419 18276 2430 se
rect 18276 2419 18339 2430
tri 18339 2419 18351 2431 nw
tri 14556 1635 14569 1648 sw
tri 4183 1583 4193 1593 ne
rect 4193 1583 8254 1593
rect 14441 1583 14447 1635
rect 14499 1583 14511 1635
rect 14563 1583 14569 1635
tri 4193 1579 4197 1583 ne
rect 4197 1579 8254 1583
tri 5323 1567 5335 1579 ne
rect 5335 1567 8254 1579
tri 5335 1556 5346 1567 ne
rect 5346 1556 8254 1567
rect 793 1546 2822 1552
rect 845 1494 1735 1546
rect 1787 1494 2770 1546
rect 4488 1538 4494 1542
rect 793 1482 2822 1494
rect 3880 1486 3886 1538
rect 3938 1486 3950 1538
rect 4002 1503 4494 1538
rect 4002 1486 4008 1503
rect 4488 1490 4494 1503
rect 4546 1490 4558 1542
rect 4610 1490 4616 1542
rect 845 1430 1735 1482
rect 1787 1430 2770 1482
rect 793 1424 2822 1430
rect 3832 1398 3838 1450
rect 3890 1398 3902 1450
rect 3954 1444 4537 1450
rect 3954 1398 4485 1444
rect 4485 1380 4537 1392
rect 317 1314 3340 1366
rect 3392 1314 3406 1366
rect 3458 1314 3675 1366
rect 3727 1314 3739 1366
rect 3791 1314 4327 1366
rect 4379 1314 4391 1366
rect 4443 1314 4449 1366
rect 4485 1322 4537 1328
tri 4303 1282 4305 1284 se
rect 4305 1282 4357 1284
rect 793 1276 2822 1282
tri 4299 1278 4303 1282 se
rect 4303 1278 4357 1282
rect 845 1224 1735 1276
rect 1787 1224 2770 1276
tri 4285 1264 4299 1278 se
rect 4299 1264 4305 1278
rect 793 1212 2822 1224
rect 3606 1212 3612 1264
rect 3664 1212 3678 1264
rect 3730 1226 4305 1264
rect 17366 1243 17401 2419
tri 17401 2411 17409 2419 nw
tri 17789 2411 17797 2419 se
rect 17797 2411 17872 2419
tri 17872 2411 17880 2419 nw
tri 18257 2411 18265 2419 se
rect 18265 2411 18304 2419
tri 17473 2396 17488 2411 se
rect 17488 2396 17857 2411
tri 17857 2396 17872 2411 nw
tri 18242 2396 18257 2411 se
rect 18257 2396 18304 2411
tri 17444 2367 17473 2396 se
rect 17473 2376 17837 2396
tri 17837 2376 17857 2396 nw
tri 18230 2384 18242 2396 se
rect 18242 2384 18304 2396
tri 18304 2384 18339 2419 nw
rect 17473 2367 17492 2376
tri 17492 2367 17501 2376 nw
rect 18230 2367 18287 2384
tri 18287 2367 18304 2384 nw
tri 18394 2367 18397 2370 se
rect 18397 2367 18449 2946
tri 17440 2363 17444 2367 se
rect 17444 2363 17488 2367
tri 17488 2363 17492 2367 nw
rect 3730 1214 4357 1226
rect 3730 1212 4305 1214
rect 845 1160 1735 1212
rect 1787 1160 2770 1212
tri 4285 1192 4305 1212 ne
rect 793 1154 2822 1160
rect 4305 1156 4357 1162
rect 17125 1208 17401 1243
tri 17431 2354 17440 2363 se
rect 17440 2354 17479 2363
tri 17479 2354 17488 2363 nw
rect 17431 2342 17467 2354
tri 17467 2342 17479 2354 nw
rect 3298 1011 3304 1063
rect 3356 1011 3368 1063
rect 3420 1011 3426 1063
rect 3866 951 3872 1003
rect 3924 951 3938 1003
rect 3990 1000 6069 1003
tri 6069 1000 6072 1003 sw
rect 3990 968 6072 1000
tri 6072 968 6104 1000 sw
rect 3990 951 6104 968
tri 6044 923 6072 951 ne
rect 6072 923 6104 951
tri 6104 923 6149 968 sw
rect 3864 871 3870 923
rect 3922 871 3934 923
rect 3986 871 3992 923
rect 5460 871 5466 923
rect 5518 871 5530 923
rect 5582 871 5588 923
tri 6072 871 6124 923 ne
rect 6124 871 6637 923
rect 6689 871 6703 923
rect 6755 871 8168 923
rect 3454 833 3506 839
rect 4035 787 4041 839
rect 4093 787 4107 839
rect 4159 787 5333 839
rect 5385 787 5399 839
rect 5451 787 6498 839
rect 6550 787 6564 839
rect 6616 787 8350 839
rect 15675 787 16983 806
tri 16983 787 17002 806 sw
rect 3454 767 3506 781
rect 15675 776 17002 787
tri 17002 776 17013 787 sw
rect 15675 772 17013 776
tri 16939 758 16953 772 ne
rect 16953 758 17013 772
tri 16953 755 16956 758 ne
rect 16956 755 17013 758
rect 3506 715 4733 755
rect 3454 703 4733 715
rect 4785 703 4797 755
rect 4849 703 6246 755
rect 6298 703 6312 755
rect 6364 703 8150 755
tri 16956 750 16961 755 ne
rect 15673 738 15931 742
tri 15931 738 15935 742 sw
rect 15673 716 15935 738
tri 15935 716 15957 738 sw
rect 15673 708 15957 716
tri 15877 703 15882 708 ne
rect 15882 703 15957 708
tri 15882 680 15905 703 ne
rect 3846 616 3852 668
rect 3904 616 3918 668
rect 3970 616 4658 668
rect 4710 616 4722 668
rect 4774 616 5216 668
rect 5268 616 5282 668
rect 5334 616 5340 668
rect 15905 587 15957 703
rect 3506 443 3512 495
rect 3564 443 3576 495
rect 3628 443 3634 495
rect 6374 469 6380 521
rect 6432 469 6446 521
rect 6498 469 6766 521
rect 6818 469 6832 521
rect 6884 469 6890 521
rect 15905 520 15957 535
rect 16961 587 17013 755
rect 15905 462 15957 468
rect 15992 517 16309 523
rect 16044 488 16257 517
tri 16044 467 16065 488 nw
tri 16235 467 16256 488 ne
rect 16256 467 16257 488
tri 16256 466 16257 467 ne
rect 15992 451 16044 465
rect 6199 395 6251 401
rect 1295 345 1347 351
rect 16961 520 17013 535
rect 16257 451 16309 465
rect 15992 393 16044 399
rect 16162 431 16214 437
rect 16257 393 16309 399
rect 16609 487 16926 493
rect 16661 458 16874 487
rect 16661 437 16662 458
tri 16662 437 16683 458 nw
tri 16853 437 16874 458 ne
tri 16661 436 16662 437 nw
rect 16609 421 16661 435
tri 16156 369 16162 375 se
rect 16162 369 16214 379
tri 16154 367 16156 369 se
rect 16156 367 16214 369
tri 16132 345 16154 367 se
rect 16154 345 16162 367
rect 6199 322 6251 343
rect 1347 313 3422 319
rect 1347 293 3370 313
rect 1295 281 3370 293
rect 1347 266 3370 281
rect 1295 223 1347 229
rect 3686 264 3692 316
rect 3744 264 3756 316
rect 3808 264 4575 316
rect 4627 264 4639 316
rect 4691 270 6199 316
rect 15681 315 16162 345
rect 16609 363 16661 369
rect 16961 462 17013 468
rect 16874 421 16926 435
rect 16874 363 16926 369
rect 15681 309 16214 315
rect 4691 264 6251 270
rect 16516 280 16568 286
rect 3370 249 3422 261
rect 3370 191 3422 197
rect 4305 226 6630 232
rect 4357 180 6630 226
rect 6682 180 6694 232
rect 6746 180 8166 232
tri 16508 216 16516 224 se
rect 16516 216 16568 228
tri 16486 194 16508 216 se
rect 16508 194 16516 216
rect 4305 162 4357 174
rect 3259 132 3311 138
rect 2191 33 2197 85
rect 2249 33 2299 85
rect 2351 33 2357 85
rect 2191 16 2357 33
rect 15681 164 16516 194
rect 15681 158 16568 164
rect 4305 104 4357 110
rect 4396 145 4448 151
rect 3259 68 3311 80
tri 2357 16 2362 21 sw
rect 4448 93 7107 144
rect 4396 92 7107 93
rect 7159 92 7171 144
rect 7223 92 7231 144
tri 7779 121 7795 137 se
rect 7795 121 8153 137
tri 7767 109 7779 121 se
rect 7779 109 8153 121
tri 7750 92 7767 109 se
rect 7767 101 8153 109
rect 7767 92 7795 101
rect 4396 81 4448 92
tri 7725 67 7750 92 se
rect 7750 67 7795 92
tri 7795 67 7829 101 nw
tri 7720 62 7725 67 se
rect 7725 62 7790 67
tri 7790 62 7795 67 nw
rect 4396 23 4448 29
rect 2191 10 2362 16
tri 2362 10 2368 16 sw
rect 3259 10 3311 16
tri 3311 10 3315 14 sw
rect 4485 10 4491 62
rect 4543 10 4555 62
rect 4607 10 6794 62
rect 6846 10 6860 62
rect 6912 57 7785 62
tri 7785 57 7790 62 nw
rect 8589 60 8645 69
rect 6912 10 7738 57
tri 7738 10 7785 57 nw
rect 2191 6 2368 10
tri 2368 6 2372 10 sw
tri 3255 6 3259 10 se
rect 3259 6 3315 10
tri 2162 -23 2191 6 se
rect 2191 -23 2372 6
tri 2372 -23 2401 6 sw
tri 3226 -23 3255 6 se
rect 3255 -23 3315 6
tri 3315 -23 3348 10 sw
rect 2162 -74 3348 -23
rect 8589 -20 8645 4
rect 8211 -55 8267 -46
rect 8211 -135 8267 -111
rect 8211 -269 8267 -191
rect 8337 -54 8393 -45
rect 8337 -134 8393 -110
rect 8337 -197 8393 -190
rect 8463 -52 8519 -43
rect 8463 -132 8519 -108
rect 17125 -36 17160 1208
rect 17431 1178 17466 2342
tri 17466 2341 17467 2342 nw
rect 17662 2061 17668 2113
rect 17720 2061 17738 2113
rect 17790 2061 17796 2113
tri 17881 2061 17933 2113 se
rect 17933 2061 18025 2113
rect 18077 2061 18095 2113
rect 18147 2061 18153 2113
rect 17703 1198 17751 2061
tri 17878 2058 17881 2061 se
rect 17881 2058 17947 2061
tri 17947 2058 17950 2061 nw
tri 17873 2053 17878 2058 se
rect 17878 2053 17942 2058
tri 17942 2053 17947 2058 nw
tri 17864 2044 17873 2053 se
rect 17873 2044 17933 2053
tri 17933 2044 17942 2053 nw
tri 17821 2001 17864 2044 se
rect 17864 2001 17890 2044
tri 17890 2001 17933 2044 nw
tri 17809 1989 17821 2001 se
rect 17821 1989 17878 2001
tri 17878 1989 17890 2001 nw
tri 17795 1975 17809 1989 se
rect 17809 1975 17864 1989
tri 17864 1975 17878 1989 nw
tri 17781 1961 17795 1975 se
rect 17795 1961 17850 1975
tri 17850 1961 17864 1975 nw
rect 17781 1335 17830 1961
tri 17830 1941 17850 1961 nw
rect 18230 1369 18282 2367
tri 18282 2362 18287 2367 nw
tri 18389 2362 18394 2367 se
rect 18394 2362 18449 2367
tri 18369 2342 18389 2362 se
rect 18389 2348 18449 2362
rect 18389 2343 18444 2348
tri 18444 2343 18449 2348 nw
rect 18389 2342 18443 2343
tri 18443 2342 18444 2343 nw
tri 18488 2342 18489 2343 se
rect 18489 2342 18541 3013
rect 18701 2453 18753 3035
tri 21995 3029 22028 3062 ne
rect 22028 3029 22066 3062
tri 22066 3029 22102 3065 sw
rect 21584 2977 21590 3029
rect 21642 2977 21662 3029
rect 21714 3019 21780 3029
tri 21780 3019 21790 3029 sw
tri 22028 3019 22038 3029 ne
rect 22038 3019 22102 3029
tri 22102 3019 22112 3029 sw
rect 21714 2983 21790 3019
tri 21790 2983 21826 3019 sw
rect 21714 2977 21826 2983
tri 22038 2977 22080 3019 ne
rect 22080 2977 22112 3019
tri 22112 2977 22154 3019 sw
tri 21750 2967 21760 2977 ne
rect 21760 2967 21826 2977
tri 22080 2967 22090 2977 ne
rect 22090 2967 22154 2977
tri 22154 2967 22164 2977 sw
rect 19542 2915 19548 2967
rect 19600 2915 19620 2967
rect 19672 2915 19756 2967
tri 19756 2915 19808 2967 sw
rect 19868 2915 19874 2967
rect 19926 2915 19946 2967
rect 19998 2965 20034 2967
tri 20034 2965 20036 2967 sw
tri 21760 2965 21762 2967 ne
rect 21762 2965 21826 2967
tri 22090 2965 22092 2967 ne
rect 22092 2965 22164 2967
tri 22164 2965 22166 2967 sw
rect 19998 2915 20036 2965
tri 20036 2915 20086 2965 sw
tri 21762 2959 21768 2965 ne
tri 19734 2841 19808 2915 ne
tri 19808 2841 19882 2915 sw
tri 20012 2891 20036 2915 ne
rect 20036 2913 20086 2915
tri 20086 2913 20088 2915 sw
tri 19808 2821 19828 2841 ne
rect 19828 2821 19882 2841
tri 19882 2821 19902 2841 sw
tri 19828 2767 19882 2821 ne
rect 19882 2767 19902 2821
tri 19902 2767 19956 2821 sw
rect 20036 2769 20088 2913
tri 20088 2769 20110 2791 sw
rect 20278 2779 20287 2835
rect 20343 2779 20368 2835
rect 20424 2779 20449 2835
tri 20036 2767 20038 2769 ne
rect 20038 2767 20110 2769
tri 19882 2742 19907 2767 ne
rect 19907 2742 19956 2767
tri 19956 2742 19981 2767 sw
tri 20038 2742 20063 2767 ne
rect 20063 2742 20110 2767
tri 20110 2742 20137 2769 sw
rect 20278 2755 20449 2779
tri 19907 2736 19913 2742 ne
rect 19913 2736 19981 2742
tri 19981 2736 19987 2742 sw
tri 20063 2736 20069 2742 ne
rect 20069 2736 20137 2742
tri 20137 2736 20143 2742 sw
tri 19913 2725 19924 2736 ne
rect 19924 2725 19987 2736
tri 19987 2725 19998 2736 sw
tri 20069 2725 20080 2736 ne
rect 20080 2725 20143 2736
tri 20143 2725 20154 2736 sw
tri 19924 2708 19941 2725 ne
rect 19941 2708 19998 2725
tri 19998 2708 20015 2725 sw
tri 20080 2708 20097 2725 ne
rect 20097 2708 20154 2725
tri 20154 2708 20171 2725 sw
tri 19941 2705 19944 2708 ne
rect 19944 2705 20015 2708
tri 20015 2705 20018 2708 sw
tri 20097 2705 20100 2708 ne
rect 20100 2705 20171 2708
tri 20171 2705 20174 2708 sw
tri 19944 2700 19949 2705 ne
rect 19949 2700 20018 2705
tri 20018 2700 20023 2705 sw
tri 20100 2700 20105 2705 ne
rect 20105 2700 20174 2705
tri 20174 2700 20179 2705 sw
tri 19949 2693 19956 2700 ne
rect 19956 2693 20023 2700
tri 20023 2693 20030 2700 sw
tri 20105 2695 20110 2700 ne
rect 20110 2695 20179 2700
tri 20179 2695 20184 2700 sw
rect 20278 2699 20287 2755
rect 20343 2699 20368 2755
rect 20424 2699 20449 2755
rect 20665 2827 20674 2835
tri 20674 2827 20682 2835 sw
rect 20665 2821 21159 2827
rect 20665 2705 20848 2821
rect 21156 2705 21159 2821
rect 21379 2764 21385 2816
rect 21437 2764 21449 2816
rect 21501 2764 21507 2816
tri 21391 2752 21403 2764 ne
rect 21403 2753 21485 2764
tri 21485 2753 21496 2764 nw
rect 21403 2752 21484 2753
tri 21484 2752 21485 2753 nw
tri 21403 2742 21413 2752 ne
rect 21413 2742 21474 2752
tri 21474 2742 21484 2752 nw
tri 21413 2736 21419 2742 ne
rect 21419 2740 21472 2742
tri 21472 2740 21474 2742 nw
rect 21419 2736 21468 2740
tri 21468 2736 21472 2740 nw
tri 21419 2730 21425 2736 ne
rect 20665 2699 21159 2705
tri 21421 2702 21425 2706 se
rect 21425 2702 21462 2736
tri 21462 2730 21468 2736 nw
tri 21591 2725 21592 2726 se
rect 21592 2725 21598 2752
tri 21574 2708 21591 2725 se
rect 21591 2708 21598 2725
tri 21568 2702 21574 2708 se
rect 21574 2702 21598 2708
tri 21419 2700 21421 2702 se
rect 21421 2700 21462 2702
tri 21566 2700 21568 2702 se
rect 21568 2700 21598 2702
rect 21650 2700 21662 2752
rect 21714 2700 21720 2752
tri 21418 2699 21419 2700 se
rect 21419 2699 21462 2700
tri 20563 2695 20567 2699 ne
rect 20567 2695 20755 2699
tri 20755 2695 20759 2699 nw
tri 21414 2695 21418 2699 se
rect 21418 2695 21462 2699
tri 21561 2695 21566 2700 se
rect 21566 2695 21611 2700
tri 21611 2695 21616 2700 nw
tri 20110 2693 20112 2695 ne
rect 20112 2693 20184 2695
tri 19956 2680 19969 2693 ne
rect 19969 2680 20030 2693
tri 20030 2680 20043 2693 sw
tri 20112 2680 20125 2693 ne
rect 20125 2680 20184 2693
tri 20184 2680 20199 2695 sw
tri 20567 2680 20582 2695 ne
rect 20582 2684 20744 2695
tri 20744 2684 20755 2695 nw
tri 21403 2684 21414 2695 se
rect 21414 2691 21462 2695
rect 21414 2684 21455 2691
tri 21455 2684 21462 2691 nw
tri 21550 2684 21561 2695 se
rect 21561 2684 21600 2695
tri 21600 2684 21611 2695 nw
rect 20582 2680 20740 2684
tri 20740 2680 20744 2684 nw
tri 21399 2680 21403 2684 se
rect 21403 2680 21451 2684
tri 21451 2680 21455 2684 nw
tri 21546 2680 21550 2684 se
rect 21550 2680 21596 2684
tri 21596 2680 21600 2684 nw
tri 19969 2673 19976 2680 ne
rect 19976 2673 20043 2680
tri 20043 2673 20050 2680 sw
tri 20125 2673 20132 2680 ne
rect 20132 2673 20199 2680
tri 20199 2673 20206 2680 sw
tri 20582 2673 20589 2680 ne
rect 20589 2673 20733 2680
tri 20733 2673 20740 2680 nw
tri 21392 2673 21399 2680 se
rect 21399 2673 21444 2680
tri 21444 2673 21451 2680 nw
tri 21539 2673 21546 2680 se
rect 21546 2673 21589 2680
tri 21589 2673 21596 2680 nw
tri 19976 2646 20003 2673 ne
rect 20003 2646 20050 2673
tri 20050 2646 20077 2673 sw
tri 20132 2646 20159 2673 ne
rect 20159 2646 20206 2673
tri 20206 2646 20233 2673 sw
tri 20589 2670 20592 2673 ne
rect 20592 2670 20730 2673
tri 20730 2670 20733 2673 nw
tri 21389 2670 21392 2673 se
rect 21392 2670 21425 2673
tri 20592 2665 20597 2670 ne
tri 20725 2665 20730 2670 nw
tri 21384 2665 21389 2670 se
rect 21389 2665 21425 2670
tri 21373 2654 21384 2665 se
rect 21384 2654 21425 2665
tri 21425 2654 21444 2673 nw
tri 21520 2654 21539 2673 se
rect 21539 2654 21562 2673
tri 21365 2646 21373 2654 se
rect 21373 2646 21417 2654
tri 21417 2646 21425 2654 nw
tri 21512 2646 21520 2654 se
rect 21520 2646 21562 2654
tri 21562 2646 21589 2673 nw
tri 20003 2619 20030 2646 ne
rect 20030 2619 20077 2646
tri 20077 2619 20104 2646 sw
tri 20159 2621 20184 2646 ne
rect 20184 2621 20496 2646
tri 20496 2621 20521 2646 sw
tri 21353 2634 21365 2646 se
rect 21365 2634 21405 2646
tri 21405 2634 21417 2646 nw
tri 21500 2634 21512 2646 se
rect 21512 2634 21550 2646
tri 21550 2634 21562 2646 nw
tri 21340 2621 21353 2634 se
rect 21353 2621 21392 2634
tri 21392 2621 21405 2634 nw
tri 21487 2621 21500 2634 se
rect 21500 2621 21537 2634
tri 21537 2621 21550 2634 nw
tri 20184 2619 20186 2621 ne
rect 20186 2619 20521 2621
tri 20030 2545 20104 2619 ne
tri 20104 2549 20174 2619 sw
tri 20186 2594 20211 2619 ne
rect 20211 2617 20521 2619
tri 20521 2617 20525 2621 sw
tri 21336 2617 21340 2621 se
rect 21340 2617 21388 2621
tri 21388 2617 21392 2621 nw
tri 21483 2617 21487 2621 se
rect 21487 2617 21533 2621
tri 21533 2617 21537 2621 nw
rect 20211 2594 20525 2617
tri 20525 2594 20548 2617 sw
tri 21321 2602 21336 2617 se
rect 21336 2602 21373 2617
tri 21373 2602 21388 2617 nw
tri 21468 2602 21483 2617 se
rect 21483 2602 21510 2617
tri 21313 2594 21321 2602 se
rect 21321 2594 21365 2602
tri 21365 2594 21373 2602 nw
tri 21460 2594 21468 2602 se
rect 21468 2594 21510 2602
tri 21510 2594 21533 2617 nw
tri 20474 2549 20519 2594 ne
rect 20519 2584 20548 2594
tri 20548 2584 20558 2594 sw
tri 21303 2584 21313 2594 se
rect 21313 2584 21355 2594
tri 21355 2584 21365 2594 nw
tri 21450 2584 21460 2594 se
rect 21460 2584 21500 2594
tri 21500 2584 21510 2594 nw
rect 20519 2550 20909 2584
tri 20909 2550 20943 2584 sw
tri 21269 2550 21303 2584 se
rect 21303 2550 21321 2584
tri 21321 2550 21355 2584 nw
tri 21416 2550 21450 2584 se
rect 20519 2549 20943 2550
rect 20104 2545 20460 2549
tri 20460 2545 20464 2549 sw
tri 20519 2545 20523 2549 ne
rect 20523 2545 20943 2549
tri 20104 2522 20127 2545 ne
rect 20127 2543 20464 2545
tri 20464 2543 20466 2545 sw
tri 20523 2543 20525 2545 ne
rect 20525 2543 20943 2545
rect 20127 2522 20466 2543
rect 18798 2470 18804 2522
rect 18856 2470 18868 2522
rect 18920 2470 18926 2522
tri 20127 2511 20138 2522 ne
rect 20138 2511 20466 2522
tri 20466 2511 20498 2543 sw
tri 20876 2528 20891 2543 ne
rect 20891 2511 20943 2543
tri 21253 2534 21269 2550 se
rect 21269 2534 21305 2550
tri 21305 2534 21321 2550 nw
tri 21400 2534 21416 2550 se
rect 21416 2534 21450 2550
tri 21450 2534 21500 2584 nw
tri 21230 2511 21253 2534 se
rect 21253 2511 21282 2534
tri 21282 2511 21305 2534 nw
tri 21377 2511 21400 2534 se
rect 21400 2511 21427 2534
tri 21427 2511 21450 2534 nw
tri 20138 2497 20152 2511 ne
rect 20152 2497 20716 2511
tri 20438 2470 20465 2497 ne
rect 20465 2470 20716 2497
rect 18798 2459 18876 2470
tri 20465 2464 20471 2470 ne
rect 20471 2464 20716 2470
tri 19426 2459 19431 2464 se
rect 19431 2459 20421 2464
tri 20421 2459 20426 2464 sw
tri 20471 2459 20476 2464 ne
rect 20476 2459 20716 2464
rect 20768 2459 20780 2511
rect 20832 2459 20838 2511
rect 20891 2459 20897 2511
rect 20949 2459 20961 2511
rect 21013 2459 21019 2511
tri 21217 2498 21230 2511 se
rect 21230 2498 21269 2511
tri 21269 2498 21282 2511 nw
tri 21364 2498 21377 2511 se
rect 21377 2498 21400 2511
tri 21203 2484 21217 2498 se
rect 21217 2484 21255 2498
tri 21255 2484 21269 2498 nw
tri 21350 2484 21364 2498 se
rect 21364 2484 21400 2498
tri 21400 2484 21427 2511 nw
tri 21178 2459 21203 2484 se
rect 21203 2459 21230 2484
tri 21230 2459 21255 2484 nw
tri 21325 2459 21350 2484 se
rect 21350 2459 21375 2484
tri 21375 2459 21400 2484 nw
tri 18798 2457 18800 2459 ne
rect 18800 2457 18876 2459
tri 18753 2453 18757 2457 sw
tri 18800 2453 18804 2457 ne
rect 18804 2453 18876 2457
tri 19420 2453 19426 2459 se
rect 19426 2453 20426 2459
tri 20426 2453 20432 2459 sw
tri 21172 2453 21178 2459 se
rect 21178 2453 21224 2459
tri 21224 2453 21230 2459 nw
tri 21319 2453 21325 2459 se
rect 21325 2453 21369 2459
tri 21369 2453 21375 2459 nw
rect 18701 2435 18757 2453
tri 18701 2427 18709 2435 ne
rect 18709 2433 18757 2435
tri 18757 2433 18777 2453 sw
tri 18804 2433 18824 2453 ne
rect 18709 2427 18777 2433
tri 18777 2427 18783 2433 sw
tri 18709 2419 18717 2427 ne
rect 18717 2419 18783 2427
tri 18717 2405 18731 2419 ne
tri 17830 1335 17851 1356 sw
tri 17781 1317 17799 1335 ne
rect 17799 1317 17851 1335
tri 17851 1317 17869 1335 sw
tri 17799 1305 17811 1317 ne
rect 17811 1305 17869 1317
tri 17869 1305 17881 1317 sw
rect 18230 1305 18282 1317
tri 17811 1265 17851 1305 ne
rect 17851 1265 17881 1305
tri 17881 1265 17921 1305 sw
tri 17851 1253 17863 1265 ne
rect 17863 1253 17921 1265
tri 17921 1253 17933 1265 sw
tri 17863 1241 17875 1253 ne
rect 17875 1241 17933 1253
tri 17933 1241 17945 1253 sw
rect 18230 1241 18282 1253
tri 18326 2299 18369 2342 se
rect 18369 2317 18418 2342
tri 18418 2317 18443 2342 nw
tri 18463 2317 18488 2342 se
rect 18488 2319 18541 2342
rect 18488 2317 18512 2319
rect 18369 2299 18400 2317
tri 18400 2299 18418 2317 nw
tri 18445 2299 18463 2317 se
rect 18463 2299 18512 2317
rect 18326 2290 18391 2299
tri 18391 2290 18400 2299 nw
tri 18436 2290 18445 2299 se
rect 18445 2290 18512 2299
tri 18512 2290 18541 2319 nw
rect 18575 2290 18581 2342
rect 18633 2290 18645 2342
rect 18697 2290 18703 2342
rect 18326 1322 18378 2290
tri 18378 2277 18391 2290 nw
tri 18423 2277 18436 2290 se
rect 18436 2277 18494 2290
tri 18418 2272 18423 2277 se
rect 18423 2272 18494 2277
tri 18494 2272 18512 2290 nw
rect 18418 2245 18467 2272
tri 18467 2245 18494 2272 nw
rect 18418 2153 18463 2245
tri 18463 2241 18467 2245 nw
rect 18418 2101 18424 2153
rect 18476 2101 18488 2153
rect 18540 2101 18546 2153
rect 18326 1258 18378 1270
tri 17875 1206 17910 1241 ne
rect 17910 1206 17945 1241
tri 17945 1206 17980 1241 sw
tri 17910 1200 17916 1206 ne
rect 17916 1200 17980 1206
tri 17980 1200 17986 1206 sw
rect 18326 1200 18378 1206
tri 17916 1198 17918 1200 ne
rect 17918 1198 17986 1200
tri 9561 -50 9575 -36 se
rect 9575 -50 17160 -36
tri 9540 -71 9561 -50 se
rect 9561 -71 17160 -50
rect 17188 1143 17466 1178
rect 17662 1146 17668 1198
rect 17720 1146 17738 1198
rect 17790 1165 17796 1198
tri 17918 1197 17919 1198 ne
rect 17919 1197 17986 1198
tri 17986 1197 17989 1200 sw
tri 17919 1195 17921 1197 ne
rect 17921 1195 18025 1197
tri 17921 1170 17946 1195 ne
rect 17946 1170 18025 1195
tri 17796 1165 17801 1170 sw
tri 17946 1165 17951 1170 ne
rect 17951 1165 18025 1170
rect 17790 1146 17801 1165
tri 17801 1146 17820 1165 sw
tri 17951 1146 17970 1165 ne
rect 17970 1146 18025 1165
tri 17752 1145 17753 1146 ne
rect 17753 1145 17820 1146
tri 17820 1145 17821 1146 sw
tri 17970 1145 17971 1146 ne
rect 17971 1145 18025 1146
rect 18077 1145 18095 1197
rect 18147 1157 18278 1197
tri 18278 1157 18318 1197 sw
rect 18147 1145 18318 1157
tri 18318 1145 18330 1157 sw
tri 17753 1143 17755 1145 ne
rect 17755 1143 17821 1145
tri 17821 1143 17823 1145 sw
tri 18245 1143 18247 1145 ne
rect 18247 1143 18330 1145
tri 18330 1143 18332 1145 sw
rect 8589 -85 8645 -76
tri 8645 -85 8659 -71 sw
tri 9526 -85 9540 -71 se
rect 9540 -85 9575 -71
rect 8589 -99 8659 -85
tri 8659 -99 8673 -85 sw
tri 9512 -99 9526 -85 se
rect 9526 -99 9575 -85
tri 9575 -99 9603 -71 nw
rect 8589 -101 8673 -99
tri 8673 -101 8675 -99 sw
tri 9510 -101 9512 -99 se
rect 9512 -101 9573 -99
tri 9573 -101 9575 -99 nw
rect 17188 -101 17223 1143
tri 17755 1105 17793 1143 ne
rect 17793 1133 17823 1143
tri 17823 1133 17833 1143 sw
tri 18247 1133 18257 1143 ne
rect 18257 1133 18332 1143
tri 18332 1133 18342 1143 sw
rect 17793 1112 17833 1133
tri 17833 1112 17854 1133 sw
tri 18257 1112 18278 1133 ne
rect 18278 1112 18342 1133
rect 17793 1105 17854 1112
tri 17854 1105 17861 1112 sw
tri 18278 1105 18285 1112 ne
rect 18285 1105 18342 1112
tri 17793 1097 17801 1105 ne
rect 17801 1100 17861 1105
tri 17861 1100 17866 1105 sw
tri 18285 1100 18290 1105 ne
rect 17801 1097 17866 1100
tri 17866 1097 17869 1100 sw
tri 17801 1090 17808 1097 ne
rect 17808 1090 18144 1097
tri 18144 1090 18151 1097 sw
tri 17808 1077 17821 1090 ne
rect 17821 1077 18151 1090
tri 18151 1077 18164 1090 sw
tri 17821 1049 17849 1077 ne
rect 17849 1049 18164 1077
tri 18124 1025 18148 1049 ne
rect 18148 1025 18164 1049
tri 18164 1025 18216 1077 sw
tri 18148 1022 18151 1025 ne
rect 18151 1022 18216 1025
tri 18216 1022 18219 1025 sw
tri 18151 1006 18167 1022 ne
rect 18167 1006 18219 1022
tri 18167 1002 18171 1006 ne
rect 17277 859 18078 894
rect 17277 553 17309 859
tri 17933 842 17950 859 ne
rect 17344 813 17407 814
tri 17407 813 17408 814 sw
rect 17344 810 17408 813
tri 17408 810 17411 813 sw
rect 17344 796 17411 810
tri 17411 796 17425 810 sw
tri 17599 796 17613 810 se
rect 17613 796 17635 810
rect 17344 793 17425 796
tri 17425 793 17428 796 sw
tri 17596 793 17599 796 se
rect 17599 793 17635 796
rect 17344 758 17635 793
rect 17687 758 17699 810
rect 17751 758 17757 810
rect 17950 802 18078 859
rect 17344 750 17410 758
tri 17410 750 17418 758 nw
rect 17950 750 17956 802
rect 18008 750 18020 802
rect 18072 750 18078 802
rect 17344 738 17398 750
tri 17398 738 17410 750 nw
rect 17344 668 17397 738
tri 17397 737 17398 738 nw
tri 17344 650 17362 668 ne
rect 8589 -102 8675 -101
tri 8675 -102 8676 -101 sw
tri 9509 -102 9510 -101 se
rect 9510 -102 9572 -101
tri 9572 -102 9573 -101 nw
tri 9618 -102 9619 -101 se
rect 9619 -102 17223 -101
rect 8589 -108 8676 -102
tri 8676 -108 8682 -102 sw
tri 9503 -108 9509 -102 se
rect 9509 -108 9566 -102
tri 9566 -108 9572 -102 nw
tri 9612 -108 9618 -102 se
rect 9618 -108 17223 -102
rect 8589 -114 9560 -108
tri 9560 -114 9566 -108 nw
tri 9606 -114 9612 -108 se
rect 9612 -114 17223 -108
rect 8589 -130 9544 -114
tri 9544 -130 9560 -114 nw
tri 9590 -130 9606 -114 se
rect 9606 -130 17223 -114
tri 8589 -135 8594 -130 ne
rect 8594 -135 9530 -130
tri 8519 -149 8533 -135 sw
tri 8594 -144 8603 -135 ne
rect 8603 -144 9530 -135
tri 9530 -144 9544 -130 nw
tri 9576 -144 9590 -130 se
rect 9590 -134 17223 -130
rect 17252 521 17309 553
rect 9590 -144 9634 -134
tri 9571 -149 9576 -144 se
rect 9576 -149 9634 -144
tri 9634 -149 9649 -134 nw
rect 8519 -163 8533 -149
tri 8533 -163 8547 -149 sw
tri 9557 -163 9571 -149 se
rect 9571 -163 9620 -149
tri 9620 -163 9634 -149 nw
rect 17252 -163 17284 521
rect 17362 481 17397 668
rect 18171 568 18219 1006
rect 18126 516 18132 568
rect 18184 516 18196 568
rect 18248 516 18254 568
rect 8519 -164 8547 -163
tri 8547 -164 8548 -163 sw
tri 9556 -164 9557 -163 se
rect 9557 -164 9619 -163
tri 9619 -164 9620 -163 nw
tri 9664 -164 9665 -163 se
rect 9665 -164 17284 -163
rect 8519 -173 8548 -164
tri 8548 -173 8557 -164 sw
tri 9547 -173 9556 -164 se
rect 9556 -173 9610 -164
tri 9610 -173 9619 -164 nw
tri 9655 -173 9664 -164 se
rect 9664 -173 17284 -164
rect 8519 -188 9586 -173
tri 8393 -197 8395 -195 sw
rect 8463 -197 9586 -188
tri 9586 -197 9610 -173 nw
tri 9631 -197 9655 -173 se
rect 9655 -196 17284 -173
rect 17313 446 17397 481
rect 18290 506 18342 1105
rect 18639 968 18675 2290
tri 18715 2252 18731 2268 se
rect 18731 2252 18783 2419
rect 18715 2246 18783 2252
rect 18715 2245 18782 2246
tri 18782 2245 18783 2246 nw
rect 18715 2232 18769 2245
tri 18769 2232 18782 2245 nw
rect 18715 2053 18767 2232
tri 18767 2230 18769 2232 nw
rect 18715 1989 18767 2001
rect 18715 1931 18767 1937
tri 18797 2202 18824 2229 se
rect 18824 2207 18876 2453
tri 19391 2424 19420 2453 se
rect 19420 2446 20432 2453
tri 20432 2446 20439 2453 sw
tri 21165 2446 21172 2453 se
rect 21172 2446 21217 2453
tri 21217 2446 21224 2453 nw
tri 21312 2446 21319 2453 se
rect 21319 2446 21350 2453
rect 19420 2434 20439 2446
tri 20439 2434 20451 2446 sw
tri 21153 2434 21165 2446 se
rect 21165 2434 21205 2446
tri 21205 2434 21217 2446 nw
tri 21300 2434 21312 2446 se
rect 21312 2434 21350 2446
tri 21350 2434 21369 2453 nw
rect 19420 2424 19439 2434
tri 19439 2424 19449 2434 nw
tri 20400 2424 20410 2434 ne
rect 20410 2424 20451 2434
tri 20451 2424 20461 2434 sw
tri 21143 2424 21153 2434 se
rect 21153 2424 21195 2434
tri 21195 2424 21205 2434 nw
tri 21290 2424 21300 2434 se
rect 21300 2424 21335 2434
tri 19386 2419 19391 2424 se
rect 19391 2419 19434 2424
tri 19434 2419 19439 2424 nw
tri 20410 2419 20415 2424 ne
rect 20415 2419 21190 2424
tri 21190 2419 21195 2424 nw
tri 21285 2419 21290 2424 se
rect 21290 2419 21335 2424
tri 21335 2419 21350 2434 nw
tri 19383 2416 19386 2419 se
rect 19386 2416 19431 2419
tri 19431 2416 19434 2419 nw
tri 20415 2416 20418 2419 ne
rect 20418 2416 21184 2419
tri 19371 2404 19383 2416 se
rect 19383 2404 19419 2416
tri 19419 2404 19431 2416 nw
tri 20418 2413 20421 2416 ne
rect 20421 2413 21184 2416
tri 21184 2413 21190 2419 nw
tri 21279 2413 21285 2419 se
rect 21285 2413 21300 2419
tri 20421 2404 20430 2413 ne
rect 20430 2404 21165 2413
tri 19351 2384 19371 2404 se
rect 19371 2384 19399 2404
tri 19399 2384 19419 2404 nw
tri 19464 2384 19484 2404 se
rect 19484 2384 20324 2404
tri 20324 2384 20344 2404 sw
tri 20430 2394 20440 2404 ne
rect 20440 2394 21165 2404
tri 21165 2394 21184 2413 nw
tri 21260 2394 21279 2413 se
rect 21279 2394 21300 2413
tri 21250 2384 21260 2394 se
rect 21260 2384 21300 2394
tri 21300 2384 21335 2419 nw
rect 18824 2202 18871 2207
tri 18871 2202 18876 2207 nw
tri 19346 2379 19351 2384 se
rect 19351 2379 19394 2384
tri 19394 2379 19399 2384 nw
tri 19459 2379 19464 2384 se
rect 19464 2379 20344 2384
rect 19346 2374 19389 2379
tri 19389 2374 19394 2379 nw
tri 19454 2374 19459 2379 se
rect 19459 2374 20344 2379
tri 20344 2374 20354 2384 sw
tri 21240 2374 21250 2384 se
rect 21250 2374 21290 2384
tri 21290 2374 21300 2384 nw
rect 19346 2367 19382 2374
tri 19382 2367 19389 2374 nw
tri 19447 2367 19454 2374 se
rect 19454 2367 19503 2374
tri 19503 2367 19510 2374 nw
tri 20304 2367 20311 2374 ne
rect 20311 2367 20354 2374
tri 20354 2367 20361 2374 sw
tri 21233 2367 21240 2374 se
rect 21240 2367 21283 2374
tri 21283 2367 21290 2374 nw
rect 18547 916 18553 968
rect 18605 916 18617 968
rect 18669 916 18675 968
tri 18761 1875 18797 1911 se
rect 18797 1889 18849 2202
tri 18849 2180 18871 2202 nw
rect 18797 1875 18835 1889
tri 18835 1875 18849 1889 nw
rect 18878 2100 18884 2152
rect 18936 2100 18948 2152
rect 19000 2100 19006 2152
rect 18290 454 18296 506
rect 18348 454 18360 506
rect 18412 454 18418 506
rect 9655 -197 9690 -196
rect 8337 -199 8395 -197
tri 8395 -199 8397 -197 sw
rect 8463 -199 9584 -197
tri 9584 -199 9586 -197 nw
tri 9629 -199 9631 -197 se
rect 9631 -199 9690 -197
rect 8337 -200 8397 -199
tri 8397 -200 8398 -199 sw
rect 8463 -200 9583 -199
tri 9583 -200 9584 -199 nw
tri 9628 -200 9629 -199 se
rect 9629 -200 9690 -199
rect 8337 -201 8398 -200
tri 8398 -201 8399 -200 sw
rect 8463 -201 9582 -200
tri 9582 -201 9583 -200 nw
tri 9627 -201 9628 -200 se
rect 9628 -201 9690 -200
tri 9690 -201 9695 -196 nw
rect 8337 -226 8399 -201
tri 8399 -226 8424 -201 sw
rect 8463 -209 9574 -201
tri 9574 -209 9582 -201 nw
tri 9619 -209 9627 -201 se
rect 9627 -209 9665 -201
tri 9602 -226 9619 -209 se
rect 9619 -226 9665 -209
tri 9665 -226 9690 -201 nw
rect 17313 -226 17348 446
rect 8337 -237 8424 -226
tri 8424 -237 8435 -226 sw
tri 9591 -237 9602 -226 se
rect 9602 -237 9654 -226
tri 9654 -237 9665 -226 nw
tri 9704 -237 9715 -226 se
rect 9715 -237 17348 -226
rect 8337 -239 9652 -237
tri 9652 -239 9654 -237 nw
tri 9702 -239 9704 -237 se
rect 9704 -239 17348 -237
rect 8337 -254 9637 -239
tri 9637 -254 9652 -239 nw
tri 9687 -254 9702 -239 se
rect 9702 -254 17348 -239
tri 8337 -261 8344 -254 ne
rect 8344 -261 9622 -254
tri 8267 -269 8275 -261 sw
tri 8344 -269 8352 -261 ne
rect 8352 -269 9622 -261
tri 9622 -269 9637 -254 nw
tri 9672 -269 9687 -254 se
rect 9687 -261 17348 -254
rect 17386 278 17392 330
rect 17444 278 17456 330
rect 17508 278 17514 330
rect 9687 -269 9715 -261
rect 8211 -289 8275 -269
tri 8275 -289 8295 -269 sw
tri 9652 -289 9672 -269 se
rect 9672 -289 9715 -269
tri 9715 -289 9743 -261 nw
rect 8211 -298 8295 -289
tri 8295 -298 8304 -289 sw
tri 9643 -298 9652 -289 se
rect 9652 -290 9714 -289
tri 9714 -290 9715 -289 nw
rect 17386 -290 17421 278
rect 9652 -298 9706 -290
tri 9706 -298 9714 -290 nw
tri 9760 -298 9768 -290 se
rect 9768 -298 17421 -290
rect 8211 -299 9705 -298
tri 9705 -299 9706 -298 nw
tri 9759 -299 9760 -298 se
rect 9760 -299 17421 -298
rect 8211 -303 9701 -299
tri 9701 -303 9705 -299 nw
tri 9755 -303 9759 -299 se
rect 9759 -303 17421 -299
tri 8211 -334 8242 -303 ne
rect 8242 -334 9670 -303
tri 9670 -334 9701 -303 nw
tri 9724 -334 9755 -303 se
rect 9755 -325 17421 -303
rect 17477 173 17529 179
rect 17477 109 17529 121
rect 17477 41 17529 57
rect 9755 -334 9768 -325
tri 9705 -353 9724 -334 se
rect 9724 -353 9768 -334
tri 9768 -353 9796 -325 nw
tri 9696 -362 9705 -353 se
rect 9705 -362 9759 -353
tri 9759 -362 9768 -353 nw
rect 17477 -355 17512 41
tri 17512 24 17529 41 nw
rect 18547 -50 18583 916
tri 18742 790 18761 809 se
rect 18761 790 18813 1875
tri 18813 1853 18835 1875 nw
rect 18878 1157 18924 2100
rect 18846 1105 18852 1157
rect 18904 1105 18916 1157
rect 18968 1105 18974 1157
rect 18878 923 18924 1105
tri 18924 923 18937 936 sw
rect 18878 916 18937 923
tri 18878 911 18883 916 ne
rect 18883 911 18937 916
tri 18937 911 18949 923 sw
tri 18883 891 18903 911 ne
tri 18664 738 18716 790 se
rect 18716 738 18741 790
rect 18793 738 18805 790
rect 18857 738 18863 790
tri 18662 736 18664 738 se
rect 18664 736 18733 738
tri 18733 736 18735 738 nw
tri 18645 719 18662 736 se
rect 18662 719 18716 736
tri 18716 719 18733 736 nw
tri 18886 719 18903 736 se
rect 18903 719 18949 911
rect 18455 -102 18461 -50
rect 18513 -102 18525 -50
rect 18577 -102 18583 -50
tri 18625 699 18645 719 se
rect 18645 699 18696 719
tri 18696 699 18716 719 nw
tri 18866 699 18886 719 se
rect 18886 716 18949 719
rect 18886 699 18903 716
rect 18625 -149 18677 699
tri 18677 680 18696 699 nw
tri 18847 680 18866 699 se
rect 18866 680 18903 699
tri 18837 670 18847 680 se
rect 18847 670 18903 680
tri 18903 670 18949 716 nw
tri 18809 642 18837 670 se
rect 18837 642 18875 670
tri 18875 642 18903 670 nw
tri 19325 642 19346 663 se
rect 19346 642 19376 2367
tri 19376 2361 19382 2367 nw
tri 19441 2361 19447 2367 se
rect 19447 2361 19492 2367
tri 19436 2356 19441 2361 se
rect 19441 2356 19492 2361
tri 19492 2356 19503 2367 nw
tri 20311 2356 20322 2367 ne
rect 20322 2364 20361 2367
tri 20361 2364 20364 2367 sw
tri 21230 2364 21233 2367 se
rect 21233 2364 21253 2367
rect 20322 2356 21253 2364
tri 19422 2342 19436 2356 se
rect 19436 2342 19478 2356
tri 19478 2342 19492 2356 nw
tri 20322 2342 20336 2356 ne
rect 20336 2342 21253 2356
rect 18809 629 18862 642
tri 18862 629 18875 642 nw
tri 19312 629 19325 642 se
rect 19325 629 19376 642
rect 18809 -62 18855 629
tri 18855 622 18862 629 nw
rect 19248 577 19254 629
rect 19306 577 19318 629
rect 19370 577 19376 629
tri 19406 2326 19422 2342 se
rect 19422 2326 19436 2342
tri 19396 526 19406 536 se
rect 19406 526 19436 2326
tri 19436 2300 19478 2342 nw
rect 19964 2290 19970 2342
rect 20022 2290 20034 2342
rect 20086 2290 20092 2342
tri 20336 2337 20341 2342 ne
rect 20341 2337 21253 2342
tri 21253 2337 21283 2367 nw
tri 20341 2334 20344 2337 ne
rect 20344 2334 21250 2337
tri 21250 2334 21253 2337 nw
rect 19634 2100 19640 2152
rect 19692 2100 19704 2152
rect 19756 2100 19762 2152
rect 19647 942 19693 2100
rect 20040 2058 20092 2290
tri 21231 2245 21283 2297 se
rect 21283 2245 21365 2297
rect 21417 2245 21429 2297
rect 21481 2245 21487 2297
tri 21224 2238 21231 2245 se
rect 21231 2238 21273 2245
rect 20213 2232 20265 2238
tri 21207 2221 21224 2238 se
rect 21224 2221 21273 2238
tri 21273 2221 21297 2245 nw
tri 21195 2209 21207 2221 se
rect 21207 2209 21261 2221
tri 21261 2209 21273 2221 nw
tri 21193 2207 21195 2209 se
rect 21195 2207 21259 2209
tri 21259 2207 21261 2209 nw
tri 21190 2204 21193 2207 se
rect 21193 2204 21256 2207
tri 21256 2204 21259 2207 nw
tri 21170 2184 21190 2204 se
rect 21190 2184 21207 2204
rect 20265 2180 21207 2184
rect 20213 2168 21207 2180
rect 20265 2155 21207 2168
tri 21207 2155 21256 2204 nw
rect 20265 2143 21195 2155
tri 21195 2143 21207 2155 nw
rect 20265 2138 21190 2143
tri 21190 2138 21195 2143 nw
rect 20213 2110 20265 2116
tri 20092 2058 20098 2064 sw
rect 20501 2058 20507 2110
rect 20559 2058 20571 2110
rect 20623 2058 20931 2110
rect 20969 2058 20975 2110
rect 21027 2058 21039 2110
rect 21091 2058 21097 2110
rect 20040 2047 20098 2058
tri 20098 2047 20109 2058 sw
rect 20040 2042 20109 2047
tri 20040 1973 20109 2042 ne
tri 20109 1973 20183 2047 sw
rect 20892 2013 20931 2058
rect 20892 1974 20970 2013
tri 20109 1899 20183 1973 ne
tri 20183 1899 20257 1973 sw
tri 20183 1877 20205 1899 ne
tri 19693 942 19701 950 sw
rect 19647 936 19701 942
tri 19701 936 19707 942 sw
rect 19647 930 19707 936
tri 19647 923 19654 930 ne
rect 19654 923 19707 930
tri 19707 923 19720 936 sw
tri 19654 895 19682 923 ne
rect 19682 895 19720 923
tri 19720 895 19748 923 sw
tri 19682 892 19685 895 ne
rect 19685 892 20014 895
tri 20014 892 20017 895 sw
tri 19685 890 19687 892 ne
rect 19687 890 20017 892
tri 20017 890 20019 892 sw
tri 19687 884 19693 890 ne
rect 19693 884 20019 890
tri 19693 877 19700 884 ne
rect 19700 877 20019 884
tri 20019 877 20032 890 sw
tri 19700 860 19717 877 ne
rect 19717 860 20032 877
tri 19983 826 20017 860 ne
rect 20017 826 20032 860
tri 20032 826 20083 877 sw
tri 20017 825 20018 826 ne
rect 20018 825 20084 826
tri 20018 813 20030 825 ne
rect 20030 813 20084 825
tri 20030 805 20038 813 ne
tri 20027 642 20038 653 se
rect 20038 642 20084 813
tri 20014 629 20027 642 se
rect 20027 629 20084 642
rect 19248 474 19254 526
rect 19306 474 19318 526
rect 19370 510 19436 526
rect 19370 488 19414 510
tri 19414 488 19436 510 nw
tri 20007 622 20014 629 se
rect 20014 628 20084 629
rect 20014 622 20078 628
tri 20078 622 20084 628 nw
rect 20007 612 20068 622
tri 20068 612 20078 622 nw
rect 19370 474 19400 488
tri 19400 474 19414 488 nw
rect 20007 175 20053 612
tri 20053 597 20068 612 nw
rect 20205 259 20257 1899
rect 20751 1818 20868 1820
rect 20740 1791 20868 1818
rect 20740 1739 20746 1791
rect 20798 1739 20810 1791
rect 20862 1739 20868 1791
rect 20740 1712 20868 1739
rect 20751 488 20868 1712
rect 20931 1629 20970 1974
rect 21034 1705 21073 2058
rect 21034 1666 21691 1705
rect 20931 1590 21622 1629
tri 21577 890 21583 896 se
rect 21583 890 21622 1590
tri 21570 883 21577 890 se
rect 21577 883 21622 890
rect 21570 877 21622 883
rect 21570 813 21622 825
rect 21570 755 21622 761
rect 21652 890 21691 1666
rect 21768 1666 21826 2965
tri 22092 2945 22112 2965 ne
rect 22112 2945 22166 2965
tri 22166 2945 22186 2965 sw
tri 22112 2929 22128 2945 ne
rect 21768 1614 21771 1666
rect 21823 1614 21826 1666
rect 21768 1594 21826 1614
rect 21768 1542 21771 1594
rect 21823 1542 21826 1594
rect 21768 1536 21826 1542
rect 22128 1678 22186 2945
rect 22983 2742 22989 2794
rect 23041 2742 23053 2794
rect 23105 2742 23111 2794
tri 23038 2736 23044 2742 ne
rect 23044 2736 23111 2742
tri 23044 2732 23048 2736 ne
rect 23048 2732 23111 2736
rect 22731 2680 22737 2732
rect 22789 2680 22801 2732
rect 22853 2680 22859 2732
tri 23048 2725 23055 2732 ne
rect 23055 2725 23111 2732
tri 23055 2708 23072 2725 ne
tri 22786 2673 22793 2680 ne
rect 22793 2673 22859 2680
tri 22793 2646 22820 2673 ne
rect 22820 2459 22859 2673
rect 23072 2459 23111 2725
rect 22820 2453 22872 2459
rect 22407 2367 22413 2419
rect 22465 2367 22477 2419
rect 22529 2367 22535 2419
rect 23072 2407 23078 2459
rect 23130 2407 23142 2459
rect 23194 2407 23200 2459
rect 22820 2389 22872 2401
rect 22820 2331 22872 2337
tri 22929 2331 22953 2355 se
rect 22953 2331 23217 2355
tri 23217 2331 23241 2355 sw
tri 22903 2305 22929 2331 se
rect 22929 2305 23241 2331
rect 22903 2303 23241 2305
rect 22903 2296 22968 2303
tri 22968 2296 22975 2303 nw
tri 23195 2296 23202 2303 ne
rect 23202 2296 23241 2303
tri 23241 2296 23276 2331 sw
rect 22903 2273 22955 2296
tri 22955 2283 22968 2296 nw
tri 23202 2283 23215 2296 ne
rect 23215 2283 23276 2296
tri 23215 2281 23217 2283 ne
rect 23217 2281 23276 2283
tri 23217 2274 23224 2281 ne
rect 22903 2207 22955 2221
rect 22903 2149 22955 2155
rect 23084 2261 23136 2267
rect 23084 2195 23136 2209
tri 23016 2010 23084 2078 se
rect 23084 2056 23136 2143
rect 23084 2010 23090 2056
tri 23090 2010 23136 2056 nw
tri 22942 1811 23016 1885 se
rect 23016 1867 23072 2010
tri 23072 1992 23090 2010 nw
tri 23016 1811 23072 1867 nw
tri 22868 1737 22942 1811 se
tri 22942 1737 23016 1811 nw
tri 22853 1722 22868 1737 se
rect 22868 1722 22927 1737
tri 22927 1722 22942 1737 nw
tri 22186 1678 22189 1681 sw
rect 22853 1678 22905 1722
tri 22905 1700 22927 1722 nw
rect 22128 1661 22189 1678
tri 22189 1661 22206 1678 sw
rect 22128 1655 22206 1661
rect 22128 1603 22154 1655
tri 22821 1626 22853 1658 se
tri 22807 1612 22821 1626 se
rect 22821 1612 22905 1626
rect 22128 1583 22206 1603
tri 22793 1598 22807 1612 se
rect 22807 1598 22853 1612
rect 22128 1531 22154 1583
tri 22511 1560 22549 1598 se
rect 22549 1560 22853 1598
tri 22497 1546 22511 1560 se
rect 22511 1546 22905 1560
rect 23224 1585 23276 2281
tri 23276 1585 23310 1619 sw
rect 22128 1525 22206 1531
rect 22469 1536 22549 1546
tri 22549 1536 22559 1546 nw
rect 22469 1533 22546 1536
tri 22546 1533 22549 1536 nw
rect 23224 1533 23230 1585
rect 23282 1533 23294 1585
rect 23346 1533 23352 1585
tri 22468 1517 22469 1518 se
rect 22469 1517 22530 1533
tri 22530 1517 22546 1533 nw
rect 23224 1525 23284 1533
tri 23284 1525 23292 1533 nw
rect 23224 1517 23276 1525
tri 23276 1517 23284 1525 nw
tri 22430 1479 22468 1517 se
rect 22468 1479 22492 1517
tri 22492 1479 22530 1517 nw
rect 23224 1515 23274 1517
tri 23274 1515 23276 1517 nw
tri 23188 1479 23224 1515 se
rect 23224 1479 23238 1515
tri 23238 1479 23274 1515 nw
tri 22427 1476 22430 1479 se
rect 22430 1476 22489 1479
tri 22489 1476 22492 1479 nw
tri 23185 1476 23188 1479 se
rect 23188 1476 23232 1479
tri 22425 1474 22427 1476 se
rect 22427 1474 22487 1476
tri 22487 1474 22489 1476 nw
tri 22424 1473 22425 1474 se
rect 22425 1473 22486 1474
tri 22486 1473 22487 1474 nw
tri 22421 1470 22424 1473 se
rect 22424 1470 22483 1473
tri 22483 1470 22486 1473 nw
rect 22950 1470 23002 1476
tri 23182 1473 23185 1476 se
rect 23185 1473 23232 1476
tri 23232 1473 23238 1479 nw
rect 23327 1473 23379 1479
tri 22369 1418 22421 1470 se
rect 22421 1418 22431 1470
tri 22431 1418 22483 1470 nw
tri 23174 1465 23182 1473 se
rect 23182 1465 23224 1473
tri 23224 1465 23232 1473 nw
tri 23130 1421 23174 1465 se
rect 23174 1421 23180 1465
tri 23180 1421 23224 1465 nw
tri 22363 1412 22369 1418 se
rect 22369 1412 22425 1418
tri 22425 1412 22431 1418 nw
tri 22360 1409 22363 1412 se
rect 22363 1409 22422 1412
tri 22422 1409 22425 1412 nw
tri 22357 1406 22360 1409 se
rect 22360 1406 22419 1409
tri 22419 1406 22422 1409 nw
rect 22950 1406 23002 1418
tri 23124 1415 23130 1421 se
rect 23130 1415 23174 1421
tri 23174 1415 23180 1421 nw
tri 23118 1409 23124 1415 se
rect 23124 1409 23168 1415
tri 23168 1409 23174 1415 nw
rect 23327 1409 23379 1421
tri 22353 1402 22357 1406 se
rect 22357 1402 22415 1406
tri 22415 1402 22419 1406 nw
tri 22279 1123 22353 1197 se
rect 22353 1167 22397 1402
tri 22397 1384 22415 1402 nw
tri 23074 1365 23118 1409 se
rect 23118 1365 23124 1409
tri 23124 1365 23168 1409 nw
tri 23066 1357 23074 1365 se
rect 23074 1357 23116 1365
tri 23116 1357 23124 1365 nw
tri 22889 1287 22950 1348 se
rect 22950 1339 23002 1354
tri 23060 1351 23066 1357 se
rect 23066 1351 23110 1357
tri 23110 1351 23116 1357 nw
rect 22950 1315 22978 1339
tri 22978 1315 23002 1339 nw
tri 23024 1315 23060 1351 se
rect 23060 1315 23074 1351
tri 23074 1315 23110 1351 nw
rect 22950 1311 22974 1315
tri 22974 1311 22978 1315 nw
tri 23020 1311 23024 1315 se
tri 22950 1287 22974 1311 nw
tri 22996 1287 23020 1311 se
rect 23020 1287 23024 1311
tri 22879 1277 22889 1287 se
rect 22889 1277 22940 1287
tri 22940 1277 22950 1287 nw
tri 22986 1277 22996 1287 se
rect 22996 1277 23024 1287
tri 22353 1123 22397 1167 nw
tri 22590 1227 22640 1277 se
rect 22640 1265 22928 1277
tri 22928 1265 22940 1277 nw
tri 22974 1265 22986 1277 se
rect 22986 1265 23024 1277
tri 23024 1265 23074 1315 nw
rect 23327 1286 23379 1357
rect 23327 1284 23377 1286
tri 23377 1284 23379 1286 nw
tri 23308 1265 23327 1284 se
rect 22640 1261 22924 1265
tri 22924 1261 22928 1265 nw
tri 22970 1261 22974 1265 se
rect 22640 1241 22904 1261
tri 22904 1241 22924 1261 nw
tri 22950 1241 22970 1261 se
rect 22970 1241 22974 1261
rect 22640 1227 22648 1241
tri 22648 1227 22662 1241 nw
tri 22936 1227 22950 1241 se
rect 22950 1227 22974 1241
tri 22252 1096 22279 1123 se
rect 22279 1096 22287 1123
rect 21720 1077 21862 1096
rect 21720 1025 21726 1077
rect 21778 1025 21804 1077
rect 21856 1025 21862 1077
tri 22213 1057 22252 1096 se
rect 22252 1057 22287 1096
tri 22287 1057 22353 1123 nw
tri 22205 1049 22213 1057 se
rect 22213 1049 22279 1057
tri 22279 1049 22287 1057 nw
tri 22582 1049 22590 1057 se
rect 22590 1049 22626 1227
tri 22626 1205 22648 1227 nw
tri 22924 1215 22936 1227 se
rect 22936 1215 22974 1227
tri 22974 1215 23024 1265 nw
tri 23277 1234 23308 1265 se
rect 23308 1234 23327 1265
tri 23327 1234 23377 1284 nw
tri 23258 1215 23277 1234 se
tri 22914 1205 22924 1215 se
rect 22924 1205 22956 1215
tri 22906 1197 22914 1205 se
rect 22914 1197 22956 1205
tri 22956 1197 22974 1215 nw
tri 23240 1197 23258 1215 se
rect 23258 1197 23277 1215
rect 21720 937 21862 1025
tri 22168 1012 22205 1049 se
rect 22205 1012 22242 1049
tri 22242 1012 22279 1049 nw
tri 22545 1012 22582 1049 se
rect 22582 1043 22626 1049
rect 22582 1012 22595 1043
tri 22595 1012 22626 1043 nw
tri 22660 1165 22692 1197 se
rect 22692 1165 22924 1197
tri 22924 1165 22956 1197 nw
tri 23227 1184 23240 1197 se
rect 23240 1184 23277 1197
tri 23277 1184 23327 1234 nw
tri 23208 1165 23227 1184 se
rect 22660 1161 22920 1165
tri 22920 1161 22924 1165 nw
tri 23204 1161 23208 1165 se
rect 23208 1161 23227 1165
tri 22646 1012 22660 1026 se
rect 22660 1012 22696 1161
tri 22696 1151 22706 1161 nw
tri 23194 1151 23204 1161 se
rect 23204 1151 23227 1161
tri 23177 1134 23194 1151 se
rect 23194 1134 23227 1151
tri 23227 1134 23277 1184 nw
tri 23166 1123 23177 1134 se
rect 23177 1123 23216 1134
tri 23216 1123 23227 1134 nw
tri 22728 1073 22778 1123 se
rect 22778 1087 23180 1123
tri 23180 1087 23216 1123 nw
tri 22778 1073 22792 1087 nw
tri 22162 1006 22168 1012 se
rect 22168 1006 22236 1012
tri 22236 1006 22242 1012 nw
rect 22543 1006 22595 1012
tri 22131 975 22162 1006 se
rect 22162 975 22205 1006
tri 22205 975 22236 1006 nw
tri 22110 954 22131 975 se
rect 22131 954 22184 975
tri 22184 954 22205 975 nw
tri 22098 942 22110 954 se
rect 22110 942 22172 954
tri 22172 942 22184 954 nw
rect 22543 942 22595 954
tri 21720 915 21742 937 ne
tri 21691 890 21697 896 sw
rect 21652 883 21697 890
tri 21697 883 21704 890 sw
rect 21652 877 21704 883
rect 21652 813 21704 825
rect 21652 755 21704 761
rect 20740 308 20746 488
rect 20862 308 20868 488
tri 21718 653 21742 677 se
rect 21742 653 21862 937
rect 21718 612 21862 653
rect 21770 560 21810 612
rect 21718 523 21862 560
rect 21770 471 21810 523
rect 21718 465 21862 471
tri 22087 931 22098 942 se
rect 22098 931 22161 942
tri 22161 931 22172 942 nw
rect 22087 479 22139 931
tri 22139 909 22161 931 nw
rect 22543 884 22595 890
tri 22626 992 22646 1012 se
rect 22646 992 22676 1012
tri 22676 992 22696 1012 nw
tri 22724 1069 22728 1073 se
rect 22728 1069 22774 1073
tri 22774 1069 22778 1073 nw
tri 22623 869 22626 872 se
rect 22626 869 22663 992
tri 22663 979 22676 992 nw
tri 22711 979 22724 992 se
rect 22724 979 22760 1069
tri 22760 1055 22774 1069 nw
tri 22611 857 22623 869 se
rect 22623 859 22663 869
rect 22623 857 22661 859
tri 22661 857 22663 859 nw
tri 22693 961 22711 979 se
rect 22711 978 22760 979
rect 22711 961 22745 978
tri 22745 963 22760 978 nw
rect 22693 921 22745 961
rect 22693 857 22745 869
tri 22576 822 22611 857 se
rect 22611 822 22626 857
tri 22626 822 22661 857 nw
tri 22559 805 22576 822 se
rect 22576 805 22609 822
tri 22609 805 22626 822 nw
tri 22553 799 22559 805 se
rect 22559 799 22603 805
tri 22603 799 22609 805 nw
rect 22693 799 22745 805
tri 22526 772 22553 799 se
rect 22553 772 22576 799
tri 22576 772 22603 799 nw
tri 22519 765 22526 772 se
rect 22526 765 22569 772
tri 22569 765 22576 772 nw
rect 22474 713 22517 765
tri 22517 713 22569 765 nw
rect 22087 415 22139 427
rect 22087 357 22139 363
rect 20751 300 20868 308
rect 20129 207 20135 259
rect 20187 207 20199 259
rect 20251 207 20257 259
rect 19967 123 19973 175
rect 20025 123 20037 175
rect 20089 123 20095 175
rect 18751 -114 18757 -62
rect 18809 -114 18821 -62
rect 18873 -114 18879 -62
rect 18580 -201 18586 -149
rect 18638 -201 18650 -149
rect 18702 -201 18708 -149
tri 9828 -362 9835 -355 se
rect 9835 -362 17512 -355
rect 4816 -414 4822 -362
rect 4874 -414 4886 -362
rect 4938 -414 4944 -362
rect 5077 -398 9723 -362
tri 9723 -398 9759 -362 nw
tri 9792 -398 9828 -362 se
rect 9828 -390 17512 -362
rect 9828 -398 9835 -390
tri 9776 -414 9792 -398 se
rect 9792 -414 9835 -398
tri 9772 -418 9776 -414 se
rect 9776 -418 9835 -414
tri 9835 -418 9863 -390 nw
tri 9763 -427 9772 -418 se
rect 9772 -427 9826 -418
tri 9826 -427 9835 -418 nw
rect 5028 -463 9790 -427
tri 9790 -463 9826 -427 nw
<< via2 >>
rect 8589 2578 8645 2634
rect 8669 2578 8725 2634
rect 8463 2485 8519 2541
rect 8337 2402 8393 2458
rect 8211 2322 8267 2378
rect 8463 2405 8519 2461
rect 8337 2322 8393 2378
rect 8211 2242 8267 2298
rect 17863 2719 17919 2775
rect 17944 2719 18000 2775
rect 18025 2719 18081 2775
rect 18105 2719 18161 2775
rect 18185 2719 18241 2775
rect 8589 4 8645 60
rect 8211 -111 8267 -55
rect 8211 -191 8267 -135
rect 8337 -110 8393 -54
rect 8337 -190 8393 -134
rect 8463 -108 8519 -52
rect 8463 -188 8519 -132
rect 8589 -76 8645 -20
rect 20287 2779 20343 2835
rect 20368 2779 20424 2835
rect 20287 2699 20343 2755
rect 20368 2699 20424 2755
rect 20449 2699 20665 2835
<< metal3 >>
rect 20282 2835 20670 2840
rect 17858 2775 18246 2780
rect 17858 2719 17863 2775
rect 17919 2719 17944 2775
rect 18000 2719 18025 2775
rect 18081 2719 18105 2775
rect 18161 2719 18185 2775
rect 18241 2719 18246 2775
rect 8584 2634 8730 2639
rect 8584 2578 8589 2634
rect 8645 2578 8669 2634
rect 8725 2578 8730 2634
rect 8584 2573 8730 2578
rect 8458 2541 8524 2551
rect 8458 2485 8463 2541
rect 8519 2485 8524 2541
rect 8332 2458 8398 2467
rect 8332 2402 8337 2458
rect 8393 2402 8398 2458
rect 8206 2378 8272 2383
rect 8206 2322 8211 2378
rect 8267 2322 8272 2378
rect 8206 2298 8272 2322
rect 8206 2242 8211 2298
rect 8267 2242 8272 2298
rect 8206 -55 8272 2242
rect 8206 -111 8211 -55
rect 8267 -111 8272 -55
rect 8206 -135 8272 -111
rect 8206 -191 8211 -135
rect 8267 -191 8272 -135
rect 8206 -196 8272 -191
rect 8332 2378 8398 2402
rect 8332 2322 8337 2378
rect 8393 2322 8398 2378
rect 8332 -54 8398 2322
rect 8332 -110 8337 -54
rect 8393 -110 8398 -54
rect 8332 -134 8398 -110
rect 8332 -190 8337 -134
rect 8393 -190 8398 -134
rect 8332 -195 8398 -190
rect 8458 2461 8524 2485
rect 8458 2405 8463 2461
rect 8519 2405 8524 2461
rect 8458 -52 8524 2405
rect 8458 -108 8463 -52
rect 8519 -108 8524 -52
rect 8584 60 8650 2573
rect 17858 1302 18246 2719
rect 20282 2779 20287 2835
rect 20343 2779 20368 2835
rect 20424 2779 20449 2835
rect 20282 2755 20449 2779
rect 20282 2699 20287 2755
rect 20343 2699 20368 2755
rect 20424 2699 20449 2755
rect 20665 2699 20670 2835
rect 8584 4 8589 60
rect 8645 4 8650 60
rect 8584 -20 8650 4
rect 8584 -76 8589 -20
rect 8645 -76 8650 -20
rect 8584 -81 8650 -76
rect 20282 525 20670 2699
rect 20282 461 20284 525
rect 20348 461 20364 525
rect 20428 461 20444 525
rect 20508 461 20524 525
rect 20588 461 20604 525
rect 20668 461 20670 525
rect 20282 439 20670 461
rect 20282 375 20284 439
rect 20348 375 20364 439
rect 20428 375 20444 439
rect 20508 375 20524 439
rect 20588 375 20604 439
rect 20668 375 20670 439
rect 20282 353 20670 375
rect 20282 289 20284 353
rect 20348 289 20364 353
rect 20428 289 20444 353
rect 20508 289 20524 353
rect 20588 289 20604 353
rect 20668 289 20670 353
rect 20282 267 20670 289
rect 20282 203 20284 267
rect 20348 203 20364 267
rect 20428 203 20444 267
rect 20508 203 20524 267
rect 20588 203 20604 267
rect 20668 203 20670 267
rect 20282 181 20670 203
rect 20282 117 20284 181
rect 20348 117 20364 181
rect 20428 117 20444 181
rect 20508 117 20524 181
rect 20588 117 20604 181
rect 20668 117 20670 181
rect 20282 95 20670 117
rect 20282 31 20284 95
rect 20348 31 20364 95
rect 20428 31 20444 95
rect 20508 31 20524 95
rect 20588 31 20604 95
rect 20668 31 20670 95
rect 20282 9 20670 31
rect 20282 -55 20284 9
rect 20348 -55 20364 9
rect 20428 -55 20444 9
rect 20508 -55 20524 9
rect 20588 -55 20604 9
rect 20668 -55 20670 9
rect 20282 -78 20670 -55
rect 8458 -132 8524 -108
rect 8458 -188 8463 -132
rect 8519 -188 8524 -132
rect 8458 -193 8524 -188
rect 20282 -142 20284 -78
rect 20348 -142 20364 -78
rect 20428 -142 20444 -78
rect 20508 -142 20524 -78
rect 20588 -142 20604 -78
rect 20668 -142 20670 -78
rect 20282 -165 20670 -142
rect 20282 -229 20284 -165
rect 20348 -229 20364 -165
rect 20428 -229 20444 -165
rect 20508 -229 20524 -165
rect 20588 -229 20604 -165
rect 20668 -229 20670 -165
rect 20282 -252 20670 -229
rect 20282 -316 20284 -252
rect 20348 -316 20364 -252
rect 20428 -316 20444 -252
rect 20508 -316 20524 -252
rect 20588 -316 20604 -252
rect 20668 -316 20670 -252
rect 20282 -339 20670 -316
rect 20282 -403 20284 -339
rect 20348 -403 20364 -339
rect 20428 -403 20444 -339
rect 20508 -403 20524 -339
rect 20588 -403 20604 -339
rect 20668 -403 20670 -339
rect 20282 -409 20670 -403
<< via3 >>
rect 20284 461 20348 525
rect 20364 461 20428 525
rect 20444 461 20508 525
rect 20524 461 20588 525
rect 20604 461 20668 525
rect 20284 375 20348 439
rect 20364 375 20428 439
rect 20444 375 20508 439
rect 20524 375 20588 439
rect 20604 375 20668 439
rect 20284 289 20348 353
rect 20364 289 20428 353
rect 20444 289 20508 353
rect 20524 289 20588 353
rect 20604 289 20668 353
rect 20284 203 20348 267
rect 20364 203 20428 267
rect 20444 203 20508 267
rect 20524 203 20588 267
rect 20604 203 20668 267
rect 20284 117 20348 181
rect 20364 117 20428 181
rect 20444 117 20508 181
rect 20524 117 20588 181
rect 20604 117 20668 181
rect 20284 31 20348 95
rect 20364 31 20428 95
rect 20444 31 20508 95
rect 20524 31 20588 95
rect 20604 31 20668 95
rect 20284 -55 20348 9
rect 20364 -55 20428 9
rect 20444 -55 20508 9
rect 20524 -55 20588 9
rect 20604 -55 20668 9
rect 20284 -142 20348 -78
rect 20364 -142 20428 -78
rect 20444 -142 20508 -78
rect 20524 -142 20588 -78
rect 20604 -142 20668 -78
rect 20284 -229 20348 -165
rect 20364 -229 20428 -165
rect 20444 -229 20508 -165
rect 20524 -229 20588 -165
rect 20604 -229 20668 -165
rect 20284 -316 20348 -252
rect 20364 -316 20428 -252
rect 20444 -316 20508 -252
rect 20524 -316 20588 -252
rect 20604 -316 20668 -252
rect 20284 -403 20348 -339
rect 20364 -403 20428 -339
rect 20444 -403 20508 -339
rect 20524 -403 20588 -339
rect 20604 -403 20668 -339
<< metal4 >>
rect 20281 525 20671 526
rect 20281 461 20284 525
rect 20348 461 20364 525
rect 20428 461 20444 525
rect 20508 461 20524 525
rect 20588 461 20604 525
rect 20668 461 20671 525
rect 20281 439 20671 461
rect 20281 375 20284 439
rect 20348 375 20364 439
rect 20428 375 20444 439
rect 20508 375 20524 439
rect 20588 375 20604 439
rect 20668 375 20671 439
rect 20281 353 20671 375
rect 20281 289 20284 353
rect 20348 289 20364 353
rect 20428 289 20444 353
rect 20508 289 20524 353
rect 20588 289 20604 353
rect 20668 289 20671 353
rect 20281 267 20671 289
rect 20281 203 20284 267
rect 20348 203 20364 267
rect 20428 203 20444 267
rect 20508 203 20524 267
rect 20588 203 20604 267
rect 20668 203 20671 267
rect 20281 181 20671 203
rect 20281 117 20284 181
rect 20348 117 20364 181
rect 20428 117 20444 181
rect 20508 117 20524 181
rect 20588 117 20604 181
rect 20668 117 20671 181
rect 20281 95 20671 117
rect 20281 31 20284 95
rect 20348 31 20364 95
rect 20428 31 20444 95
rect 20508 31 20524 95
rect 20588 31 20604 95
rect 20668 31 20671 95
rect 20281 9 20671 31
rect 20281 -55 20284 9
rect 20348 -55 20364 9
rect 20428 -55 20444 9
rect 20508 -55 20524 9
rect 20588 -55 20604 9
rect 20668 -55 20671 9
rect 20281 -78 20671 -55
rect 20281 -142 20284 -78
rect 20348 -142 20364 -78
rect 20428 -142 20444 -78
rect 20508 -142 20524 -78
rect 20588 -142 20604 -78
rect 20668 -142 20671 -78
rect 20281 -165 20671 -142
rect 20281 -229 20284 -165
rect 20348 -229 20364 -165
rect 20428 -229 20444 -165
rect 20508 -229 20524 -165
rect 20588 -229 20604 -165
rect 20668 -229 20671 -165
rect 20281 -252 20671 -229
rect 20281 -316 20284 -252
rect 20348 -316 20364 -252
rect 20428 -316 20444 -252
rect 20508 -316 20524 -252
rect 20588 -316 20604 -252
rect 20668 -316 20671 -252
rect 20281 -339 20671 -316
rect 20281 -403 20284 -339
rect 20348 -403 20364 -339
rect 20428 -403 20444 -339
rect 20508 -403 20524 -339
rect 20588 -403 20604 -339
rect 20668 -403 20671 -339
rect 20281 -404 20671 -403
use sky130_fd_io__gpio_ovtv2_amux_drvr_lshv2hv_1  sky130_fd_io__gpio_ovtv2_amux_drvr_lshv2hv_1_0
timestamp 1640697850
transform 1 0 6 0 1 0
box -43 1398 15108 3122
use sky130_fd_io__gpio_ovtv2_amux_drvr_lshv2hv  sky130_fd_io__gpio_ovtv2_amux_drvr_lshv2hv_0
timestamp 1640697850
transform 1 0 9 0 1 -14
box -6 52 14977 2964
use sky130_fd_io__gpio_ovtv2_amux_drvr_ls_1  sky130_fd_io__gpio_ovtv2_amux_drvr_ls_1_0
timestamp 1640697850
transform 1 0 1252 0 1 49
box 0 10 6326 2677
use sky130_fd_io__gpio_ovtv2_amux_drvr_ls  sky130_fd_io__gpio_ovtv2_amux_drvr_ls_0
timestamp 1640697850
transform 1 0 1252 0 1 49
box 0 -208 4912 2661
use sky130_fd_pr__nfet_01v8__example_55959141808511  sky130_fd_pr__nfet_01v8__example_55959141808511_0
timestamp 1640697850
transform 0 1 3632 -1 0 906
box -28 0 324 29
use sky130_fd_pr__nfet_01v8__example_55959141808511  sky130_fd_pr__nfet_01v8__example_55959141808511_1
timestamp 1640697850
transform 0 1 3418 -1 0 906
box -28 0 324 29
use sky130_fd_pr__nfet_01v8__example_55959141808511  sky130_fd_pr__nfet_01v8__example_55959141808511_2
timestamp 1640697850
transform 0 1 3880 1 0 144
box -28 0 324 29
use sky130_fd_pr__nfet_01v8__example_55959141808511  sky130_fd_pr__nfet_01v8__example_55959141808511_3
timestamp 1640697850
transform 0 1 3880 1 0 496
box -28 0 324 29
use sky130_fd_pr__nfet_01v8__example_55959141808509  sky130_fd_pr__nfet_01v8__example_55959141808509_0
timestamp 1640697850
transform 1 0 3349 0 1 1120
box -28 0 128 63
use sky130_fd_pr__nfet_01v8__example_55959141808509  sky130_fd_pr__nfet_01v8__example_55959141808509_1
timestamp 1640697850
transform -1 0 3918 0 -1 1270
box -28 0 128 63
use sky130_fd_pr__nfet_01v8__example_55959141808509  sky130_fd_pr__nfet_01v8__example_55959141808509_2
timestamp 1640697850
transform 1 0 3662 0 -1 1270
box -28 0 128 63
use sky130_fd_pr__nfet_01v8__example_55959141808503  sky130_fd_pr__nfet_01v8__example_55959141808503_0
timestamp 1640697850
transform 1 0 3347 0 1 1521
box -28 0 284 131
use sky130_fd_pr__nfet_01v8__example_55959141808485  sky130_fd_pr__nfet_01v8__example_55959141808485_0
timestamp 1640697850
transform 0 1 3798 1 0 1560
box -28 0 284 97
use sky130_fd_pr__nfet_01v8__example_55959141808485  sky130_fd_pr__nfet_01v8__example_55959141808485_1
timestamp 1640697850
transform 0 -1 3998 -1 0 2296
box -28 0 284 97
use sky130_fd_pr__nfet_01v8__example_55959141808474  sky130_fd_pr__nfet_01v8__example_55959141808474_0
timestamp 1640697850
transform 0 -1 3998 -1 0 2575
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808472  sky130_fd_pr__nfet_01v8__example_55959141808472_0
timestamp 1640697850
transform 1 0 22877 0 -1 2471
box -28 0 148 63
use sky130_fd_pr__nfet_01v8__example_55959141808472  sky130_fd_pr__nfet_01v8__example_55959141808472_1
timestamp 1640697850
transform -1 0 23173 0 -1 2471
box -28 0 148 63
use sky130_fd_pr__nfet_01v8__example_55959141808472  sky130_fd_pr__nfet_01v8__example_55959141808472_2
timestamp 1640697850
transform -1 0 22945 0 1 1336
box -28 0 148 63
use sky130_fd_pr__nfet_01v8__example_55959141808472  sky130_fd_pr__nfet_01v8__example_55959141808472_3
timestamp 1640697850
transform -1 0 23701 0 1 1336
box -28 0 148 63
use sky130_fd_pr__pfet_01v8__example_55959141808470  sky130_fd_pr__pfet_01v8__example_55959141808470_0
timestamp 1640697850
transform 0 -1 6411 1 0 -184
box -28 0 324 97
use sky130_fd_pr__pfet_01v8__example_55959141808470  sky130_fd_pr__pfet_01v8__example_55959141808470_1
timestamp 1640697850
transform 0 -1 6411 1 0 168
box -28 0 324 97
use sky130_fd_pr__pfet_01v8__example_55959141808470  sky130_fd_pr__pfet_01v8__example_55959141808470_2
timestamp 1640697850
transform 0 1 5258 1 0 -184
box -28 0 324 97
use sky130_fd_pr__pfet_01v8__example_55959141808470  sky130_fd_pr__pfet_01v8__example_55959141808470_3
timestamp 1640697850
transform 0 1 5258 1 0 168
box -28 0 324 97
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_0
timestamp 1640697850
transform 0 1 6626 1 0 233
box -28 0 128 131
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_1
timestamp 1640697850
transform 0 1 6626 1 0 -47
box -28 0 128 131
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_2
timestamp 1640697850
transform 0 1 6626 -1 0 -103
box -28 0 128 131
use sky130_fd_pr__pfet_01v8__example_55959141808508  sky130_fd_pr__pfet_01v8__example_55959141808508_0
timestamp 1640697850
transform 0 1 7385 -1 0 206
box -28 0 428 63
use sky130_fd_pr__pfet_01v8__example_55959141808508  sky130_fd_pr__pfet_01v8__example_55959141808508_1
timestamp 1640697850
transform 0 1 7105 -1 0 206
box -28 0 428 63
use sky130_fd_pr__pfet_01v8__example_55959141808469  sky130_fd_pr__pfet_01v8__example_55959141808469_0
timestamp 1640697850
transform -1 0 22997 0 1 1959
box -28 0 324 97
use sky130_fd_pr__pfet_01v8__example_55959141808469  sky130_fd_pr__pfet_01v8__example_55959141808469_1
timestamp 1640697850
transform 1 0 23053 0 1 1959
box -28 0 324 97
use sky130_fd_pr__pfet_01v8__example_55959141808507  sky130_fd_pr__pfet_01v8__example_55959141808507_0
timestamp 1640697850
transform 1 0 23405 0 1 1647
box -130 0 324 97
use sky130_fd_pr__pfet_01v8__example_55959141808505  sky130_fd_pr__pfet_01v8__example_55959141808505_0
timestamp 1640697850
transform 1 0 22825 0 1 1647
box -28 0 450 97
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_0
timestamp 1640697850
transform -1 0 16550 0 -1 865
box 0 24 534 1116
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_1
timestamp 1640697850
transform -1 0 16902 0 -1 865
box 0 24 534 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1640697850
transform 1 0 16720 0 -1 865
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1640697850
transform -1 0 16198 0 -1 865
box -46 24 399 1116
use sky130_fd_io__gpio_ovtv2_amux_drvr_ls_2  sky130_fd_io__gpio_ovtv2_amux_drvr_ls_2_0
timestamp 1640697850
transform 1 0 2826 0 1 51
box -31 -4 3247 2661
use sky130_fd_io__gpio_ovtv2_amux_guardring  sky130_fd_io__gpio_ovtv2_amux_guardring_0
timestamp 1640697850
transform 1 0 -142 0 1 -188
box -120 -120 4512 3350
use sky130_fd_io__gpio_ovtv2_amux_drvr_ls_i2c_fix_3  sky130_fd_io__gpio_ovtv2_amux_drvr_ls_i2c_fix_3_0
timestamp 1640697850
transform -1 0 21208 0 -1 2725
box 32 -167 1862 1132
use sky130_fd_io__gpio_ovtv2_amux_drvr_ls_i2c_fix_3  sky130_fd_io__gpio_ovtv2_amux_drvr_ls_i2c_fix_3_1
timestamp 1640697850
transform 1 0 17440 0 -1 2725
box 32 -167 1862 1132
use sky130_fd_io__gpio_ovtv2_amux_inv4_i2c_fix  sky130_fd_io__gpio_ovtv2_amux_inv4_i2c_fix_0
timestamp 1640697850
transform -1 0 22586 0 1 1099
box 50 -8 584 869
use sky130_fd_io__gpio_ovtv2_amux_inv4_i2c_fix  sky130_fd_io__gpio_ovtv2_amux_inv4_i2c_fix_1
timestamp 1640697850
transform -1 0 22234 0 1 1099
box 50 -8 584 869
use sky130_fd_io__gpio_ovtv2_amux_drvr_ls_i2c_fix_4  sky130_fd_io__gpio_ovtv2_amux_drvr_ls_i2c_fix_4_0
timestamp 1640697850
transform 1 0 17440 0 1 533
box 13 -167 1862 1138
use sky130_fd_io__gpio_ovtv2_amx_pucsd_buf_i2c_fix  sky130_fd_io__gpio_ovtv2_amx_pucsd_buf_i2c_fix_0
timestamp 1640697850
transform 1 0 21239 0 1 1876
box 1 -294 1490 797
<< labels >>
flabel metal2 s 4632 617 4732 667 3 FreeSans 400 0 0 0 NGB_AMX_VSWITCH_H
port 1 nsew
flabel metal2 s 4078 787 4159 839 3 FreeSans 400 0 0 0 NGB_PAD_VSWITCH_H
port 2 nsew
flabel metal2 s 4072 951 4160 1003 3 FreeSans 400 0 0 0 NGB_PAD_VSWITCH_H_N
port 3 nsew
flabel metal2 s 4629 264 4718 316 3 FreeSans 400 0 0 0 NGA_AMX_VSWITCH_H
port 4 nsew
flabel metal2 s 4642 705 4734 754 3 FreeSans 400 0 0 0 NGA_PAD_VSWITCH_H
port 5 nsew
flabel metal2 s 4629 181 4718 230 3 FreeSans 400 0 0 0 NGA_PAD_VSWITCH_H_N
port 6 nsew
flabel metal2 s 4629 92 4717 144 3 FreeSans 400 0 0 0 PD_CSD_VSWITCH_H
port 7 nsew
flabel metal2 s 4628 10 4711 62 3 FreeSans 400 0 0 0 PD_CSD_VSWITCH_H_N
port 8 nsew
flabel metal2 s 6593 2584 6692 2633 3 FreeSans 400 0 0 0 AMUXBUSA_ON
port 9 nsew
flabel metal2 s 6596 2499 6681 2549 3 FreeSans 400 0 0 0 AMUXBUSA_ON_N
port 10 nsew
flabel metal2 s 6589 2349 6683 2387 3 FreeSans 400 0 0 0 AMUXBUSB_ON
port 11 nsew
flabel metal2 s 6596 2417 6682 2466 3 FreeSans 400 0 0 0 AMUXBUSB_ON_N
port 12 nsew
flabel metal2 s 9566 2673 9647 2725 3 FreeSans 400 0 0 0 PD_ON
port 13 nsew
flabel metal2 s 9574 2755 9652 2798 3 FreeSans 400 0 0 0 PD_ON_N
port 14 nsew
flabel metal2 s 16264 450 16301 495 3 FreeSans 400 90 0 0 NMIDA_VCCD
port 15 nsew
flabel metal2 s 15756 708 15798 742 3 FreeSans 400 0 0 0 NMIDA_VCCD_N
port 16 nsew
flabel metal2 s 16622 363 16646 403 3 FreeSans 400 90 0 0 D_B
port 17 nsew
flabel metal2 s 15756 772 15798 806 3 FreeSans 400 0 0 0 D_B
port 17 nsew
flabel metal2 s 875 1609 918 1642 3 FreeSans 400 0 0 0 AMUX_EN_VDDA_H_N
port 18 nsew
flabel metal2 s 21745 733 21788 769 3 FreeSans 400 0 0 0 VSSD
port 19 nsew
flabel metal1 s 1262 1934 1308 1980 3 FreeSans 400 90 0 0 AMUX_EN_VSWITCH_H_N
port 20 nsew
flabel metal1 s 2255 88 2297 144 3 FreeSans 400 90 0 0 AMUX_EN_VSWITCH_H
port 21 nsew
flabel metal1 s 18915 -23 18991 29 3 FreeSans 400 0 0 0 AMUX_EN_VDDIO_H
port 22 nsew
flabel metal1 s -31 2105 2 2150 3 FreeSans 400 90 0 0 AMUX_EN_VDDA_H
port 23 nsew
flabel metal1 s 16175 320 16203 363 3 FreeSans 400 90 0 0 NMIDA_ON_N
port 24 nsew
flabel metal1 s 16523 192 16558 241 3 FreeSans 400 90 0 0 D_B
port 17 nsew
flabel metal1 s 20746 2462 20780 2509 3 FreeSans 400 90 0 0 PU_ON
port 25 nsew
flabel metal1 s 20898 2467 20936 2509 3 FreeSans 400 90 0 0 PU_ON_N
port 26 nsew
flabel metal1 s 15873 -105 15915 -69 3 FreeSans 400 0 0 0 VCCD
port 27 nsew
flabel metal1 s 5278 1973 5313 2013 3 FreeSans 400 90 0 0 VDDA
port 28 nsew
flabel metal1 s 21309 1749 21347 1789 3 FreeSans 400 90 0 0 VDDIO_Q
port 29 nsew
flabel metal1 s 798 1437 834 1476 3 FreeSans 400 90 0 0 VSSA
port 30 nsew
flabel metal1 s 6839 475 6878 515 3 FreeSans 400 0 0 0 VSWITCH
port 31 nsew
flabel metal1 s 978 2629 1024 2684 3 FreeSans 400 90 0 0 PGA_AMX_VDDA_H_N
port 32 nsew
flabel metal1 s 22246 1435 22290 1496 3 FreeSans 400 90 0 0 PGA_PAD_VDDIOQ_H_N
port 33 nsew
flabel metal1 s 890 1978 942 2040 3 FreeSans 400 90 0 0 PGB_AMX_VDDA_H_N
port 34 nsew
flabel metal1 s 21890 1452 21944 1515 3 FreeSans 400 90 0 0 PGB_PAD_VDDIOQ_H_N
port 35 nsew
flabel metal1 s 22360 2135 22413 2196 3 FreeSans 400 90 0 0 PU_CSD_VDDIOQ_H_N
port 36 nsew
flabel metal1 s 8208 1678 8244 1720 3 FreeSans 400 90 0 0 VCCD
port 27 nsew
flabel comment s 4307 650 4307 650 0 FreeSans 400 0 0 0 NGB_AMX_VSWITCH_H
flabel comment s 7845 817 7845 817 0 FreeSans 400 0 0 0 NGB_PAD_VSWITCH_H
flabel comment s 7843 901 7843 901 0 FreeSans 400 0 0 0 NGB_PAD_VSWITCH_H_N
flabel comment s 7846 734 7846 734 0 FreeSans 400 0 0 0 NGA_PAD_VSWITCH_H
flabel comment s 7838 217 7838 217 0 FreeSans 400 0 0 0 NGA_PAD_VSWITCH_H_N
flabel comment s 6856 126 6856 126 0 FreeSans 400 0 0 0 PD_CSD_VSWITCH_H
flabel comment s 7913 42 7913 42 0 FreeSans 400 0 0 0 PD_CSD_VSWITCH_H_N
flabel comment s 4040 1348 4040 1348 0 FreeSans 400 0 0 0 PD_CSD_VSWITCH_H
flabel comment s 7961 2370 7961 2370 0 FreeSans 400 0 0 0 AMUXBUSB_ON
flabel comment s 18507 3040 18507 3040 0 FreeSans 280 0 0 0 NET258(IN)
flabel comment s 9316 2782 9316 2782 0 FreeSans 400 0 0 0 PD_ON_N
flabel comment s 9328 2706 9328 2706 0 FreeSans 400 0 0 0 PD_ON
flabel comment s 7966 2523 7966 2523 0 FreeSans 400 0 0 0 AMUXBUSA_ON_N
flabel comment s 7960 2612 7960 2612 0 FreeSans 400 0 0 0 AMUXBUSA_ON
flabel comment s 7969 2446 7969 2446 0 FreeSans 400 0 0 0 AMUXBUSB_ON_N
flabel comment s 18518 3106 18518 3106 0 FreeSans 280 0 0 0 INB
flabel comment s 1171 2285 1171 2285 0 FreeSans 280 90 0 0 AMUX_EN_VDDA_H_N
flabel comment s 6 1631 6 1631 0 FreeSans 280 180 0 0 AMUX_EN_VDDA_H_N
flabel comment s 22432 2400 22432 2400 0 FreeSans 280 0 0 0 PU_CSD_VDDIOQ_H_N
flabel comment s 288 2771 288 2771 0 FreeSans 280 90 0 0 CONDIODE
flabel comment s 22651 1576 22651 1576 0 FreeSans 600 0 0 0 HLD_I_H_N
flabel comment s 18704 -3 18704 -3 0 FreeSans 280 0 0 0 AMUX_EN_VDDIO_H
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 48684136
string GDS_START 48538128
<< end >>
