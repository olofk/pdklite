magic
tech sky130A
magscale 1 2
timestamp 1640697977
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 827 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 315 47 345 177
rect 399 47 429 177
rect 515 47 545 177
rect 599 47 629 177
rect 705 47 735 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 315 297 345 497
rect 399 297 429 497
rect 515 297 545 497
rect 599 297 629 497
rect 705 297 735 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 161 163 177
rect 109 127 119 161
rect 153 127 163 161
rect 109 93 163 127
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 161 315 177
rect 193 127 235 161
rect 269 127 315 161
rect 193 93 315 127
rect 193 59 235 93
rect 269 59 315 93
rect 193 47 315 59
rect 345 161 399 177
rect 345 127 355 161
rect 389 127 399 161
rect 345 93 399 127
rect 345 59 355 93
rect 389 59 399 93
rect 345 47 399 59
rect 429 93 515 177
rect 429 59 455 93
rect 489 59 515 93
rect 429 47 515 59
rect 545 161 599 177
rect 545 127 555 161
rect 589 127 599 161
rect 545 93 599 127
rect 545 59 555 93
rect 589 59 599 93
rect 545 47 599 59
rect 629 161 705 177
rect 629 127 655 161
rect 689 127 705 161
rect 629 47 705 127
rect 735 161 801 177
rect 735 127 745 161
rect 779 127 801 161
rect 735 93 801 127
rect 735 59 745 93
rect 779 59 801 93
rect 735 47 801 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 475 315 497
rect 193 441 203 475
rect 237 441 271 475
rect 305 441 315 475
rect 193 297 315 441
rect 345 297 399 497
rect 429 297 515 497
rect 545 485 599 497
rect 545 451 555 485
rect 589 451 599 485
rect 545 417 599 451
rect 545 383 555 417
rect 589 383 599 417
rect 545 297 599 383
rect 629 297 705 497
rect 735 485 801 497
rect 735 451 745 485
rect 779 451 801 485
rect 735 417 801 451
rect 735 383 745 417
rect 779 383 801 417
rect 735 349 801 383
rect 735 315 745 349
rect 779 315 801 349
rect 735 297 801 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 127 153 161
rect 119 59 153 93
rect 235 127 269 161
rect 235 59 269 93
rect 355 127 389 161
rect 355 59 389 93
rect 455 59 489 93
rect 555 127 589 161
rect 555 59 589 93
rect 655 127 689 161
rect 745 127 779 161
rect 745 59 779 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 441 237 475
rect 271 441 305 475
rect 555 451 589 485
rect 555 383 589 417
rect 745 451 779 485
rect 745 383 779 417
rect 745 315 779 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 315 497 345 523
rect 399 497 429 523
rect 515 497 545 523
rect 599 497 629 523
rect 705 497 735 523
rect 79 265 109 297
rect 163 265 193 297
rect 315 265 345 297
rect 399 265 429 297
rect 515 265 545 297
rect 599 265 629 297
rect 79 249 247 265
rect 79 215 203 249
rect 237 215 247 249
rect 79 199 247 215
rect 289 249 345 265
rect 289 215 299 249
rect 333 215 345 249
rect 289 199 345 215
rect 387 249 441 265
rect 387 215 397 249
rect 431 215 441 249
rect 387 199 441 215
rect 483 249 545 265
rect 483 215 493 249
rect 527 215 545 249
rect 483 199 545 215
rect 587 249 641 265
rect 587 215 597 249
rect 631 215 641 249
rect 587 199 641 215
rect 705 261 735 297
rect 705 249 807 261
rect 705 215 755 249
rect 789 215 807 249
rect 705 203 807 215
rect 79 177 109 199
rect 163 177 193 199
rect 315 177 345 199
rect 399 177 429 199
rect 515 177 545 199
rect 599 177 629 199
rect 705 177 735 203
rect 79 21 109 47
rect 163 21 193 47
rect 315 21 345 47
rect 399 21 429 47
rect 515 21 545 47
rect 599 21 629 47
rect 705 21 735 47
<< polycont >>
rect 203 215 237 249
rect 299 215 333 249
rect 397 215 431 249
rect 493 215 527 249
rect 597 215 631 249
rect 755 215 789 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 485 69 527
rect 17 451 35 485
rect 17 417 69 451
rect 17 383 35 417
rect 17 349 69 383
rect 17 315 35 349
rect 17 299 69 315
rect 103 485 169 493
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 203 475 305 527
rect 237 441 271 475
rect 203 425 305 441
rect 539 485 605 493
rect 539 451 555 485
rect 589 451 605 485
rect 103 383 119 417
rect 153 383 169 417
rect 539 417 605 451
rect 539 391 555 417
rect 103 349 169 383
rect 103 315 119 349
rect 153 315 169 349
rect 17 161 69 177
rect 17 127 35 161
rect 17 93 69 127
rect 17 59 35 93
rect 17 17 69 59
rect 103 161 169 315
rect 203 383 555 391
rect 589 391 605 417
rect 739 485 811 527
rect 739 451 745 485
rect 779 451 811 485
rect 739 417 811 451
rect 589 383 705 391
rect 203 357 705 383
rect 203 249 265 357
rect 237 215 265 249
rect 203 199 265 215
rect 299 249 343 323
rect 333 215 343 249
rect 299 199 343 215
rect 397 249 432 323
rect 431 215 432 249
rect 397 199 432 215
rect 483 249 527 323
rect 483 215 493 249
rect 483 199 527 215
rect 582 249 631 323
rect 582 215 597 249
rect 582 199 631 215
rect 665 165 705 357
rect 739 383 745 417
rect 779 383 811 417
rect 739 349 811 383
rect 739 315 745 349
rect 779 315 811 349
rect 739 299 811 315
rect 745 249 811 265
rect 739 215 755 249
rect 789 215 811 249
rect 103 127 119 161
rect 153 127 169 161
rect 103 93 169 127
rect 103 59 119 93
rect 153 59 169 93
rect 103 51 169 59
rect 219 161 285 165
rect 219 127 235 161
rect 269 127 285 161
rect 219 93 285 127
rect 219 59 235 93
rect 269 59 285 93
rect 219 17 285 59
rect 339 161 605 165
rect 339 127 355 161
rect 389 131 555 161
rect 389 127 405 131
rect 339 93 405 127
rect 539 127 555 131
rect 589 127 605 161
rect 339 59 355 93
rect 389 59 405 93
rect 339 51 405 59
rect 439 93 505 97
rect 439 59 455 93
rect 489 59 505 93
rect 439 17 505 59
rect 539 93 605 127
rect 639 161 705 165
rect 639 127 655 161
rect 689 127 705 161
rect 639 119 705 127
rect 739 161 811 181
rect 739 127 745 161
rect 779 127 811 161
rect 539 59 555 93
rect 589 85 605 93
rect 739 93 811 127
rect 739 85 745 93
rect 589 59 745 85
rect 779 59 811 93
rect 539 51 811 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 766 221 800 255 0 FreeSans 250 0 0 0 B1
port 4 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 250 0 0 0 B2
port 5 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 122 85 156 119 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel locali s 122 153 156 187 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel locali s 122 289 156 323 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel locali s 122 357 156 391 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel locali s 122 425 156 459 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o32a_2
rlabel metal1 s 0 -48 828 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 1487078
string GDS_START 1479344
string path 0.000 0.000 4.140 0.000 
<< end >>
