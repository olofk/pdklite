magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1239 -1236 1373 1288
<< labels >>
flabel comment s 50 27 50 27 0 FreeSans 50 0 0 0 A
flabel comment s 86 27 86 27 0 FreeSans 50 0 0 0 B
flabel comment s 59 25 59 25 2 FreeSans 50 0 0 0 EM1S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 39964234
string GDS_START 39963530
<< end >>
