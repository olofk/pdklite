magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect 24595 -17719 43320 3236
<< nwell >>
rect 25915 1200 26081 1914
rect 26557 1200 27193 1316
rect 25915 1131 27193 1200
rect 25974 1090 27193 1131
<< pwell >>
rect 27322 -992 28068 -696
rect 28699 -992 29757 -696
rect 27573 -1740 27847 -1119
rect 28088 -3500 28368 -2914
<< psubdiff >>
rect 27322 -698 28068 -696
rect 27322 -732 27346 -698
rect 27380 -732 27420 -698
rect 27454 -732 27494 -698
rect 27528 -732 27568 -698
rect 27602 -732 27642 -698
rect 27676 -732 27716 -698
rect 27750 -732 27790 -698
rect 27824 -732 27864 -698
rect 27898 -732 27937 -698
rect 27971 -732 28010 -698
rect 28044 -732 28068 -698
rect 27322 -784 28068 -732
rect 27322 -818 27346 -784
rect 27380 -818 27420 -784
rect 27454 -818 27494 -784
rect 27528 -818 27568 -784
rect 27602 -818 27642 -784
rect 27676 -818 27716 -784
rect 27750 -818 27790 -784
rect 27824 -818 27864 -784
rect 27898 -818 27937 -784
rect 27971 -818 28010 -784
rect 28044 -818 28068 -784
rect 27322 -870 28068 -818
rect 27322 -904 27346 -870
rect 27380 -904 27420 -870
rect 27454 -904 27494 -870
rect 27528 -904 27568 -870
rect 27602 -904 27642 -870
rect 27676 -904 27716 -870
rect 27750 -904 27790 -870
rect 27824 -904 27864 -870
rect 27898 -904 27937 -870
rect 27971 -904 28010 -870
rect 28044 -904 28068 -870
rect 27322 -956 28068 -904
rect 27322 -990 27346 -956
rect 27380 -990 27420 -956
rect 27454 -990 27494 -956
rect 27528 -990 27568 -956
rect 27602 -990 27642 -956
rect 27676 -990 27716 -956
rect 27750 -990 27790 -956
rect 27824 -990 27864 -956
rect 27898 -990 27937 -956
rect 27971 -990 28010 -956
rect 28044 -990 28068 -956
rect 27322 -992 28068 -990
rect 28699 -698 29757 -696
rect 28699 -732 28723 -698
rect 28757 -732 28793 -698
rect 28827 -732 28863 -698
rect 28897 -732 28933 -698
rect 28967 -732 29003 -698
rect 29037 -732 29073 -698
rect 29107 -732 29143 -698
rect 29177 -732 29213 -698
rect 29247 -732 29283 -698
rect 29317 -732 29353 -698
rect 29387 -732 29423 -698
rect 29457 -732 29492 -698
rect 29526 -732 29561 -698
rect 29595 -732 29630 -698
rect 29664 -732 29699 -698
rect 29733 -732 29757 -698
rect 28699 -784 29757 -732
rect 28699 -818 28723 -784
rect 28757 -818 28793 -784
rect 28827 -818 28863 -784
rect 28897 -818 28933 -784
rect 28967 -818 29003 -784
rect 29037 -818 29073 -784
rect 29107 -818 29143 -784
rect 29177 -818 29213 -784
rect 29247 -818 29283 -784
rect 29317 -818 29353 -784
rect 29387 -818 29423 -784
rect 29457 -818 29492 -784
rect 29526 -818 29561 -784
rect 29595 -818 29630 -784
rect 29664 -818 29699 -784
rect 29733 -818 29757 -784
rect 28699 -870 29757 -818
rect 28699 -904 28723 -870
rect 28757 -904 28793 -870
rect 28827 -904 28863 -870
rect 28897 -904 28933 -870
rect 28967 -904 29003 -870
rect 29037 -904 29073 -870
rect 29107 -904 29143 -870
rect 29177 -904 29213 -870
rect 29247 -904 29283 -870
rect 29317 -904 29353 -870
rect 29387 -904 29423 -870
rect 29457 -904 29492 -870
rect 29526 -904 29561 -870
rect 29595 -904 29630 -870
rect 29664 -904 29699 -870
rect 29733 -904 29757 -870
rect 28699 -956 29757 -904
rect 28699 -990 28723 -956
rect 28757 -990 28793 -956
rect 28827 -990 28863 -956
rect 28897 -990 28933 -956
rect 28967 -990 29003 -956
rect 29037 -990 29073 -956
rect 29107 -990 29143 -956
rect 29177 -990 29213 -956
rect 29247 -990 29283 -956
rect 29317 -990 29353 -956
rect 29387 -990 29423 -956
rect 29457 -990 29492 -956
rect 29526 -990 29561 -956
rect 29595 -990 29630 -956
rect 29664 -990 29699 -956
rect 29733 -990 29757 -956
rect 28699 -992 29757 -990
rect 27573 -1143 27847 -1119
rect 27607 -1177 27653 -1143
rect 27687 -1177 27733 -1143
rect 27767 -1177 27813 -1143
rect 27573 -1220 27847 -1177
rect 27607 -1254 27653 -1220
rect 27687 -1254 27733 -1220
rect 27767 -1254 27813 -1220
rect 27573 -1297 27847 -1254
rect 27607 -1331 27653 -1297
rect 27687 -1331 27733 -1297
rect 27767 -1331 27813 -1297
rect 27573 -1374 27847 -1331
rect 27607 -1408 27653 -1374
rect 27687 -1408 27733 -1374
rect 27767 -1408 27813 -1374
rect 27573 -1451 27847 -1408
rect 27607 -1485 27653 -1451
rect 27687 -1485 27733 -1451
rect 27767 -1485 27813 -1451
rect 27573 -1528 27847 -1485
rect 27607 -1562 27653 -1528
rect 27687 -1562 27733 -1528
rect 27767 -1562 27813 -1528
rect 27573 -1605 27847 -1562
rect 27607 -1639 27653 -1605
rect 27687 -1639 27733 -1605
rect 27767 -1639 27813 -1605
rect 27573 -1682 27847 -1639
rect 27607 -1716 27653 -1682
rect 27687 -1716 27733 -1682
rect 27767 -1716 27813 -1682
rect 27573 -1740 27847 -1716
rect 28088 -2948 28368 -2914
rect 28122 -2982 28170 -2948
rect 28204 -2982 28252 -2948
rect 28286 -2982 28334 -2948
rect 28088 -3017 28368 -2982
rect 28122 -3051 28170 -3017
rect 28204 -3051 28252 -3017
rect 28286 -3051 28334 -3017
rect 28088 -3086 28368 -3051
rect 28122 -3120 28170 -3086
rect 28204 -3120 28252 -3086
rect 28286 -3120 28334 -3086
rect 28088 -3155 28368 -3120
rect 28122 -3189 28170 -3155
rect 28204 -3189 28252 -3155
rect 28286 -3189 28334 -3155
rect 28088 -3224 28368 -3189
rect 28122 -3258 28170 -3224
rect 28204 -3258 28252 -3224
rect 28286 -3258 28334 -3224
rect 28088 -3293 28368 -3258
rect 28122 -3327 28170 -3293
rect 28204 -3327 28252 -3293
rect 28286 -3327 28334 -3293
rect 28088 -3362 28368 -3327
rect 28122 -3396 28170 -3362
rect 28204 -3396 28252 -3362
rect 28286 -3396 28334 -3362
rect 28088 -3432 28368 -3396
rect 28122 -3466 28170 -3432
rect 28204 -3466 28252 -3432
rect 28286 -3466 28334 -3432
rect 28088 -3500 28368 -3466
<< mvnsubdiff >>
rect 25981 1824 26015 1848
rect 25981 1753 26015 1790
rect 25981 1682 26015 1719
rect 25981 1611 26015 1648
rect 25981 1540 26015 1577
rect 25981 1469 26015 1506
rect 25981 1398 26015 1435
rect 25981 1327 26015 1364
rect 25981 1255 26015 1293
rect 25981 1197 26015 1221
<< psubdiffcont >>
rect 27346 -732 27380 -698
rect 27420 -732 27454 -698
rect 27494 -732 27528 -698
rect 27568 -732 27602 -698
rect 27642 -732 27676 -698
rect 27716 -732 27750 -698
rect 27790 -732 27824 -698
rect 27864 -732 27898 -698
rect 27937 -732 27971 -698
rect 28010 -732 28044 -698
rect 27346 -818 27380 -784
rect 27420 -818 27454 -784
rect 27494 -818 27528 -784
rect 27568 -818 27602 -784
rect 27642 -818 27676 -784
rect 27716 -818 27750 -784
rect 27790 -818 27824 -784
rect 27864 -818 27898 -784
rect 27937 -818 27971 -784
rect 28010 -818 28044 -784
rect 27346 -904 27380 -870
rect 27420 -904 27454 -870
rect 27494 -904 27528 -870
rect 27568 -904 27602 -870
rect 27642 -904 27676 -870
rect 27716 -904 27750 -870
rect 27790 -904 27824 -870
rect 27864 -904 27898 -870
rect 27937 -904 27971 -870
rect 28010 -904 28044 -870
rect 27346 -990 27380 -956
rect 27420 -990 27454 -956
rect 27494 -990 27528 -956
rect 27568 -990 27602 -956
rect 27642 -990 27676 -956
rect 27716 -990 27750 -956
rect 27790 -990 27824 -956
rect 27864 -990 27898 -956
rect 27937 -990 27971 -956
rect 28010 -990 28044 -956
rect 28723 -732 28757 -698
rect 28793 -732 28827 -698
rect 28863 -732 28897 -698
rect 28933 -732 28967 -698
rect 29003 -732 29037 -698
rect 29073 -732 29107 -698
rect 29143 -732 29177 -698
rect 29213 -732 29247 -698
rect 29283 -732 29317 -698
rect 29353 -732 29387 -698
rect 29423 -732 29457 -698
rect 29492 -732 29526 -698
rect 29561 -732 29595 -698
rect 29630 -732 29664 -698
rect 29699 -732 29733 -698
rect 28723 -818 28757 -784
rect 28793 -818 28827 -784
rect 28863 -818 28897 -784
rect 28933 -818 28967 -784
rect 29003 -818 29037 -784
rect 29073 -818 29107 -784
rect 29143 -818 29177 -784
rect 29213 -818 29247 -784
rect 29283 -818 29317 -784
rect 29353 -818 29387 -784
rect 29423 -818 29457 -784
rect 29492 -818 29526 -784
rect 29561 -818 29595 -784
rect 29630 -818 29664 -784
rect 29699 -818 29733 -784
rect 28723 -904 28757 -870
rect 28793 -904 28827 -870
rect 28863 -904 28897 -870
rect 28933 -904 28967 -870
rect 29003 -904 29037 -870
rect 29073 -904 29107 -870
rect 29143 -904 29177 -870
rect 29213 -904 29247 -870
rect 29283 -904 29317 -870
rect 29353 -904 29387 -870
rect 29423 -904 29457 -870
rect 29492 -904 29526 -870
rect 29561 -904 29595 -870
rect 29630 -904 29664 -870
rect 29699 -904 29733 -870
rect 28723 -990 28757 -956
rect 28793 -990 28827 -956
rect 28863 -990 28897 -956
rect 28933 -990 28967 -956
rect 29003 -990 29037 -956
rect 29073 -990 29107 -956
rect 29143 -990 29177 -956
rect 29213 -990 29247 -956
rect 29283 -990 29317 -956
rect 29353 -990 29387 -956
rect 29423 -990 29457 -956
rect 29492 -990 29526 -956
rect 29561 -990 29595 -956
rect 29630 -990 29664 -956
rect 29699 -990 29733 -956
rect 27573 -1177 27607 -1143
rect 27653 -1177 27687 -1143
rect 27733 -1177 27767 -1143
rect 27813 -1177 27847 -1143
rect 27573 -1254 27607 -1220
rect 27653 -1254 27687 -1220
rect 27733 -1254 27767 -1220
rect 27813 -1254 27847 -1220
rect 27573 -1331 27607 -1297
rect 27653 -1331 27687 -1297
rect 27733 -1331 27767 -1297
rect 27813 -1331 27847 -1297
rect 27573 -1408 27607 -1374
rect 27653 -1408 27687 -1374
rect 27733 -1408 27767 -1374
rect 27813 -1408 27847 -1374
rect 27573 -1485 27607 -1451
rect 27653 -1485 27687 -1451
rect 27733 -1485 27767 -1451
rect 27813 -1485 27847 -1451
rect 27573 -1562 27607 -1528
rect 27653 -1562 27687 -1528
rect 27733 -1562 27767 -1528
rect 27813 -1562 27847 -1528
rect 27573 -1639 27607 -1605
rect 27653 -1639 27687 -1605
rect 27733 -1639 27767 -1605
rect 27813 -1639 27847 -1605
rect 27573 -1716 27607 -1682
rect 27653 -1716 27687 -1682
rect 27733 -1716 27767 -1682
rect 27813 -1716 27847 -1682
rect 28088 -2982 28122 -2948
rect 28170 -2982 28204 -2948
rect 28252 -2982 28286 -2948
rect 28334 -2982 28368 -2948
rect 28088 -3051 28122 -3017
rect 28170 -3051 28204 -3017
rect 28252 -3051 28286 -3017
rect 28334 -3051 28368 -3017
rect 28088 -3120 28122 -3086
rect 28170 -3120 28204 -3086
rect 28252 -3120 28286 -3086
rect 28334 -3120 28368 -3086
rect 28088 -3189 28122 -3155
rect 28170 -3189 28204 -3155
rect 28252 -3189 28286 -3155
rect 28334 -3189 28368 -3155
rect 28088 -3258 28122 -3224
rect 28170 -3258 28204 -3224
rect 28252 -3258 28286 -3224
rect 28334 -3258 28368 -3224
rect 28088 -3327 28122 -3293
rect 28170 -3327 28204 -3293
rect 28252 -3327 28286 -3293
rect 28334 -3327 28368 -3293
rect 28088 -3396 28122 -3362
rect 28170 -3396 28204 -3362
rect 28252 -3396 28286 -3362
rect 28334 -3396 28368 -3362
rect 28088 -3466 28122 -3432
rect 28170 -3466 28204 -3432
rect 28252 -3466 28286 -3432
rect 28334 -3466 28368 -3432
<< mvnsubdiffcont >>
rect 25981 1790 26015 1824
rect 25981 1719 26015 1753
rect 25981 1648 26015 1682
rect 25981 1577 26015 1611
rect 25981 1506 26015 1540
rect 25981 1435 26015 1469
rect 25981 1364 26015 1398
rect 25981 1293 26015 1327
rect 25981 1221 26015 1255
<< locali >>
rect 25981 1824 26015 1848
rect 25981 1753 26015 1790
rect 25981 1718 26015 1719
rect 25981 1682 26015 1684
rect 25981 1646 26015 1648
rect 25981 1611 26015 1612
rect 25981 1574 26015 1577
rect 25981 1502 26015 1506
rect 25981 1430 26015 1435
rect 25981 1327 26015 1364
rect 25981 1255 26015 1293
rect 25981 1197 26015 1221
rect 27322 -698 28068 -696
rect 27322 -732 27346 -698
rect 27380 -732 27420 -698
rect 27454 -732 27494 -698
rect 27528 -732 27568 -698
rect 27602 -732 27642 -698
rect 27676 -732 27716 -698
rect 27750 -732 27790 -698
rect 27824 -732 27864 -698
rect 27898 -732 27937 -698
rect 27971 -732 28010 -698
rect 28044 -732 28068 -698
rect 27322 -784 28068 -732
rect 27322 -818 27346 -784
rect 27380 -818 27420 -784
rect 27454 -818 27494 -784
rect 27528 -818 27568 -784
rect 27602 -818 27642 -784
rect 27676 -818 27716 -784
rect 27750 -818 27790 -784
rect 27824 -818 27864 -784
rect 27898 -818 27937 -784
rect 27971 -818 28010 -784
rect 28044 -818 28068 -784
rect 27322 -856 28068 -818
rect 27322 -890 27339 -856
rect 27373 -870 27414 -856
rect 27448 -870 27489 -856
rect 27523 -870 27564 -856
rect 27598 -870 27639 -856
rect 27673 -870 27714 -856
rect 27748 -870 27789 -856
rect 27823 -870 27864 -856
rect 27898 -870 27939 -856
rect 27973 -870 28013 -856
rect 27380 -890 27414 -870
rect 27454 -890 27489 -870
rect 27528 -890 27564 -870
rect 27602 -890 27639 -870
rect 27676 -890 27714 -870
rect 27750 -890 27789 -870
rect 27322 -904 27346 -890
rect 27380 -904 27420 -890
rect 27454 -904 27494 -890
rect 27528 -904 27568 -890
rect 27602 -904 27642 -890
rect 27676 -904 27716 -890
rect 27750 -904 27790 -890
rect 27824 -904 27864 -870
rect 27898 -904 27937 -870
rect 27973 -890 28010 -870
rect 28047 -890 28068 -856
rect 27971 -904 28010 -890
rect 28044 -904 28068 -890
rect 27322 -956 28068 -904
rect 27322 -990 27346 -956
rect 27380 -990 27420 -956
rect 27454 -990 27494 -956
rect 27528 -990 27568 -956
rect 27602 -990 27642 -956
rect 27676 -990 27716 -956
rect 27750 -990 27790 -956
rect 27824 -990 27864 -956
rect 27898 -990 27937 -956
rect 27971 -990 28010 -956
rect 28044 -990 28068 -956
rect 27322 -992 28068 -990
rect 28699 -698 29757 -696
rect 28699 -732 28723 -698
rect 28757 -732 28793 -698
rect 28827 -699 28863 -698
rect 28897 -699 28933 -698
rect 28967 -699 29003 -698
rect 29037 -699 29073 -698
rect 29107 -699 29143 -698
rect 28830 -732 28863 -699
rect 28905 -732 28933 -699
rect 28980 -732 29003 -699
rect 29054 -732 29073 -699
rect 29128 -732 29143 -699
rect 29177 -732 29213 -698
rect 29247 -732 29283 -698
rect 29317 -732 29353 -698
rect 29387 -732 29423 -698
rect 29457 -732 29492 -698
rect 29526 -732 29561 -698
rect 29595 -732 29630 -698
rect 29664 -732 29699 -698
rect 29733 -732 29757 -698
rect 28699 -733 28796 -732
rect 28830 -733 28871 -732
rect 28905 -733 28946 -732
rect 28980 -733 29020 -732
rect 29054 -733 29094 -732
rect 29128 -733 29757 -732
rect 28699 -783 29757 -733
rect 28699 -784 28796 -783
rect 28830 -784 28871 -783
rect 28905 -784 28946 -783
rect 28980 -784 29020 -783
rect 29054 -784 29094 -783
rect 29128 -784 29757 -783
rect 28699 -818 28723 -784
rect 28757 -818 28793 -784
rect 28830 -817 28863 -784
rect 28905 -817 28933 -784
rect 28980 -817 29003 -784
rect 29054 -817 29073 -784
rect 29128 -817 29143 -784
rect 28827 -818 28863 -817
rect 28897 -818 28933 -817
rect 28967 -818 29003 -817
rect 29037 -818 29073 -817
rect 29107 -818 29143 -817
rect 29177 -818 29213 -784
rect 29247 -818 29283 -784
rect 29317 -818 29353 -784
rect 29387 -818 29423 -784
rect 29457 -818 29492 -784
rect 29526 -818 29561 -784
rect 29595 -818 29630 -784
rect 29664 -818 29699 -784
rect 29733 -818 29757 -784
rect 28699 -867 29757 -818
rect 28699 -870 28796 -867
rect 28830 -870 28871 -867
rect 28905 -870 28946 -867
rect 28980 -870 29020 -867
rect 29054 -870 29094 -867
rect 29128 -870 29757 -867
rect 28699 -904 28723 -870
rect 28757 -904 28793 -870
rect 28830 -901 28863 -870
rect 28905 -901 28933 -870
rect 28980 -901 29003 -870
rect 29054 -901 29073 -870
rect 29128 -901 29143 -870
rect 28827 -904 28863 -901
rect 28897 -904 28933 -901
rect 28967 -904 29003 -901
rect 29037 -904 29073 -901
rect 29107 -904 29143 -901
rect 29177 -904 29213 -870
rect 29247 -904 29283 -870
rect 29317 -904 29353 -870
rect 29387 -904 29423 -870
rect 29457 -904 29492 -870
rect 29526 -904 29561 -870
rect 29595 -904 29630 -870
rect 29664 -904 29699 -870
rect 29733 -904 29757 -870
rect 28699 -951 29757 -904
rect 28699 -956 28796 -951
rect 28830 -956 28871 -951
rect 28905 -956 28946 -951
rect 28980 -956 29020 -951
rect 29054 -956 29094 -951
rect 29128 -956 29757 -951
rect 28699 -990 28723 -956
rect 28757 -990 28793 -956
rect 28830 -985 28863 -956
rect 28905 -985 28933 -956
rect 28980 -985 29003 -956
rect 29054 -985 29073 -956
rect 29128 -985 29143 -956
rect 28827 -990 28863 -985
rect 28897 -990 28933 -985
rect 28967 -990 29003 -985
rect 29037 -990 29073 -985
rect 29107 -990 29143 -985
rect 29177 -990 29213 -956
rect 29247 -990 29283 -956
rect 29317 -990 29353 -956
rect 29387 -990 29423 -956
rect 29457 -990 29492 -956
rect 29526 -990 29561 -956
rect 29595 -990 29630 -956
rect 29664 -990 29699 -956
rect 29733 -990 29757 -956
rect 28699 -992 29757 -990
rect 27573 -1143 27847 -1119
rect 27607 -1164 27653 -1143
rect 27687 -1164 27733 -1143
rect 27767 -1164 27813 -1143
rect 27607 -1177 27652 -1164
rect 27687 -1177 27732 -1164
rect 27767 -1177 27811 -1164
rect 27606 -1198 27652 -1177
rect 27686 -1198 27732 -1177
rect 27766 -1198 27811 -1177
rect 27845 -1198 27847 -1177
rect 27572 -1220 27847 -1198
rect 27572 -1254 27573 -1220
rect 27607 -1254 27653 -1220
rect 27687 -1254 27733 -1220
rect 27767 -1254 27813 -1220
rect 27572 -1297 27847 -1254
rect 27572 -1304 27573 -1297
rect 27607 -1304 27653 -1297
rect 27687 -1304 27733 -1297
rect 27767 -1304 27813 -1297
rect 27607 -1331 27652 -1304
rect 27687 -1331 27732 -1304
rect 27767 -1331 27811 -1304
rect 27606 -1338 27652 -1331
rect 27686 -1338 27732 -1331
rect 27766 -1338 27811 -1331
rect 27845 -1338 27847 -1331
rect 27573 -1374 27847 -1338
rect 27607 -1408 27653 -1374
rect 27687 -1408 27733 -1374
rect 27767 -1408 27813 -1374
rect 27573 -1451 27847 -1408
rect 27607 -1485 27653 -1451
rect 27687 -1485 27733 -1451
rect 27767 -1485 27813 -1451
rect 27573 -1528 27847 -1485
rect 27607 -1562 27653 -1528
rect 27687 -1562 27733 -1528
rect 27767 -1562 27813 -1528
rect 27573 -1605 27847 -1562
rect 27607 -1639 27653 -1605
rect 27687 -1639 27733 -1605
rect 27767 -1639 27813 -1605
rect 27573 -1682 27847 -1639
rect 27607 -1685 27653 -1682
rect 27687 -1685 27733 -1682
rect 27767 -1685 27813 -1682
rect 27573 -1719 27578 -1716
rect 27612 -1719 27653 -1685
rect 27687 -1719 27728 -1685
rect 27767 -1716 27803 -1685
rect 27762 -1719 27803 -1716
rect 27837 -1719 27847 -1716
rect 27573 -1740 27847 -1719
rect 30266 -1890 30328 -1858
rect 30266 -1924 30280 -1890
rect 30314 -1924 30328 -1890
rect 30266 -1964 30328 -1924
rect 30266 -1998 30280 -1964
rect 30314 -1998 30328 -1964
rect 30266 -2039 30328 -1998
rect 30266 -2073 30280 -2039
rect 30314 -2073 30328 -2039
rect 30266 -2114 30328 -2073
rect 30266 -2148 30280 -2114
rect 30314 -2148 30328 -2114
rect 30266 -2180 30328 -2148
rect 30076 -2226 30124 -2192
rect 30158 -2226 30206 -2192
rect 30240 -2226 30288 -2192
rect 30042 -2267 30322 -2226
rect 30076 -2301 30124 -2267
rect 30158 -2301 30206 -2267
rect 30240 -2301 30288 -2267
rect 30042 -2342 30322 -2301
rect 30076 -2376 30124 -2342
rect 30158 -2376 30206 -2342
rect 30240 -2376 30288 -2342
rect 30042 -2417 30322 -2376
rect 30076 -2451 30124 -2417
rect 30158 -2451 30206 -2417
rect 30240 -2451 30288 -2417
rect 30042 -2493 30322 -2451
rect 30076 -2527 30124 -2493
rect 30158 -2527 30206 -2493
rect 30240 -2527 30288 -2493
rect 30042 -2569 30322 -2527
rect 30076 -2603 30124 -2569
rect 30158 -2603 30206 -2569
rect 30240 -2603 30288 -2569
rect 30042 -2645 30322 -2603
rect 30076 -2679 30124 -2645
rect 30158 -2679 30206 -2645
rect 30240 -2679 30288 -2645
rect 30042 -2721 30322 -2679
rect 30076 -2755 30124 -2721
rect 30158 -2755 30206 -2721
rect 30240 -2755 30288 -2721
rect 30042 -2797 30322 -2755
rect 30076 -2831 30124 -2797
rect 30158 -2831 30206 -2797
rect 30240 -2831 30288 -2797
rect 30042 -2873 30322 -2831
rect 30076 -2907 30124 -2873
rect 30158 -2907 30206 -2873
rect 30240 -2907 30288 -2873
rect 28088 -2945 28368 -2914
rect 28088 -2948 28098 -2945
rect 28132 -2948 28218 -2945
rect 28132 -2979 28170 -2948
rect 28122 -2982 28170 -2979
rect 28204 -2979 28218 -2948
rect 28252 -2948 28368 -2945
rect 28204 -2982 28252 -2979
rect 28286 -2982 28334 -2948
rect 28088 -3017 28368 -2982
rect 30042 -2949 30322 -2907
rect 30076 -2983 30124 -2949
rect 30158 -2983 30206 -2949
rect 30240 -2983 30288 -2949
rect 28122 -3022 28170 -3017
rect 28132 -3051 28170 -3022
rect 28204 -3022 28252 -3017
rect 28204 -3051 28218 -3022
rect 28088 -3056 28098 -3051
rect 28132 -3056 28218 -3051
rect 28286 -3051 28334 -3017
rect 28252 -3056 28368 -3051
rect 28088 -3086 28368 -3056
rect 28122 -3099 28170 -3086
rect 28132 -3120 28170 -3099
rect 28204 -3099 28252 -3086
rect 28204 -3120 28218 -3099
rect 28088 -3133 28098 -3120
rect 28132 -3133 28218 -3120
rect 28286 -3120 28334 -3086
rect 28252 -3133 28368 -3120
rect 28088 -3155 28368 -3133
rect 28122 -3176 28170 -3155
rect 28132 -3189 28170 -3176
rect 28204 -3176 28252 -3155
rect 28204 -3189 28218 -3176
rect 28088 -3210 28098 -3189
rect 28132 -3210 28218 -3189
rect 28286 -3189 28334 -3155
rect 28252 -3210 28368 -3189
rect 28088 -3224 28368 -3210
rect 28122 -3254 28170 -3224
rect 28132 -3258 28170 -3254
rect 28204 -3254 28252 -3224
rect 28204 -3258 28218 -3254
rect 28088 -3288 28098 -3258
rect 28132 -3288 28218 -3258
rect 28286 -3258 28334 -3224
rect 28252 -3288 28368 -3258
rect 28088 -3293 28368 -3288
rect 28122 -3327 28170 -3293
rect 28204 -3327 28252 -3293
rect 28286 -3327 28334 -3293
rect 28088 -3332 28368 -3327
rect 28088 -3362 28098 -3332
rect 28132 -3362 28218 -3332
rect 28132 -3366 28170 -3362
rect 28122 -3396 28170 -3366
rect 28204 -3366 28218 -3362
rect 28252 -3362 28368 -3332
rect 28204 -3396 28252 -3366
rect 28286 -3396 28334 -3362
rect 28088 -3410 28368 -3396
rect 28088 -3432 28098 -3410
rect 28132 -3432 28218 -3410
rect 28132 -3444 28170 -3432
rect 28122 -3466 28170 -3444
rect 28204 -3444 28218 -3432
rect 28252 -3432 28368 -3410
rect 28204 -3466 28252 -3444
rect 28286 -3466 28334 -3432
rect 28088 -3500 28368 -3466
rect 34118 -3909 34152 -3871
rect 32564 -4815 32629 -4496
rect 32751 -4815 32814 -4496
<< viali >>
rect 25981 1684 26015 1718
rect 25981 1612 26015 1646
rect 25981 1540 26015 1574
rect 25981 1469 26015 1502
rect 25981 1468 26015 1469
rect 25981 1398 26015 1430
rect 25981 1396 26015 1398
rect 27339 -870 27373 -856
rect 27414 -870 27448 -856
rect 27489 -870 27523 -856
rect 27564 -870 27598 -856
rect 27639 -870 27673 -856
rect 27714 -870 27748 -856
rect 27789 -870 27823 -856
rect 27864 -870 27898 -856
rect 27939 -870 27973 -856
rect 28013 -870 28047 -856
rect 27339 -890 27346 -870
rect 27346 -890 27373 -870
rect 27414 -890 27420 -870
rect 27420 -890 27448 -870
rect 27489 -890 27494 -870
rect 27494 -890 27523 -870
rect 27564 -890 27568 -870
rect 27568 -890 27598 -870
rect 27639 -890 27642 -870
rect 27642 -890 27673 -870
rect 27714 -890 27716 -870
rect 27716 -890 27748 -870
rect 27789 -890 27790 -870
rect 27790 -890 27823 -870
rect 27864 -890 27898 -870
rect 27939 -890 27971 -870
rect 27971 -890 27973 -870
rect 28013 -890 28044 -870
rect 28044 -890 28047 -870
rect 28796 -732 28827 -699
rect 28827 -732 28830 -699
rect 28871 -732 28897 -699
rect 28897 -732 28905 -699
rect 28946 -732 28967 -699
rect 28967 -732 28980 -699
rect 29020 -732 29037 -699
rect 29037 -732 29054 -699
rect 29094 -732 29107 -699
rect 29107 -732 29128 -699
rect 28796 -733 28830 -732
rect 28871 -733 28905 -732
rect 28946 -733 28980 -732
rect 29020 -733 29054 -732
rect 29094 -733 29128 -732
rect 28796 -784 28830 -783
rect 28871 -784 28905 -783
rect 28946 -784 28980 -783
rect 29020 -784 29054 -783
rect 29094 -784 29128 -783
rect 28796 -817 28827 -784
rect 28827 -817 28830 -784
rect 28871 -817 28897 -784
rect 28897 -817 28905 -784
rect 28946 -817 28967 -784
rect 28967 -817 28980 -784
rect 29020 -817 29037 -784
rect 29037 -817 29054 -784
rect 29094 -817 29107 -784
rect 29107 -817 29128 -784
rect 28796 -870 28830 -867
rect 28871 -870 28905 -867
rect 28946 -870 28980 -867
rect 29020 -870 29054 -867
rect 29094 -870 29128 -867
rect 28796 -901 28827 -870
rect 28827 -901 28830 -870
rect 28871 -901 28897 -870
rect 28897 -901 28905 -870
rect 28946 -901 28967 -870
rect 28967 -901 28980 -870
rect 29020 -901 29037 -870
rect 29037 -901 29054 -870
rect 29094 -901 29107 -870
rect 29107 -901 29128 -870
rect 28796 -956 28830 -951
rect 28871 -956 28905 -951
rect 28946 -956 28980 -951
rect 29020 -956 29054 -951
rect 29094 -956 29128 -951
rect 28796 -985 28827 -956
rect 28827 -985 28830 -956
rect 28871 -985 28897 -956
rect 28897 -985 28905 -956
rect 28946 -985 28967 -956
rect 28967 -985 28980 -956
rect 29020 -985 29037 -956
rect 29037 -985 29054 -956
rect 29094 -985 29107 -956
rect 29107 -985 29128 -956
rect 27572 -1177 27573 -1164
rect 27573 -1177 27606 -1164
rect 27652 -1177 27653 -1164
rect 27653 -1177 27686 -1164
rect 27732 -1177 27733 -1164
rect 27733 -1177 27766 -1164
rect 27811 -1177 27813 -1164
rect 27813 -1177 27845 -1164
rect 27572 -1198 27606 -1177
rect 27652 -1198 27686 -1177
rect 27732 -1198 27766 -1177
rect 27811 -1198 27845 -1177
rect 27572 -1331 27573 -1304
rect 27573 -1331 27606 -1304
rect 27652 -1331 27653 -1304
rect 27653 -1331 27686 -1304
rect 27732 -1331 27733 -1304
rect 27733 -1331 27766 -1304
rect 27811 -1331 27813 -1304
rect 27813 -1331 27845 -1304
rect 27572 -1338 27606 -1331
rect 27652 -1338 27686 -1331
rect 27732 -1338 27766 -1331
rect 27811 -1338 27845 -1331
rect 27578 -1716 27607 -1685
rect 27607 -1716 27612 -1685
rect 27578 -1719 27612 -1716
rect 27653 -1716 27687 -1685
rect 27653 -1719 27687 -1716
rect 27728 -1716 27733 -1685
rect 27733 -1716 27762 -1685
rect 27803 -1716 27813 -1685
rect 27813 -1716 27837 -1685
rect 27728 -1719 27762 -1716
rect 27803 -1719 27837 -1716
rect 30280 -1924 30314 -1890
rect 30280 -1998 30314 -1964
rect 30280 -2073 30314 -2039
rect 30280 -2148 30314 -2114
rect 30042 -2226 30076 -2192
rect 30124 -2226 30158 -2192
rect 30206 -2226 30240 -2192
rect 30288 -2226 30322 -2192
rect 30042 -2301 30076 -2267
rect 30124 -2301 30158 -2267
rect 30206 -2301 30240 -2267
rect 30288 -2301 30322 -2267
rect 30042 -2376 30076 -2342
rect 30124 -2376 30158 -2342
rect 30206 -2376 30240 -2342
rect 30288 -2376 30322 -2342
rect 30042 -2451 30076 -2417
rect 30124 -2451 30158 -2417
rect 30206 -2451 30240 -2417
rect 30288 -2451 30322 -2417
rect 30042 -2527 30076 -2493
rect 30124 -2527 30158 -2493
rect 30206 -2527 30240 -2493
rect 30288 -2527 30322 -2493
rect 30042 -2603 30076 -2569
rect 30124 -2603 30158 -2569
rect 30206 -2603 30240 -2569
rect 30288 -2603 30322 -2569
rect 30042 -2679 30076 -2645
rect 30124 -2679 30158 -2645
rect 30206 -2679 30240 -2645
rect 30288 -2679 30322 -2645
rect 30042 -2755 30076 -2721
rect 30124 -2755 30158 -2721
rect 30206 -2755 30240 -2721
rect 30288 -2755 30322 -2721
rect 30042 -2831 30076 -2797
rect 30124 -2831 30158 -2797
rect 30206 -2831 30240 -2797
rect 30288 -2831 30322 -2797
rect 30042 -2907 30076 -2873
rect 30124 -2907 30158 -2873
rect 30206 -2907 30240 -2873
rect 30288 -2907 30322 -2873
rect 28098 -2948 28132 -2945
rect 28098 -2979 28122 -2948
rect 28122 -2979 28132 -2948
rect 28218 -2979 28252 -2945
rect 30042 -2983 30076 -2949
rect 30124 -2983 30158 -2949
rect 30206 -2983 30240 -2949
rect 30288 -2983 30322 -2949
rect 28098 -3051 28122 -3022
rect 28122 -3051 28132 -3022
rect 28098 -3056 28132 -3051
rect 28218 -3056 28252 -3022
rect 28098 -3120 28122 -3099
rect 28122 -3120 28132 -3099
rect 28098 -3133 28132 -3120
rect 28218 -3133 28252 -3099
rect 28098 -3189 28122 -3176
rect 28122 -3189 28132 -3176
rect 28098 -3210 28132 -3189
rect 28218 -3210 28252 -3176
rect 28098 -3258 28122 -3254
rect 28122 -3258 28132 -3254
rect 28098 -3288 28132 -3258
rect 28218 -3288 28252 -3254
rect 28098 -3362 28132 -3332
rect 28098 -3366 28122 -3362
rect 28122 -3366 28132 -3362
rect 28218 -3366 28252 -3332
rect 28098 -3432 28132 -3410
rect 28098 -3444 28122 -3432
rect 28122 -3444 28132 -3432
rect 28218 -3444 28252 -3410
rect 34118 -3871 34152 -3837
rect 34118 -3943 34152 -3909
<< metal1 >>
rect 25969 1718 26131 1730
rect 25969 1684 25981 1718
rect 26015 1684 26131 1718
rect 25969 1646 26131 1684
rect 25969 1612 25981 1646
rect 26015 1612 26131 1646
rect 25969 1574 26131 1612
rect 26296 1600 26324 1628
rect 25969 1540 25981 1574
rect 26015 1540 26131 1574
rect 25969 1502 26131 1540
rect 25969 1468 25981 1502
rect 26015 1468 26131 1502
rect 25969 1430 26131 1468
rect 25969 1396 25981 1430
rect 26015 1396 26131 1430
rect 25969 1384 26131 1396
rect 26743 885 26771 913
rect 26499 327 26551 333
rect 26499 263 26551 275
rect 26499 205 26551 211
rect 26872 327 26924 333
rect 26872 263 26924 275
tri 26924 234 27014 324 sw
rect 26924 211 27014 234
rect 26872 205 27014 211
tri 27014 205 27043 234 sw
tri 26964 155 27014 205 ne
rect 27014 155 27043 205
tri 27043 155 27093 205 sw
tri 27014 103 27066 155 ne
rect 27066 133 27849 155
tri 27849 133 27871 155 sw
rect 27066 103 27871 133
tri 27871 103 27901 133 sw
tri 27827 59 27871 103 ne
rect 27871 81 27901 103
tri 27901 81 27923 103 sw
rect 27871 33 27923 81
rect 27871 -31 27923 -19
rect 27871 -89 27923 -83
rect 26856 -555 28669 -547
tri 28669 -555 28677 -547 sw
rect 26856 -579 28677 -555
tri 28677 -579 28701 -555 sw
tri 28655 -601 28677 -579 ne
rect 28677 -601 28701 -579
tri 28701 -601 28723 -579 sw
tri 28677 -615 28691 -601 ne
rect 26218 -721 26270 -715
rect 26218 -787 26270 -773
rect 28205 -769 28257 -763
rect 26514 -819 26542 -791
rect 26218 -845 26270 -839
rect 26660 -842 26666 -790
rect 26718 -842 26746 -790
rect 26798 -842 26825 -790
rect 26877 -842 26883 -790
rect 26660 -868 26883 -842
rect 28363 -819 28391 -791
rect 28205 -833 28257 -821
tri 27981 -850 27984 -847 se
rect 27984 -850 27990 -847
rect 26660 -920 26666 -868
rect 26718 -920 26746 -868
rect 26798 -920 26825 -868
rect 26877 -920 26883 -868
rect 27327 -856 27990 -850
rect 28042 -856 28054 -847
rect 27327 -890 27339 -856
rect 27373 -890 27414 -856
rect 27448 -890 27489 -856
rect 27523 -890 27564 -856
rect 27598 -890 27639 -856
rect 27673 -890 27714 -856
rect 27748 -890 27789 -856
rect 27823 -890 27864 -856
rect 27898 -890 27939 -856
rect 27973 -890 27990 -856
rect 28047 -890 28054 -856
rect 27327 -896 27990 -890
tri 27981 -899 27984 -896 ne
rect 27984 -899 27990 -896
rect 28042 -899 28054 -890
rect 28106 -899 28112 -847
rect 28205 -891 28257 -885
rect 28691 -1037 28723 -601
rect 28784 -699 29140 -692
rect 28784 -714 28796 -699
rect 28830 -714 28871 -699
rect 28905 -714 28946 -699
rect 28784 -766 28786 -714
rect 28838 -733 28871 -714
rect 28938 -733 28946 -714
rect 28980 -714 29020 -699
rect 29054 -714 29094 -699
rect 29128 -714 29140 -699
rect 28980 -733 28986 -714
rect 29054 -733 29086 -714
rect 28838 -766 28886 -733
rect 28938 -766 28986 -733
rect 29038 -766 29086 -733
rect 29138 -766 29140 -714
rect 28784 -778 29140 -766
rect 28784 -830 28786 -778
rect 28838 -783 28886 -778
rect 28938 -783 28986 -778
rect 29038 -783 29086 -778
rect 28838 -817 28871 -783
rect 28938 -817 28946 -783
rect 28980 -817 28986 -783
rect 29054 -817 29086 -783
rect 28838 -830 28886 -817
rect 28938 -830 28986 -817
rect 29038 -830 29086 -817
rect 29138 -830 29140 -778
rect 28784 -867 29140 -830
rect 28784 -901 28796 -867
rect 28830 -901 28871 -867
rect 28905 -901 28946 -867
rect 28980 -901 29020 -867
rect 29054 -901 29094 -867
rect 29128 -901 29140 -867
rect 28784 -951 29140 -901
rect 29756 -923 29762 -871
rect 29814 -923 29826 -871
rect 29878 -923 29884 -871
rect 30241 -892 30771 -864
rect 28784 -985 28796 -951
rect 28830 -985 28871 -951
rect 28905 -985 28946 -951
rect 28980 -985 29020 -951
rect 29054 -985 29094 -951
rect 29128 -985 29140 -951
rect 28784 -992 29140 -985
tri 28691 -1057 28711 -1037 ne
rect 28711 -1057 28723 -1037
tri 28723 -1057 28757 -1023 sw
tri 28711 -1062 28716 -1057 ne
rect 28716 -1062 29018 -1057
rect 27142 -1090 27170 -1062
tri 28716 -1065 28719 -1062 ne
rect 28719 -1065 29018 -1062
rect 27432 -1093 27460 -1065
tri 28719 -1069 28723 -1065 ne
rect 28723 -1069 29018 -1065
tri 28723 -1093 28747 -1069 ne
rect 28747 -1093 29018 -1069
tri 28747 -1103 28757 -1093 ne
rect 28757 -1103 29018 -1093
rect 29758 -1065 29810 -923
rect 29758 -1129 29810 -1117
rect 27560 -1164 27857 -1158
rect 27560 -1198 27572 -1164
rect 27606 -1198 27652 -1164
rect 27686 -1198 27731 -1164
rect 27560 -1216 27731 -1198
rect 27783 -1216 27805 -1164
rect 29758 -1187 29810 -1181
rect 27560 -1286 27857 -1216
rect 27560 -1304 27731 -1286
rect 27560 -1338 27572 -1304
rect 27606 -1338 27652 -1304
rect 27686 -1338 27731 -1304
rect 27783 -1338 27805 -1286
rect 27560 -1344 27857 -1338
rect 28145 -1465 28151 -1413
rect 28203 -1465 28215 -1413
rect 28267 -1465 28273 -1413
rect 27436 -1685 28196 -1661
rect 27436 -1719 27578 -1685
rect 27612 -1719 27653 -1685
rect 27687 -1719 27728 -1685
rect 27762 -1719 27803 -1685
rect 27837 -1719 28196 -1685
rect 27436 -1858 28196 -1719
rect 28787 -1747 28815 -1719
tri 30203 -1890 30235 -1858 ne
rect 30235 -1890 30328 -1858
tri 30235 -1921 30266 -1890 ne
rect 30266 -1924 30280 -1890
rect 30314 -1924 30328 -1890
tri 30328 -1921 30391 -1858 nw
rect 30266 -1964 30328 -1924
rect 30266 -1998 30280 -1964
rect 30314 -1998 30328 -1964
rect 30266 -2039 30328 -1998
rect 30266 -2073 30280 -2039
rect 30314 -2073 30328 -2039
tri 30239 -2114 30266 -2087 se
rect 30266 -2114 30328 -2073
tri 30205 -2148 30239 -2114 se
rect 30239 -2148 30280 -2114
rect 30314 -2148 30328 -2114
rect 31155 -2024 31207 -2018
rect 31155 -2088 31207 -2076
tri 30173 -2180 30205 -2148 se
rect 30205 -2180 30328 -2148
rect 30036 -2192 30328 -2180
rect 30698 -2189 30704 -2137
rect 30756 -2189 30768 -2137
rect 30820 -2189 30826 -2137
tri 36776 -2118 36784 -2110 se
rect 36784 -2118 36790 -2110
rect 31207 -2140 36790 -2118
rect 31155 -2146 36790 -2140
tri 36768 -2162 36784 -2146 ne
rect 36784 -2162 36790 -2146
rect 36842 -2162 36854 -2110
rect 36906 -2162 36912 -2110
rect 30036 -2226 30042 -2192
rect 30076 -2226 30124 -2192
rect 30158 -2226 30206 -2192
rect 30240 -2226 30288 -2192
rect 30322 -2226 30328 -2192
tri 30734 -2226 30771 -2189 ne
rect 30771 -2226 30826 -2189
rect 30036 -2267 30328 -2226
tri 30771 -2253 30798 -2226 ne
rect 30036 -2301 30042 -2267
rect 30076 -2301 30124 -2267
rect 30158 -2301 30206 -2267
rect 30240 -2301 30288 -2267
rect 30322 -2301 30328 -2267
rect 30036 -2342 30328 -2301
rect 30036 -2376 30042 -2342
rect 30076 -2376 30124 -2342
rect 30158 -2376 30206 -2342
rect 30240 -2376 30288 -2342
rect 30322 -2376 30328 -2342
rect 30036 -2417 30328 -2376
rect 30036 -2451 30042 -2417
rect 30076 -2451 30124 -2417
rect 30158 -2451 30206 -2417
rect 30240 -2451 30288 -2417
rect 30322 -2451 30328 -2417
rect 28020 -2548 28048 -2520
rect 29406 -2554 29412 -2502
rect 29464 -2554 29476 -2502
rect 29528 -2554 29534 -2502
rect 29637 -2530 29643 -2478
rect 29695 -2530 29709 -2478
rect 29761 -2530 29767 -2478
rect 30036 -2493 30328 -2451
rect 30036 -2527 30042 -2493
rect 30076 -2527 30124 -2493
rect 30158 -2527 30206 -2493
rect 30240 -2527 30288 -2493
rect 30322 -2527 30328 -2493
rect 30036 -2569 30328 -2527
rect 30036 -2603 30042 -2569
rect 30076 -2603 30124 -2569
rect 30158 -2603 30206 -2569
rect 30240 -2603 30288 -2569
rect 30322 -2603 30328 -2569
rect 30036 -2645 30328 -2603
tri 30020 -2679 30036 -2663 se
rect 30036 -2679 30042 -2645
rect 30076 -2679 30124 -2645
rect 30158 -2679 30206 -2645
rect 30240 -2679 30288 -2645
rect 30322 -2679 30328 -2645
tri 29988 -2711 30020 -2679 se
rect 30020 -2711 30328 -2679
rect 29916 -2721 30328 -2711
rect 29916 -2755 30042 -2721
rect 30076 -2755 30124 -2721
rect 30158 -2755 30206 -2721
rect 30240 -2755 30288 -2721
rect 30322 -2755 30328 -2721
rect 29916 -2797 30328 -2755
rect 29916 -2831 30042 -2797
rect 30076 -2831 30124 -2797
rect 30158 -2831 30206 -2797
rect 30240 -2831 30288 -2797
rect 30322 -2831 30328 -2797
rect 29916 -2873 30328 -2831
rect 29916 -2907 30042 -2873
rect 30076 -2907 30124 -2873
rect 30158 -2907 30206 -2873
rect 30240 -2907 30288 -2873
rect 30322 -2907 30328 -2873
rect 29916 -2925 30328 -2907
tri 29966 -2933 29974 -2925 ne
rect 29974 -2933 30328 -2925
rect 28092 -2945 28258 -2933
rect 28092 -2979 28098 -2945
rect 28132 -2979 28218 -2945
rect 28252 -2979 28258 -2945
tri 29974 -2949 29990 -2933 ne
rect 29990 -2949 30328 -2933
rect 28092 -3022 28258 -2979
tri 29990 -2983 30024 -2949 ne
rect 30024 -2983 30042 -2949
rect 30076 -2983 30124 -2949
rect 30158 -2983 30206 -2949
rect 30240 -2983 30288 -2949
rect 30322 -2983 30328 -2949
tri 30024 -2995 30036 -2983 ne
rect 30036 -2995 30328 -2983
rect 28092 -3056 28098 -3022
rect 28132 -3056 28218 -3022
rect 28252 -3056 28258 -3022
rect 28092 -3099 28258 -3056
rect 28092 -3133 28098 -3099
rect 28132 -3133 28218 -3099
rect 28252 -3133 28258 -3099
rect 28092 -3176 28258 -3133
tri 30079 -3136 30105 -3110 se
rect 30105 -3136 30491 -3110
tri 30073 -3142 30079 -3136 se
rect 30079 -3142 30491 -3136
rect 28637 -3170 28665 -3142
tri 30061 -3154 30073 -3142 se
rect 30073 -3154 30439 -3142
rect 28092 -3210 28098 -3176
rect 28132 -3210 28218 -3176
rect 28252 -3210 28258 -3176
rect 28787 -3182 28815 -3154
tri 30033 -3182 30061 -3154 se
rect 30061 -3162 30439 -3154
rect 30061 -3182 30105 -3162
tri 30031 -3184 30033 -3182 se
rect 30033 -3184 30105 -3182
tri 30105 -3184 30127 -3162 nw
rect 28092 -3254 28258 -3210
tri 29977 -3238 30031 -3184 se
rect 30031 -3238 30051 -3184
tri 30051 -3238 30105 -3184 nw
rect 30439 -3206 30491 -3194
rect 28092 -3288 28098 -3254
rect 28132 -3288 28218 -3254
rect 28252 -3288 28258 -3254
rect 29689 -3264 30025 -3238
tri 30025 -3264 30051 -3238 nw
rect 30439 -3264 30491 -3258
rect 29689 -3266 30023 -3264
tri 30023 -3266 30025 -3264 nw
rect 28092 -3332 28258 -3288
rect 28092 -3366 28098 -3332
rect 28132 -3366 28218 -3332
rect 28252 -3366 28258 -3332
rect 28092 -3410 28258 -3366
rect 28092 -3444 28098 -3410
rect 28132 -3444 28218 -3410
rect 28252 -3444 28258 -3410
rect 28092 -3456 28258 -3444
rect 30285 -3334 30337 -3328
rect 30285 -3400 30337 -3386
rect 30285 -3458 30337 -3452
rect 30377 -3371 30429 -3365
rect 30377 -3435 30429 -3423
rect 28983 -3582 29011 -3554
rect 30186 -3585 30232 -3542
rect 30377 -3585 30429 -3487
rect 30186 -3631 30429 -3585
rect 27192 -3710 27244 -3704
rect 27192 -3779 27244 -3762
rect 27326 -3826 27354 -3798
rect 27192 -3848 27244 -3831
rect 27192 -3906 27244 -3900
rect 27929 -3955 28909 -3934
rect 27929 -4007 28685 -3955
rect 28737 -4007 28768 -3955
rect 28820 -4007 28851 -3955
rect 28903 -4007 28909 -3955
rect 26087 -4027 26344 -4021
rect 26139 -4079 26292 -4027
rect 27929 -4028 28909 -4007
rect 26087 -4091 26344 -4079
rect 28136 -4088 28164 -4060
rect 26139 -4143 26292 -4091
rect 26087 -4149 26344 -4143
rect 26328 -4190 26380 -4184
rect 28361 -4216 28389 -4188
rect 26328 -4256 26380 -4242
rect 26328 -4314 26380 -4308
rect 27288 -4277 27340 -4271
tri 27254 -4371 27288 -4337 se
rect 27288 -4341 27340 -4329
tri 26936 -4399 26964 -4371 se
rect 26964 -4393 27288 -4371
rect 26964 -4399 27340 -4393
tri 26925 -4410 26936 -4399 se
rect 26936 -4410 26977 -4399
tri 26977 -4410 26988 -4399 nw
rect 26702 -4418 26969 -4410
tri 26969 -4418 26977 -4410 nw
rect 26702 -4451 26936 -4418
tri 26936 -4451 26969 -4418 nw
rect 26702 -4470 26717 -4451
tri 26717 -4470 26736 -4451 nw
rect 26702 -4477 26710 -4470
tri 26710 -4477 26717 -4470 nw
rect 26702 -4482 26705 -4477
tri 26705 -4482 26710 -4477 nw
tri 26702 -4485 26705 -4482 nw
rect 27319 -4493 27347 -4465
rect 28153 -4516 28205 -4510
rect 28153 -4580 28205 -4568
rect 28679 -4534 28685 -4482
rect 28737 -4534 28778 -4482
rect 28830 -4534 28870 -4482
rect 28922 -4534 28928 -4482
rect 28679 -4560 28928 -4534
rect 28938 -4558 28966 -4530
rect 28679 -4612 28685 -4560
rect 28737 -4612 28778 -4560
rect 28830 -4612 28870 -4560
rect 28922 -4612 28928 -4560
rect 28153 -4638 28205 -4632
rect 26773 -4692 26801 -4664
rect 27662 -4806 27668 -4754
rect 27720 -4806 27732 -4754
rect 27784 -4806 27790 -4754
rect 29152 -4932 29180 -4904
tri 27162 -5083 27192 -5053 se
rect 27192 -5059 27244 -5053
tri 27244 -5083 27274 -5053 sw
rect 27192 -5123 27244 -5111
rect 26442 -5168 26470 -5140
rect 27192 -5181 27244 -5175
rect 29480 -5263 29486 -5211
rect 29538 -5263 29550 -5211
rect 29602 -5263 29608 -5211
rect 26822 -5464 26874 -5458
rect 26110 -5521 26162 -5515
tri 26788 -5558 26822 -5524 se
rect 26822 -5528 26874 -5516
rect 26110 -5585 26162 -5573
tri 26874 -5549 26965 -5458 nw
rect 30798 -5511 30826 -2226
rect 31155 -2190 31207 -2184
rect 31881 -2226 31887 -2174
rect 31939 -2226 31951 -2174
rect 32003 -2226 32009 -2174
rect 31155 -2254 31207 -2242
tri 32128 -2255 32146 -2237 se
rect 32146 -2250 32975 -2237
tri 32975 -2250 32988 -2237 sw
rect 32146 -2255 32988 -2250
rect 31207 -2256 32988 -2255
tri 32988 -2256 32994 -2250 sw
tri 33972 -2256 33978 -2250 se
rect 33978 -2256 33984 -2250
rect 31207 -2265 33984 -2256
rect 31207 -2283 32174 -2265
tri 32174 -2283 32192 -2265 nw
tri 32910 -2283 32928 -2265 ne
rect 32928 -2283 33984 -2265
tri 32928 -2293 32938 -2283 ne
rect 32938 -2293 33984 -2283
tri 32552 -2300 32559 -2293 se
rect 32559 -2300 32852 -2293
rect 31155 -2312 31207 -2306
rect 31155 -2348 31207 -2342
rect 32232 -2352 32238 -2300
rect 32290 -2352 32302 -2300
rect 32354 -2311 32360 -2300
tri 32360 -2311 32371 -2300 sw
tri 32541 -2311 32552 -2300 se
rect 32552 -2311 32852 -2300
rect 32354 -2321 32852 -2311
rect 32354 -2330 32596 -2321
tri 32596 -2330 32605 -2321 nw
tri 32787 -2330 32796 -2321 ne
rect 32796 -2330 32852 -2321
tri 32852 -2330 32889 -2293 sw
tri 32938 -2302 32947 -2293 ne
rect 32947 -2302 33984 -2293
rect 34036 -2302 34048 -2250
rect 34100 -2302 34106 -2250
rect 32354 -2331 32595 -2330
tri 32595 -2331 32596 -2330 nw
tri 32796 -2331 32797 -2330 ne
rect 32797 -2331 35722 -2330
tri 35722 -2331 35723 -2330 sw
rect 32354 -2339 32587 -2331
tri 32587 -2339 32595 -2331 nw
tri 32797 -2339 32805 -2331 ne
rect 32805 -2339 36437 -2331
rect 32354 -2342 32370 -2339
tri 32370 -2342 32373 -2339 nw
tri 32805 -2342 32808 -2339 ne
rect 32808 -2342 36437 -2339
rect 32354 -2349 32363 -2342
tri 32363 -2349 32370 -2342 nw
tri 32808 -2349 32815 -2342 ne
rect 32815 -2349 36437 -2342
rect 32354 -2352 32360 -2349
tri 32360 -2352 32363 -2349 nw
tri 32815 -2352 32818 -2349 ne
rect 32818 -2352 36437 -2349
tri 32818 -2358 32824 -2352 ne
rect 32824 -2358 36437 -2352
tri 35693 -2359 35694 -2358 ne
rect 35694 -2359 36437 -2358
tri 36407 -2383 36431 -2359 ne
rect 36431 -2383 36437 -2359
rect 36489 -2383 36501 -2331
rect 36553 -2383 36559 -2331
rect 31155 -2412 31207 -2400
rect 36703 -2411 36731 -2383
tri 31207 -2442 31233 -2416 sw
rect 31207 -2464 34581 -2442
rect 31155 -2470 34581 -2464
rect 34575 -2494 34581 -2470
rect 34633 -2494 34645 -2442
rect 34697 -2494 34703 -2442
rect 31174 -2542 34340 -2498
rect 31174 -2550 31696 -2542
tri 31696 -2550 31704 -2542 nw
tri 34326 -2550 34334 -2542 ne
rect 34334 -2550 34340 -2542
rect 34392 -2550 34404 -2498
rect 34456 -2550 34462 -2498
rect 31174 -2580 31226 -2550
tri 31937 -2595 31961 -2571 se
rect 31961 -2595 31976 -2571
rect 31174 -2644 31226 -2632
rect 31174 -2702 31226 -2696
rect 31393 -2601 31976 -2595
rect 31445 -2604 31976 -2601
rect 31445 -2623 31961 -2604
rect 31393 -2665 31445 -2653
rect 31393 -2723 31445 -2717
rect 35376 -2739 35404 -2711
rect 32811 -2844 32825 -2792
rect 32877 -2844 32889 -2792
rect 32941 -2844 33853 -2792
rect 33905 -2844 33917 -2792
rect 33969 -2844 33975 -2792
rect 37380 -2821 37408 -2793
rect 32208 -3047 32236 -3019
rect 35760 -3047 35788 -3019
rect 32772 -3116 32824 -3110
rect 31174 -3184 31226 -3178
tri 31226 -3212 31260 -3178 sw
rect 32772 -3180 32824 -3168
rect 31226 -3232 32772 -3212
rect 31226 -3236 32824 -3232
rect 31174 -3248 32824 -3236
rect 31226 -3264 32824 -3248
tri 31226 -3298 31260 -3264 nw
rect 31174 -3306 31226 -3300
rect 35376 -3355 35404 -3327
rect 31174 -3365 31226 -3359
rect 31174 -3429 31226 -3417
tri 31226 -3458 31259 -3425 sw
tri 31682 -3458 31715 -3425 se
rect 31226 -3459 31259 -3458
tri 31259 -3459 31260 -3458 sw
tri 31681 -3459 31682 -3458 se
rect 31682 -3459 31715 -3458
tri 31767 -3458 31800 -3425 sw
tri 33001 -3458 33016 -3443 se
rect 33016 -3458 33022 -3443
rect 31767 -3459 31800 -3458
tri 31800 -3459 31801 -3458 sw
tri 33000 -3459 33001 -3458 se
rect 33001 -3459 33022 -3458
rect 31226 -3481 33022 -3459
rect 31174 -3487 33022 -3481
tri 33008 -3495 33016 -3487 ne
rect 33016 -3495 33022 -3487
rect 33074 -3495 33086 -3443
rect 33138 -3495 33144 -3443
rect 34495 -3573 34548 -3567
tri 31011 -3589 31022 -3578 se
tri 31050 -3589 31061 -3578 sw
rect 31009 -3595 31061 -3589
rect 31009 -3659 31061 -3647
rect 31009 -3717 31061 -3711
rect 31175 -3595 31963 -3589
rect 31227 -3617 31911 -3595
tri 31883 -3645 31911 -3617 ne
rect 31175 -3659 31227 -3647
rect 31175 -3717 31227 -3711
rect 34387 -3605 34439 -3599
rect 31911 -3659 31963 -3647
tri 34353 -3681 34387 -3647 se
rect 34387 -3669 34439 -3657
tri 31011 -3728 31022 -3717 ne
tri 31050 -3728 31061 -3717 nw
rect 31325 -3718 31377 -3712
rect 31911 -3717 31963 -3711
rect 33752 -3713 33780 -3685
rect 34547 -3579 34548 -3573
rect 34495 -3637 34547 -3625
tri 34439 -3681 34445 -3675 sw
rect 34495 -3709 34547 -3689
rect 34387 -3727 34439 -3721
tri 35009 -3727 35014 -3722 sw
rect 35009 -3730 35014 -3727
tri 35014 -3730 35017 -3727 sw
rect 35760 -3734 35788 -3706
rect 35009 -3764 35013 -3758
tri 35013 -3764 35019 -3758 nw
tri 35009 -3768 35013 -3764 nw
rect 31325 -3782 31377 -3770
rect 31174 -3837 31226 -3831
tri 31377 -3812 31411 -3778 sw
rect 31377 -3816 32408 -3812
tri 32408 -3816 32412 -3812 sw
rect 35878 -3816 35884 -3764
rect 35936 -3816 35948 -3764
rect 36000 -3816 36006 -3764
rect 31377 -3834 32412 -3816
rect 31325 -3837 32412 -3834
tri 32412 -3837 32433 -3816 sw
rect 34112 -3837 34158 -3825
rect 31325 -3840 32433 -3837
tri 32433 -3840 32436 -3837 sw
tri 32382 -3865 32407 -3840 ne
rect 32407 -3865 32436 -3840
tri 32436 -3865 32461 -3840 sw
tri 32407 -3866 32408 -3865 ne
rect 32408 -3866 32461 -3865
tri 32408 -3871 32413 -3866 ne
rect 32413 -3871 32461 -3866
tri 32461 -3871 32467 -3865 sw
rect 34112 -3871 34118 -3837
rect 34152 -3840 34158 -3837
tri 34158 -3840 34173 -3825 sw
rect 34152 -3853 34173 -3840
tri 34173 -3853 34186 -3840 sw
rect 34152 -3856 34482 -3853
rect 34152 -3871 34357 -3856
tri 32413 -3878 32420 -3871 ne
rect 32420 -3878 32467 -3871
tri 31226 -3888 31236 -3878 sw
tri 32420 -3888 32430 -3878 ne
rect 32430 -3888 32467 -3878
rect 31226 -3889 31236 -3888
rect 31174 -3901 31236 -3889
rect 31226 -3909 31236 -3901
tri 31236 -3909 31257 -3888 sw
tri 31774 -3909 31795 -3888 se
rect 31795 -3909 31801 -3888
rect 31226 -3912 31257 -3909
tri 31257 -3912 31260 -3909 sw
tri 31771 -3912 31774 -3909 se
rect 31774 -3912 31801 -3909
rect 31226 -3940 31801 -3912
rect 31853 -3940 31865 -3888
rect 31917 -3940 31923 -3888
tri 32430 -3909 32451 -3888 ne
rect 32451 -3903 32467 -3888
tri 32467 -3903 32499 -3871 sw
rect 32451 -3909 32499 -3903
tri 32499 -3909 32505 -3903 sw
tri 32753 -3909 32759 -3903 se
rect 32759 -3909 32765 -3903
tri 32451 -3919 32461 -3909 ne
rect 32461 -3919 32505 -3909
tri 32505 -3919 32515 -3909 sw
tri 32743 -3919 32753 -3909 se
rect 32753 -3919 32765 -3909
tri 32461 -3940 32482 -3919 ne
rect 32482 -3940 32765 -3919
rect 31226 -3943 31242 -3940
tri 31242 -3943 31245 -3940 nw
tri 32482 -3943 32485 -3940 ne
rect 32485 -3943 32765 -3940
rect 31226 -3947 31238 -3943
tri 31238 -3947 31242 -3943 nw
tri 32485 -3947 32489 -3943 ne
rect 32489 -3947 32765 -3943
rect 31226 -3953 31230 -3947
rect 31174 -3955 31230 -3953
tri 31230 -3955 31238 -3947 nw
tri 32751 -3955 32759 -3947 ne
rect 32759 -3955 32765 -3947
rect 32817 -3955 32829 -3903
rect 32881 -3955 32887 -3903
rect 34112 -3908 34357 -3871
rect 34409 -3908 34421 -3856
rect 34473 -3908 34482 -3856
rect 34112 -3909 34482 -3908
rect 34112 -3943 34118 -3909
rect 34152 -3910 34482 -3909
rect 34152 -3943 34158 -3910
rect 34112 -3955 34158 -3943
tri 34158 -3955 34203 -3910 nw
rect 31174 -3959 31226 -3955
tri 31226 -3959 31230 -3955 nw
rect 35376 -4018 35404 -3990
rect 37007 -4065 37035 -4037
tri 31126 -4088 31136 -4078 sw
rect 31126 -4112 31136 -4088
tri 31136 -4112 31160 -4088 sw
rect 35878 -4112 35884 -4088
rect 31126 -4140 35884 -4112
rect 35936 -4140 35948 -4088
rect 36000 -4140 36006 -4088
rect 31126 -4149 31151 -4140
tri 31151 -4149 31160 -4140 nw
tri 31126 -4174 31151 -4149 nw
rect 32768 -4293 32796 -4265
rect 35238 -4290 35266 -4262
tri 31532 -4418 31566 -4384 sw
rect 32724 -4470 32730 -4418
rect 32782 -4470 32794 -4418
rect 32846 -4446 34503 -4418
tri 34503 -4446 34531 -4418 sw
rect 32846 -4470 32852 -4446
tri 34457 -4470 34481 -4446 ne
rect 34481 -4467 34531 -4446
tri 34531 -4467 34552 -4446 sw
rect 34481 -4470 34559 -4467
tri 31532 -4477 31539 -4470 nw
tri 34481 -4474 34485 -4470 ne
rect 34485 -4474 34559 -4470
tri 33341 -4477 33344 -4474 se
rect 33344 -4477 34042 -4474
tri 34485 -4477 34488 -4474 ne
rect 34488 -4477 34559 -4474
tri 33310 -4508 33341 -4477 se
rect 33341 -4502 34042 -4477
rect 33341 -4508 33400 -4502
tri 33400 -4508 33406 -4502 nw
rect 32626 -4520 33388 -4508
tri 33388 -4520 33400 -4508 nw
rect 32626 -4536 33372 -4520
tri 33372 -4536 33388 -4520 nw
rect 32928 -4592 33726 -4564
rect 32928 -4691 32974 -4592
rect 34014 -4614 34042 -4502
tri 34488 -4520 34531 -4477 ne
rect 34531 -4520 34559 -4477
tri 34531 -4548 34559 -4520 ne
rect 34311 -4621 34317 -4569
rect 34369 -4621 34381 -4569
rect 34433 -4621 34439 -4569
rect 34567 -4571 34595 -4543
rect 35057 -4585 35109 -4579
rect 33618 -4634 33670 -4628
rect 33086 -4668 33114 -4640
rect 33370 -4682 33618 -4636
rect 32308 -4796 32360 -4790
rect 33370 -4804 33416 -4682
rect 34402 -4670 34430 -4642
rect 35057 -4648 35109 -4637
rect 35044 -4649 35109 -4648
rect 35044 -4676 35057 -4649
rect 33618 -4698 33670 -4686
tri 35109 -4662 35147 -4624 nw
rect 35057 -4707 35109 -4701
rect 33618 -4756 33670 -4750
rect 32308 -4860 32360 -4848
rect 32531 -4885 32559 -4857
rect 34776 -4866 34782 -4814
rect 34834 -4866 34846 -4814
rect 34898 -4866 34904 -4814
rect 34851 -4893 34879 -4866
rect 35246 -4908 35252 -4856
rect 35304 -4908 35316 -4856
rect 35368 -4908 35374 -4856
rect 35982 -4872 36010 -4859
rect 32308 -4918 32360 -4912
rect 35964 -4924 35970 -4872
rect 36022 -4924 36034 -4872
rect 36086 -4924 36092 -4872
rect 32823 -5096 32851 -5068
rect 35269 -5113 35297 -5085
rect 32991 -5280 33043 -5274
tri 32953 -5350 32991 -5312 se
rect 38006 -5292 38235 -5264
rect 32991 -5344 33043 -5332
rect 32244 -5402 32250 -5350
rect 32302 -5402 32314 -5350
rect 32366 -5396 32991 -5350
rect 32366 -5402 33043 -5396
rect 38125 -5336 38157 -5320
tri 38157 -5336 38173 -5320 sw
rect 36626 -5468 36654 -5440
rect 30774 -5517 30826 -5511
rect 26822 -5586 26874 -5580
rect 30774 -5581 30826 -5569
tri 26162 -5591 26167 -5586 sw
rect 26162 -5615 26167 -5591
tri 26167 -5615 26191 -5591 sw
rect 27681 -5615 27687 -5591
rect 26162 -5637 27687 -5615
rect 26110 -5643 27687 -5637
rect 27739 -5643 27751 -5591
rect 27803 -5643 27809 -5591
rect 30774 -5639 30826 -5633
rect 26599 -5823 26651 -5817
rect 26506 -5880 26558 -5874
rect 26386 -5946 26438 -5940
rect 26386 -6010 26438 -5998
rect 26506 -5944 26558 -5932
rect 27191 -5873 27197 -5821
rect 27249 -5873 27261 -5821
rect 27313 -5827 32351 -5821
rect 27313 -5849 32299 -5827
rect 27313 -5873 27319 -5849
rect 26599 -5887 26651 -5875
rect 32299 -5891 32351 -5879
rect 31143 -5917 31149 -5893
rect 26651 -5939 31149 -5917
rect 26599 -5945 31149 -5939
rect 31201 -5945 31213 -5893
rect 31265 -5945 31271 -5893
rect 32299 -5949 32351 -5943
rect 32416 -5829 32540 -5823
rect 32468 -5881 32488 -5829
rect 32416 -5895 32540 -5881
rect 32468 -5947 32488 -5895
rect 32863 -5897 32891 -5869
tri 38124 -5893 38125 -5892 se
rect 38125 -5893 38173 -5336
rect 38207 -5366 38235 -5292
tri 38121 -5896 38124 -5893 se
rect 38124 -5896 38173 -5893
rect 32416 -5953 32540 -5947
rect 38121 -5902 38173 -5896
rect 38121 -5966 38173 -5954
rect 26558 -5996 31311 -5973
rect 26506 -6001 31311 -5996
rect 26506 -6002 26558 -6001
rect 31305 -6025 31311 -6001
rect 31363 -6025 31375 -5973
rect 31427 -6025 31433 -5973
tri 33132 -6006 33157 -5981 se
rect 33157 -5987 33209 -5981
rect 30727 -6040 30733 -6029
rect 26438 -6062 30733 -6040
rect 26386 -6068 30733 -6062
rect 30727 -6081 30733 -6068
rect 30785 -6081 30797 -6029
rect 30849 -6081 30855 -6029
rect 32949 -6039 33157 -6006
rect 36491 -6038 36519 -6010
rect 38121 -6024 38173 -6018
rect 38207 -6019 38259 -5540
rect 32949 -6051 33209 -6039
rect 32949 -6052 33157 -6051
rect 32949 -6093 32995 -6052
tri 33126 -6083 33157 -6052 ne
rect 32633 -6099 32695 -6093
rect 32633 -6151 32643 -6099
rect 33157 -6109 33209 -6103
rect 38207 -6083 38259 -6071
rect 38207 -6141 38259 -6135
rect 32633 -6163 32695 -6151
rect 32633 -6215 32643 -6163
rect 32633 -6223 32695 -6215
rect 38044 -6278 38072 -6250
rect 27079 -6424 27107 -6396
rect 27621 -6954 27649 -6926
rect 26922 -7260 26950 -7232
rect 40211 -13346 40239 -13318
rect 41358 -13673 41386 -13645
rect 41427 -14232 41455 -14204
rect 40633 -14280 40661 -14252
rect 41023 -14572 41051 -14544
rect 40195 -14876 40223 -14848
rect 40244 -15218 40272 -15190
rect 40188 -15545 40216 -15517
<< via1 >>
rect 26499 275 26551 327
rect 26499 211 26551 263
rect 26872 275 26924 327
rect 26872 211 26924 263
rect 27871 -19 27923 33
rect 27871 -83 27923 -31
rect 26218 -773 26270 -721
rect 26218 -839 26270 -787
rect 26666 -842 26718 -790
rect 26746 -842 26798 -790
rect 26825 -842 26877 -790
rect 28205 -821 28257 -769
rect 26666 -920 26718 -868
rect 26746 -920 26798 -868
rect 26825 -920 26877 -868
rect 27990 -856 28042 -847
rect 27990 -890 28013 -856
rect 28013 -890 28042 -856
rect 27990 -899 28042 -890
rect 28054 -899 28106 -847
rect 28205 -885 28257 -833
rect 28786 -733 28796 -714
rect 28796 -733 28830 -714
rect 28830 -733 28838 -714
rect 28886 -733 28905 -714
rect 28905 -733 28938 -714
rect 28986 -733 29020 -714
rect 29020 -733 29038 -714
rect 29086 -733 29094 -714
rect 29094 -733 29128 -714
rect 29128 -733 29138 -714
rect 28786 -766 28838 -733
rect 28886 -766 28938 -733
rect 28986 -766 29038 -733
rect 29086 -766 29138 -733
rect 28786 -783 28838 -778
rect 28886 -783 28938 -778
rect 28986 -783 29038 -778
rect 29086 -783 29138 -778
rect 28786 -817 28796 -783
rect 28796 -817 28830 -783
rect 28830 -817 28838 -783
rect 28886 -817 28905 -783
rect 28905 -817 28938 -783
rect 28986 -817 29020 -783
rect 29020 -817 29038 -783
rect 29086 -817 29094 -783
rect 29094 -817 29128 -783
rect 29128 -817 29138 -783
rect 28786 -830 28838 -817
rect 28886 -830 28938 -817
rect 28986 -830 29038 -817
rect 29086 -830 29138 -817
rect 29762 -923 29814 -871
rect 29826 -923 29878 -871
rect 29758 -1117 29810 -1065
rect 27731 -1198 27732 -1164
rect 27732 -1198 27766 -1164
rect 27766 -1198 27783 -1164
rect 27731 -1216 27783 -1198
rect 27805 -1198 27811 -1164
rect 27811 -1198 27845 -1164
rect 27845 -1198 27857 -1164
rect 29758 -1181 29810 -1129
rect 27805 -1216 27857 -1198
rect 27731 -1304 27783 -1286
rect 27731 -1338 27732 -1304
rect 27732 -1338 27766 -1304
rect 27766 -1338 27783 -1304
rect 27805 -1304 27857 -1286
rect 27805 -1338 27811 -1304
rect 27811 -1338 27845 -1304
rect 27845 -1338 27857 -1304
rect 28151 -1465 28203 -1413
rect 28215 -1465 28267 -1413
rect 31155 -2076 31207 -2024
rect 30704 -2189 30756 -2137
rect 30768 -2189 30820 -2137
rect 31155 -2140 31207 -2088
rect 36790 -2162 36842 -2110
rect 36854 -2162 36906 -2110
rect 29412 -2554 29464 -2502
rect 29476 -2554 29528 -2502
rect 29643 -2530 29695 -2478
rect 29709 -2530 29761 -2478
rect 30439 -3194 30491 -3142
rect 30439 -3258 30491 -3206
rect 30285 -3386 30337 -3334
rect 30285 -3452 30337 -3400
rect 30377 -3423 30429 -3371
rect 30377 -3487 30429 -3435
rect 27192 -3762 27244 -3710
rect 27192 -3831 27244 -3779
rect 27192 -3900 27244 -3848
rect 28685 -4007 28737 -3955
rect 28768 -4007 28820 -3955
rect 28851 -4007 28903 -3955
rect 26087 -4079 26139 -4027
rect 26292 -4079 26344 -4027
rect 26087 -4143 26139 -4091
rect 26292 -4143 26344 -4091
rect 26328 -4242 26380 -4190
rect 26328 -4308 26380 -4256
rect 27288 -4329 27340 -4277
rect 27288 -4393 27340 -4341
rect 28153 -4568 28205 -4516
rect 28153 -4632 28205 -4580
rect 28685 -4534 28737 -4482
rect 28778 -4534 28830 -4482
rect 28870 -4534 28922 -4482
rect 28685 -4612 28737 -4560
rect 28778 -4612 28830 -4560
rect 28870 -4612 28922 -4560
rect 27668 -4806 27720 -4754
rect 27732 -4806 27784 -4754
rect 27192 -5111 27244 -5059
rect 27192 -5175 27244 -5123
rect 29486 -5263 29538 -5211
rect 29550 -5263 29602 -5211
rect 26110 -5573 26162 -5521
rect 26822 -5516 26874 -5464
rect 26110 -5637 26162 -5585
rect 26822 -5580 26874 -5528
rect 31155 -2242 31207 -2190
rect 31887 -2226 31939 -2174
rect 31951 -2226 32003 -2174
rect 31155 -2306 31207 -2254
rect 31155 -2400 31207 -2348
rect 32238 -2352 32290 -2300
rect 32302 -2352 32354 -2300
rect 33984 -2302 34036 -2250
rect 34048 -2302 34100 -2250
rect 36437 -2383 36489 -2331
rect 36501 -2383 36553 -2331
rect 31155 -2464 31207 -2412
rect 34581 -2494 34633 -2442
rect 34645 -2494 34697 -2442
rect 34340 -2550 34392 -2498
rect 34404 -2550 34456 -2498
rect 31174 -2632 31226 -2580
rect 31174 -2696 31226 -2644
rect 31393 -2653 31445 -2601
rect 31393 -2717 31445 -2665
rect 32825 -2844 32877 -2792
rect 32889 -2844 32941 -2792
rect 33853 -2844 33905 -2792
rect 33917 -2844 33969 -2792
rect 32772 -3168 32824 -3116
rect 31174 -3236 31226 -3184
rect 32772 -3232 32824 -3180
rect 31174 -3300 31226 -3248
rect 31174 -3417 31226 -3365
rect 31174 -3481 31226 -3429
rect 33022 -3495 33074 -3443
rect 33086 -3495 33138 -3443
rect 31009 -3647 31061 -3595
rect 31009 -3711 31061 -3659
rect 31175 -3647 31227 -3595
rect 31175 -3711 31227 -3659
rect 31911 -3647 31963 -3595
rect 31911 -3711 31963 -3659
rect 34387 -3657 34439 -3605
rect 31325 -3770 31377 -3718
rect 34387 -3721 34439 -3669
rect 34495 -3625 34547 -3573
rect 34495 -3689 34547 -3637
rect 31174 -3889 31226 -3837
rect 31325 -3834 31377 -3782
rect 35884 -3816 35936 -3764
rect 35948 -3816 36000 -3764
rect 31174 -3953 31226 -3901
rect 31801 -3940 31853 -3888
rect 31865 -3940 31917 -3888
rect 32765 -3955 32817 -3903
rect 32829 -3955 32881 -3903
rect 34357 -3908 34409 -3856
rect 34421 -3908 34473 -3856
rect 35884 -4140 35936 -4088
rect 35948 -4140 36000 -4088
rect 32730 -4470 32782 -4418
rect 32794 -4470 32846 -4418
rect 34317 -4621 34369 -4569
rect 34381 -4621 34433 -4569
rect 32308 -4848 32360 -4796
rect 33618 -4686 33670 -4634
rect 35057 -4637 35109 -4585
rect 33618 -4750 33670 -4698
rect 35057 -4701 35109 -4649
rect 32308 -4912 32360 -4860
rect 34782 -4866 34834 -4814
rect 34846 -4866 34898 -4814
rect 35252 -4908 35304 -4856
rect 35316 -4908 35368 -4856
rect 35970 -4924 36022 -4872
rect 36034 -4924 36086 -4872
rect 32991 -5332 33043 -5280
rect 32250 -5402 32302 -5350
rect 32314 -5402 32366 -5350
rect 32991 -5396 33043 -5344
rect 30774 -5569 30826 -5517
rect 27687 -5643 27739 -5591
rect 27751 -5643 27803 -5591
rect 30774 -5633 30826 -5581
rect 26506 -5932 26558 -5880
rect 26386 -5998 26438 -5946
rect 26506 -5996 26558 -5944
rect 26599 -5875 26651 -5823
rect 27197 -5873 27249 -5821
rect 27261 -5873 27313 -5821
rect 26599 -5939 26651 -5887
rect 32299 -5879 32351 -5827
rect 31149 -5945 31201 -5893
rect 31213 -5945 31265 -5893
rect 32299 -5943 32351 -5891
rect 32416 -5881 32468 -5829
rect 32488 -5881 32540 -5829
rect 32416 -5947 32468 -5895
rect 32488 -5947 32540 -5895
rect 38121 -5954 38173 -5902
rect 26386 -6062 26438 -6010
rect 31311 -6025 31363 -5973
rect 31375 -6025 31427 -5973
rect 30733 -6081 30785 -6029
rect 30797 -6081 30849 -6029
rect 33157 -6039 33209 -5987
rect 38121 -6018 38173 -5966
rect 32643 -6151 32695 -6099
rect 33157 -6103 33209 -6051
rect 38207 -6071 38259 -6019
rect 38207 -6135 38259 -6083
rect 32643 -6215 32695 -6163
<< metal2 >>
rect 26499 327 26924 333
rect 26551 275 26872 327
rect 26499 263 26924 275
rect 26551 211 26872 263
rect 26499 205 26924 211
rect 27871 33 27923 39
rect 27871 -31 27923 -19
rect 26218 -721 26444 -715
rect 26270 -766 26444 -721
tri 26444 -766 26495 -715 sw
rect 26270 -769 26495 -766
tri 26495 -769 26498 -766 sw
rect 26270 -773 26498 -769
rect 26218 -787 26498 -773
rect 26270 -790 26498 -787
tri 26498 -790 26519 -769 sw
rect 26270 -839 26666 -790
rect 26218 -842 26666 -839
rect 26718 -842 26746 -790
rect 26798 -842 26825 -790
rect 26877 -842 26924 -790
rect 26218 -845 26924 -842
tri 26390 -847 26392 -845 ne
rect 26392 -847 26924 -845
tri 26392 -868 26413 -847 ne
rect 26413 -868 26924 -847
tri 26413 -920 26465 -868 ne
rect 26465 -920 26666 -868
rect 26718 -920 26746 -868
rect 26798 -920 26825 -868
rect 26877 -920 26924 -868
rect 27871 -913 27923 -83
rect 33819 -87 33916 -78
tri 33717 -134 33721 -130 ne
rect 33721 -134 33819 -130
tri 33721 -208 33795 -134 ne
rect 33795 -143 33819 -134
rect 33875 -143 33916 -87
rect 33795 -167 33916 -143
rect 33795 -208 33819 -167
tri 33795 -232 33819 -208 ne
rect 33875 -208 33916 -167
tri 33916 -208 33990 -134 sw
rect 33875 -223 33967 -208
rect 33819 -232 33967 -223
tri 33967 -232 33990 -208 nw
rect 27984 -702 29111 -632
rect 27984 -707 28189 -702
tri 28189 -707 28194 -702 nw
tri 28270 -707 28275 -702 ne
rect 28275 -707 29111 -702
tri 29111 -707 29186 -632 sw
rect 27984 -714 28182 -707
tri 28182 -714 28189 -707 nw
tri 28275 -714 28282 -707 ne
rect 28282 -714 28324 -707
rect 27984 -763 28133 -714
tri 28133 -763 28182 -714 nw
tri 28282 -756 28324 -714 ne
rect 28784 -714 29140 -708
rect 27984 -766 28130 -763
tri 28130 -766 28133 -763 nw
rect 27984 -769 28127 -766
tri 28127 -769 28130 -766 nw
rect 28205 -769 28257 -763
rect 27984 -847 28112 -769
tri 28112 -784 28127 -769 nw
rect 27984 -899 27990 -847
rect 28042 -899 28054 -847
rect 28106 -899 28112 -847
rect 28205 -833 28257 -821
rect 28784 -766 28786 -714
rect 28838 -766 28886 -714
rect 28938 -766 28986 -714
rect 29038 -766 29086 -714
rect 29138 -766 29140 -714
rect 28784 -778 29140 -766
rect 28784 -830 28786 -778
rect 28838 -830 28886 -778
rect 28938 -830 28986 -778
rect 29038 -830 29086 -778
rect 29138 -830 29140 -778
rect 28784 -836 29140 -830
rect 28257 -885 29762 -871
tri 27871 -915 27873 -913 ne
rect 27873 -915 27923 -913
tri 27923 -915 27925 -913 sw
tri 26632 -923 26635 -920 ne
rect 26635 -923 26924 -920
tri 27873 -923 27881 -915 ne
rect 27881 -923 27925 -915
tri 27925 -923 27933 -915 sw
rect 28205 -923 29762 -885
rect 29814 -923 29826 -871
rect 29878 -923 29884 -871
tri 26635 -1060 26772 -923 ne
rect 26772 -1652 26924 -923
tri 27881 -965 27923 -923 ne
rect 27923 -965 27933 -923
tri 27923 -967 27925 -965 ne
rect 27925 -967 27933 -965
tri 27933 -967 27977 -923 sw
tri 27925 -995 27953 -967 ne
rect 27953 -995 28437 -967
rect 29758 -1065 29810 -1059
rect 29758 -1129 29810 -1117
rect 27730 -1164 27933 -1158
rect 27730 -1216 27731 -1164
rect 27783 -1216 27805 -1164
rect 27857 -1216 27933 -1164
rect 27730 -1286 27933 -1216
rect 27730 -1338 27731 -1286
rect 27783 -1338 27805 -1286
rect 27857 -1338 27933 -1286
rect 27730 -1660 27933 -1338
rect 28145 -1465 28151 -1413
rect 28203 -1465 28215 -1413
rect 28267 -1465 28273 -1413
tri 28183 -1511 28229 -1465 ne
tri 26343 -2391 26377 -2357 sw
rect 26343 -2464 26356 -2443
tri 26356 -2464 26377 -2443 nw
rect 26343 -2472 26348 -2464
tri 26348 -2472 26356 -2464 nw
tri 26667 -2472 26675 -2464 sw
tri 26343 -2477 26348 -2472 nw
tri 26634 -2477 26639 -2472 se
tri 26633 -2478 26634 -2477 se
rect 26634 -2478 26639 -2477
tri 26613 -2498 26633 -2478 se
rect 26633 -2498 26639 -2478
rect 26667 -2478 26675 -2472
tri 26675 -2478 26681 -2472 sw
rect 26667 -2498 26681 -2478
tri 26681 -2498 26701 -2478 sw
tri 26306 -4007 26315 -3998 se
rect 26315 -4007 26343 -3403
tri 26300 -4013 26306 -4007 se
rect 26306 -4013 26343 -4007
tri 26292 -4021 26300 -4013 se
rect 26300 -4015 26343 -4013
rect 27192 -3710 27244 -3704
rect 27192 -3779 27244 -3762
rect 27192 -3848 27244 -3831
tri 26343 -4015 26344 -4014 sw
rect 26300 -4021 26344 -4015
rect 26087 -4027 26139 -4021
rect 26087 -4091 26139 -4079
rect 26087 -4149 26139 -4143
rect 26292 -4027 26344 -4021
rect 26292 -4091 26344 -4079
rect 26292 -4149 26344 -4143
tri 26087 -4172 26110 -4149 ne
rect 26110 -5515 26138 -4149
tri 26138 -4150 26139 -4149 nw
rect 26324 -4190 26380 -4184
rect 26324 -4193 26328 -4190
rect 26324 -4256 26380 -4249
rect 26324 -4273 26328 -4256
rect 26324 -4338 26380 -4329
tri 26771 -4605 26773 -4603 se
rect 27192 -5059 27244 -3900
rect 27192 -5123 27244 -5111
rect 27192 -5181 27244 -5175
rect 27288 -4277 27340 -4271
rect 27288 -4341 27340 -4329
tri 27273 -5332 27288 -5317 se
rect 27288 -5332 27340 -4393
tri 28185 -4418 28229 -4374 se
rect 28229 -4418 28257 -1465
tri 28257 -1481 28273 -1465 nw
rect 29758 -2231 29810 -1181
tri 33637 -2018 33664 -1991 se
rect 33664 -2018 37134 -1991
tri 37134 -2018 37161 -1991 sw
rect 31155 -2024 31207 -2018
tri 33600 -2055 33637 -2018 se
rect 33637 -2019 37161 -2018
rect 33637 -2055 33674 -2019
tri 33674 -2055 33710 -2019 nw
tri 37096 -2049 37126 -2019 ne
rect 37126 -2049 37161 -2019
tri 36621 -2055 36627 -2049 se
rect 36627 -2055 37032 -2049
tri 37032 -2055 37038 -2049 sw
tri 37126 -2055 37132 -2049 ne
rect 37132 -2055 37161 -2049
tri 37161 -2055 37198 -2018 sw
tri 33590 -2065 33600 -2055 se
rect 33600 -2065 33664 -2055
tri 33664 -2065 33674 -2055 nw
tri 36611 -2065 36621 -2055 se
rect 36621 -2057 37038 -2055
tri 37038 -2057 37040 -2055 sw
tri 37132 -2057 37134 -2055 ne
rect 37134 -2057 37198 -2055
rect 36621 -2065 37040 -2057
tri 37040 -2065 37048 -2057 sw
tri 37134 -2065 37142 -2057 ne
rect 37142 -2065 37198 -2057
rect 31155 -2088 31207 -2076
rect 30698 -2137 31155 -2118
rect 30698 -2189 30704 -2137
rect 30756 -2189 30768 -2137
rect 30820 -2140 31155 -2137
tri 33545 -2110 33590 -2065 se
rect 33590 -2110 33619 -2065
tri 33619 -2110 33664 -2065 nw
tri 36599 -2077 36611 -2065 se
rect 36611 -2069 37048 -2065
tri 37048 -2069 37052 -2065 sw
rect 36611 -2077 37052 -2069
tri 37142 -2075 37152 -2065 ne
tri 36574 -2102 36599 -2077 se
rect 36599 -2102 36627 -2077
tri 36627 -2102 36652 -2077 nw
tri 36955 -2102 36980 -2077 ne
rect 36980 -2102 37052 -2077
tri 36566 -2110 36574 -2102 se
rect 36574 -2110 36619 -2102
tri 36619 -2110 36627 -2102 nw
tri 36980 -2110 36988 -2102 ne
rect 36988 -2110 37052 -2102
rect 30820 -2146 31207 -2140
tri 33522 -2133 33545 -2110 se
rect 33545 -2133 33596 -2110
tri 33596 -2133 33619 -2110 nw
tri 36562 -2114 36566 -2110 se
rect 36566 -2114 36574 -2110
rect 33819 -2123 34143 -2114
rect 33522 -2146 33583 -2133
tri 33583 -2146 33596 -2133 nw
rect 30820 -2162 30853 -2146
tri 30853 -2162 30869 -2146 nw
rect 30820 -2174 30841 -2162
tri 30841 -2174 30853 -2162 nw
rect 30820 -2189 30826 -2174
tri 30826 -2189 30841 -2174 nw
rect 31155 -2190 31207 -2184
rect 29758 -2242 31155 -2231
rect 29758 -2254 31207 -2242
rect 31881 -2226 31887 -2174
rect 31939 -2226 31951 -2174
rect 32003 -2226 32009 -2174
tri 31881 -2250 31905 -2226 ne
rect 31905 -2250 31985 -2226
tri 31985 -2250 32009 -2226 nw
rect 29758 -2283 31155 -2254
tri 31905 -2256 31911 -2250 ne
rect 31911 -2256 31979 -2250
tri 31979 -2256 31985 -2250 nw
rect 31155 -2312 31207 -2306
rect 31155 -2348 31207 -2342
rect 31155 -2412 31207 -2400
tri 30743 -2442 30756 -2429 se
rect 30756 -2442 31155 -2429
tri 30721 -2464 30743 -2442 se
rect 30743 -2457 31155 -2442
rect 30743 -2464 30779 -2457
tri 30779 -2464 30786 -2457 nw
tri 30707 -2478 30721 -2464 se
rect 30721 -2478 30765 -2464
tri 30765 -2478 30779 -2464 nw
rect 31155 -2470 31207 -2464
rect 29406 -2554 29412 -2502
rect 29464 -2554 29476 -2502
rect 29528 -2530 29534 -2502
tri 29534 -2530 29558 -2506 sw
rect 29637 -2530 29643 -2478
rect 29695 -2530 29709 -2478
rect 29761 -2494 30749 -2478
tri 30749 -2494 30765 -2478 nw
rect 29761 -2498 30745 -2494
tri 30745 -2498 30749 -2494 nw
rect 29761 -2506 30737 -2498
tri 30737 -2506 30745 -2498 nw
rect 29761 -2530 29767 -2506
tri 29767 -2530 29791 -2506 nw
rect 29528 -2550 29558 -2530
tri 29558 -2550 29578 -2530 sw
rect 29528 -2554 29578 -2550
tri 29578 -2554 29582 -2550 sw
tri 29530 -2574 29550 -2554 ne
rect 29550 -2574 29582 -2554
tri 29582 -2574 29602 -2554 sw
tri 29550 -2580 29556 -2574 ne
rect 29556 -2580 29602 -2574
tri 29602 -2580 29608 -2574 sw
rect 31174 -2580 31226 -2574
tri 29556 -2606 29582 -2580 ne
rect 29582 -2587 29608 -2580
tri 29608 -2587 29615 -2580 sw
rect 29582 -2606 31174 -2587
tri 29582 -2615 29591 -2606 ne
rect 29591 -2615 31174 -2606
rect 31174 -2644 31226 -2632
rect 31174 -2702 31226 -2696
rect 31393 -2601 31445 -2595
rect 31393 -2665 31445 -2653
rect 31393 -2723 31445 -2717
rect 30439 -3142 30491 -3136
rect 30439 -3206 30491 -3194
rect 31174 -3184 31226 -3178
rect 30491 -3236 31174 -3212
rect 30491 -3248 31226 -3236
rect 30491 -3258 31174 -3248
rect 30439 -3264 31174 -3258
rect 31174 -3306 31226 -3300
rect 30285 -3334 30337 -3328
rect 31174 -3365 31226 -3359
rect 30285 -3400 30337 -3386
rect 30285 -3458 30337 -3452
rect 30377 -3371 30429 -3365
rect 30429 -3417 31174 -3392
rect 30429 -3423 31226 -3417
rect 30377 -3429 31226 -3423
rect 30377 -3435 31174 -3429
rect 30304 -3889 30332 -3458
rect 30429 -3444 31174 -3435
rect 31174 -3487 31226 -3481
rect 30377 -3493 30429 -3487
rect 31009 -3595 31227 -3589
rect 31061 -3647 31175 -3595
rect 31009 -3659 31227 -3647
rect 31061 -3711 31175 -3659
rect 31009 -3717 31227 -3711
rect 31325 -3718 31377 -3712
rect 31325 -3782 31377 -3770
rect 31174 -3837 31226 -3831
tri 30332 -3889 30343 -3878 sw
rect 30304 -3901 30343 -3889
tri 30343 -3901 30355 -3889 sw
rect 31174 -3901 31226 -3889
rect 30304 -3912 30355 -3901
tri 30355 -3912 30366 -3901 sw
tri 28176 -4427 28185 -4418 se
rect 28185 -4422 28257 -4418
rect 28185 -4427 28252 -4422
tri 28252 -4427 28257 -4422 nw
rect 28679 -3955 28928 -3934
rect 30304 -3940 31174 -3912
rect 28679 -4007 28685 -3955
rect 28737 -4007 28768 -3955
rect 28820 -4007 28851 -3955
rect 28903 -4007 28928 -3955
rect 31174 -3959 31226 -3953
rect 28176 -4470 28209 -4427
tri 28209 -4470 28252 -4427 nw
tri 28153 -4510 28176 -4487 se
rect 28176 -4510 28205 -4470
tri 28205 -4474 28209 -4470 nw
rect 28153 -4516 28205 -4510
rect 28153 -4580 28205 -4568
rect 28679 -4482 28928 -4007
tri 31299 -4088 31325 -4062 se
rect 31325 -4084 31377 -3834
rect 31325 -4088 31373 -4084
tri 31373 -4088 31377 -4084 nw
tri 31251 -4136 31299 -4088 se
rect 31299 -4136 31325 -4088
tri 31325 -4136 31373 -4088 nw
tri 31247 -4140 31251 -4136 se
rect 31251 -4140 31321 -4136
tri 31321 -4140 31325 -4136 nw
rect 28679 -4534 28685 -4482
rect 28737 -4534 28778 -4482
rect 28830 -4534 28870 -4482
rect 28922 -4534 28928 -4482
rect 28679 -4560 28928 -4534
rect 28679 -4612 28685 -4560
rect 28737 -4612 28778 -4560
rect 28830 -4612 28870 -4560
rect 28922 -4612 28928 -4560
tri 31243 -4144 31247 -4140 se
rect 31247 -4144 31317 -4140
tri 31317 -4144 31321 -4140 nw
rect 28153 -4638 28205 -4632
rect 27662 -4806 27668 -4754
rect 27720 -4806 27732 -4754
rect 27784 -4806 27790 -4754
tri 27261 -5344 27273 -5332 se
rect 27273 -5339 27340 -5332
rect 27273 -5344 27335 -5339
tri 27335 -5344 27340 -5339 nw
tri 27255 -5350 27261 -5344 se
rect 27261 -5350 27329 -5344
tri 27329 -5350 27335 -5344 nw
tri 27236 -5369 27255 -5350 se
rect 27255 -5369 27310 -5350
tri 27310 -5369 27329 -5350 nw
rect 26822 -5464 26874 -5458
rect 26110 -5521 26162 -5515
rect 26110 -5585 26162 -5573
rect 26110 -5643 26162 -5637
rect 26822 -5528 26874 -5516
rect 26822 -5763 26874 -5580
rect 26599 -5823 26651 -5817
rect 27236 -5821 27288 -5369
tri 27288 -5391 27310 -5369 nw
rect 27737 -5591 27765 -4806
rect 29480 -5263 29486 -5211
rect 29538 -5263 29550 -5211
rect 29602 -5263 29608 -5211
tri 28317 -5402 28330 -5389 se
tri 28296 -5423 28317 -5402 se
rect 28317 -5423 28330 -5402
rect 30774 -5517 30826 -5511
rect 30774 -5581 30826 -5569
rect 27681 -5643 27687 -5591
rect 27739 -5643 27751 -5591
rect 27803 -5643 27809 -5591
rect 30774 -5639 30826 -5633
rect 26506 -5880 26558 -5874
rect 26384 -5923 26440 -5914
rect 26384 -5998 26386 -5979
rect 26438 -5998 26440 -5979
rect 26384 -6003 26440 -5998
rect 26506 -5944 26558 -5932
rect 27191 -5873 27197 -5821
rect 27249 -5873 27261 -5821
rect 27313 -5873 27319 -5821
rect 26599 -5887 26651 -5875
rect 26599 -5945 26651 -5939
rect 26506 -6002 26558 -5996
rect 30798 -6029 30826 -5639
rect 31243 -5893 31271 -4144
tri 31271 -4190 31317 -4144 nw
rect 31143 -5945 31149 -5893
rect 31201 -5945 31213 -5893
rect 31265 -5945 31271 -5893
rect 31405 -5973 31433 -2723
rect 31911 -3595 31963 -2256
tri 31963 -2272 31979 -2256 nw
rect 32232 -2352 32238 -2300
rect 32290 -2352 32302 -2300
rect 32354 -2352 32360 -2300
rect 31911 -3659 31963 -3647
rect 31911 -3717 31963 -3711
rect 31795 -3940 31801 -3888
rect 31853 -3940 31865 -3888
rect 31917 -3940 31923 -3888
tri 31795 -3955 31810 -3940 ne
rect 31810 -3955 31908 -3940
tri 31908 -3955 31923 -3940 nw
tri 31810 -3974 31829 -3955 ne
rect 31829 -3974 31889 -3955
tri 31889 -3974 31908 -3955 nw
tri 31829 -3982 31837 -3974 ne
rect 31837 -4912 31889 -3974
rect 32308 -4796 32360 -2352
rect 33522 -2653 33574 -2146
tri 33574 -2155 33583 -2146 nw
rect 33875 -2155 34143 -2123
tri 34143 -2155 34184 -2114 sw
tri 36521 -2155 36562 -2114 se
rect 36562 -2155 36574 -2114
tri 36574 -2155 36619 -2110 nw
rect 33875 -2162 34184 -2155
tri 34184 -2162 34191 -2155 sw
tri 36514 -2162 36521 -2155 se
rect 36521 -2162 36567 -2155
tri 36567 -2162 36574 -2155 nw
rect 36784 -2162 36790 -2110
rect 36842 -2162 36854 -2110
rect 36906 -2162 36912 -2110
tri 36988 -2122 37000 -2110 ne
rect 33875 -2166 34191 -2162
rect 33819 -2203 33875 -2179
tri 34121 -2187 34142 -2166 ne
rect 34142 -2187 34191 -2166
tri 34191 -2187 34216 -2162 sw
tri 34142 -2188 34143 -2187 ne
rect 34143 -2188 34216 -2187
tri 34143 -2209 34164 -2188 ne
rect 33819 -2268 33875 -2259
rect 33978 -2302 33984 -2250
rect 34036 -2302 34048 -2250
rect 34100 -2302 34106 -2250
tri 33574 -2653 33596 -2631 sw
tri 33522 -2727 33596 -2653 ne
tri 33596 -2727 33670 -2653 sw
tri 33596 -2749 33618 -2727 ne
rect 32772 -2844 32825 -2792
rect 32877 -2844 32889 -2792
rect 32941 -2844 32947 -2792
rect 32772 -3116 32824 -2844
rect 32772 -3180 32824 -3168
rect 32772 -3238 32824 -3232
rect 33016 -3495 33022 -3443
rect 33074 -3495 33086 -3443
rect 33138 -3472 33223 -3443
tri 33223 -3472 33252 -3443 sw
rect 33138 -3495 33252 -3472
tri 33221 -3526 33252 -3495 ne
tri 33252 -3526 33306 -3472 sw
tri 33252 -3554 33280 -3526 ne
rect 33280 -3554 33483 -3526
rect 32759 -3955 32765 -3903
rect 32817 -3955 32829 -3903
rect 32881 -3955 32887 -3903
rect 32724 -4470 32730 -4418
rect 32782 -4470 32794 -4418
rect 32846 -4470 32852 -4418
rect 32308 -4860 32360 -4848
tri 31889 -4912 31901 -4900 sw
rect 31837 -4924 31901 -4912
tri 31901 -4924 31913 -4912 sw
rect 32308 -4918 32360 -4912
rect 32748 -4900 32800 -4470
tri 32800 -4900 32813 -4887 sw
rect 32748 -4908 32813 -4900
tri 32813 -4908 32821 -4900 sw
rect 32748 -4909 32821 -4908
tri 32748 -4918 32757 -4909 ne
rect 32757 -4918 32821 -4909
tri 32757 -4924 32763 -4918 ne
rect 32763 -4924 32821 -4918
tri 32821 -4924 32837 -4908 sw
rect 31837 -4942 31913 -4924
tri 31913 -4942 31931 -4924 sw
tri 32763 -4942 32781 -4924 ne
rect 32781 -4942 32837 -4924
tri 32837 -4942 32855 -4924 sw
tri 31837 -5036 31931 -4942 ne
tri 31931 -5036 32025 -4942 sw
tri 32781 -4953 32792 -4942 ne
rect 32792 -4953 32855 -4942
tri 32855 -4953 32866 -4942 sw
tri 32792 -4961 32800 -4953 ne
rect 32800 -4961 32866 -4953
tri 32800 -4975 32814 -4961 ne
tri 31931 -5130 32025 -5036 ne
tri 32025 -5130 32119 -5036 sw
tri 32025 -5224 32119 -5130 ne
tri 32119 -5224 32213 -5130 sw
tri 32792 -5155 32814 -5133 se
rect 32814 -5155 32866 -4961
rect 33455 -5018 33483 -3554
rect 33618 -4634 33670 -2727
rect 33847 -2844 33853 -2792
rect 33905 -2844 33917 -2792
rect 33969 -2844 33975 -2792
rect 33847 -3131 33899 -2844
tri 33899 -2878 33933 -2844 nw
tri 33847 -3138 33854 -3131 ne
rect 33618 -4698 33670 -4686
rect 33618 -4756 33670 -4750
tri 33847 -3247 33854 -3240 se
rect 33854 -3247 33899 -3131
rect 33847 -4887 33899 -3247
rect 34055 -4421 34094 -2302
tri 34150 -2383 34164 -2369 se
rect 34164 -2383 34216 -2188
tri 36475 -2201 36514 -2162 se
rect 36514 -2201 36528 -2162
tri 36528 -2201 36567 -2162 nw
rect 36475 -2331 36503 -2201
tri 36503 -2226 36528 -2201 nw
rect 36431 -2383 36437 -2331
rect 36489 -2383 36501 -2331
rect 36553 -2383 36559 -2331
rect 36848 -2366 36900 -2162
rect 37000 -2367 37052 -2110
tri 34142 -2391 34150 -2383 se
rect 34150 -2391 34216 -2383
tri 34122 -2411 34142 -2391 se
rect 34142 -2411 34193 -2391
rect 34122 -2414 34193 -2411
tri 34193 -2414 34216 -2391 nw
rect 37152 -2385 37198 -2065
rect 34122 -4361 34169 -2414
tri 34169 -2438 34193 -2414 nw
tri 36660 -2438 36684 -2414 ne
rect 36684 -2438 36694 -2414
tri 36746 -2436 36768 -2414 nw
rect 37152 -2431 37906 -2385
tri 36684 -2442 36688 -2438 ne
rect 36688 -2442 36694 -2438
rect 34575 -2494 34581 -2442
rect 34633 -2494 34645 -2442
rect 34697 -2494 34703 -2442
tri 36688 -2448 36694 -2442 ne
rect 34575 -2498 34699 -2494
tri 34699 -2498 34703 -2494 nw
rect 34334 -2550 34340 -2498
rect 34392 -2550 34404 -2498
rect 34456 -2550 34462 -2498
rect 34575 -2550 34647 -2498
tri 34647 -2550 34699 -2498 nw
tri 34501 -3095 34575 -3021 se
rect 34575 -3043 34627 -2550
tri 34627 -2570 34647 -2550 nw
tri 34575 -3095 34627 -3043 nw
rect 34686 -3095 34738 -3030
tri 34738 -3095 34747 -3086 sw
tri 34495 -3101 34501 -3095 se
rect 34501 -3101 34569 -3095
tri 34569 -3101 34575 -3095 nw
rect 34686 -3101 34747 -3095
tri 34747 -3101 34753 -3095 sw
rect 34495 -3573 34547 -3101
tri 34547 -3123 34569 -3101 nw
rect 34686 -3108 34753 -3101
tri 34686 -3123 34701 -3108 ne
rect 34701 -3123 34753 -3108
tri 34753 -3123 34775 -3101 sw
tri 34701 -3142 34720 -3123 ne
rect 34720 -3142 34775 -3123
tri 34775 -3142 34794 -3123 sw
tri 34720 -3160 34738 -3142 ne
rect 34738 -3160 34794 -3142
tri 34738 -3216 34794 -3160 ne
tri 34794 -3216 34868 -3142 sw
tri 34794 -3261 34839 -3216 ne
rect 34387 -3605 34439 -3599
rect 34387 -3669 34439 -3657
rect 34495 -3637 34547 -3625
rect 34495 -3695 34547 -3689
rect 34658 -3581 34714 -3572
rect 34658 -3661 34714 -3637
rect 34387 -3727 34439 -3721
rect 34658 -3816 34714 -3717
rect 34839 -3759 34868 -3216
tri 34839 -3764 34844 -3759 ne
rect 34844 -3764 34868 -3759
tri 34868 -3764 34918 -3714 sw
tri 34844 -3788 34868 -3764 ne
rect 34868 -3788 35884 -3764
tri 34868 -3810 34890 -3788 ne
rect 34890 -3810 35884 -3788
tri 34714 -3816 34720 -3810 sw
tri 34890 -3816 34896 -3810 ne
rect 34896 -3816 35884 -3810
rect 35936 -3816 35948 -3764
rect 36000 -3816 36006 -3764
rect 34658 -3828 34720 -3816
tri 34658 -3856 34686 -3828 ne
rect 34686 -3856 34720 -3828
rect 34351 -3908 34357 -3856
rect 34409 -3908 34421 -3856
rect 34473 -3908 34479 -3856
tri 34686 -3862 34692 -3856 ne
rect 34692 -3862 34720 -3856
tri 34720 -3862 34766 -3816 sw
tri 35815 -3862 35861 -3816 ne
rect 35861 -3862 36006 -3816
tri 34692 -3868 34698 -3862 ne
rect 34698 -3868 35603 -3862
tri 35603 -3868 35609 -3862 sw
tri 35861 -3868 35867 -3862 ne
rect 35867 -3868 36006 -3862
tri 34698 -3884 34714 -3868 ne
rect 34714 -3884 35609 -3868
tri 34714 -3888 34718 -3884 ne
rect 34718 -3888 35609 -3884
tri 35609 -3888 35629 -3868 sw
tri 35867 -3879 35878 -3868 ne
tri 34718 -3903 34733 -3888 ne
rect 34733 -3903 35629 -3888
tri 35629 -3903 35644 -3888 sw
tri 34733 -3908 34738 -3903 ne
rect 34738 -3908 35644 -3903
tri 35644 -3908 35649 -3903 sw
tri 34351 -3944 34387 -3908 ne
rect 34387 -4088 34439 -3908
tri 34439 -3948 34479 -3908 nw
tri 34738 -3914 34744 -3908 ne
rect 34744 -3914 35649 -3908
tri 35581 -3942 35609 -3914 ne
rect 35609 -3942 35649 -3914
tri 35649 -3942 35683 -3908 sw
tri 35609 -3948 35615 -3942 ne
rect 35615 -3948 35683 -3942
tri 35615 -3964 35631 -3948 ne
rect 35631 -4029 35683 -3948
tri 35631 -4052 35654 -4029 ne
rect 35654 -4052 35683 -4029
tri 35683 -4052 35728 -4007 sw
tri 35654 -4072 35674 -4052 ne
rect 35674 -4072 35728 -4052
tri 35728 -4072 35748 -4052 sw
tri 34439 -4088 34455 -4072 sw
tri 35674 -4081 35683 -4072 ne
rect 35683 -4081 35748 -4072
tri 35683 -4088 35690 -4081 ne
rect 35690 -4088 35748 -4081
tri 35748 -4088 35764 -4072 sw
rect 35878 -4088 36006 -3868
rect 34387 -4090 34455 -4088
tri 34455 -4090 34457 -4088 sw
tri 35690 -4090 35692 -4088 ne
rect 35692 -4090 35764 -4088
tri 35764 -4090 35766 -4088 sw
rect 34387 -4094 34457 -4090
tri 34387 -4140 34433 -4094 ne
rect 34433 -4140 34457 -4094
tri 34457 -4140 34507 -4090 sw
tri 35692 -4126 35728 -4090 ne
rect 35728 -4126 35766 -4090
tri 35766 -4126 35802 -4090 sw
tri 35728 -4140 35742 -4126 ne
rect 35742 -4140 35802 -4126
tri 35802 -4140 35816 -4126 sw
rect 35878 -4140 35884 -4088
rect 35936 -4140 35948 -4088
rect 36000 -4140 36006 -4088
tri 34433 -4164 34457 -4140 ne
rect 34457 -4164 34507 -4140
tri 34507 -4164 34531 -4140 sw
tri 35742 -4164 35766 -4140 ne
rect 35766 -4164 35816 -4140
tri 35816 -4164 35840 -4140 sw
tri 34457 -4216 34509 -4164 ne
rect 34509 -4200 35687 -4164
tri 35687 -4200 35723 -4164 sw
tri 35766 -4200 35802 -4164 ne
rect 35802 -4200 35840 -4164
tri 35840 -4200 35876 -4164 sw
rect 34509 -4216 35723 -4200
tri 35665 -4219 35668 -4216 ne
rect 35668 -4219 35723 -4216
tri 35723 -4219 35742 -4200 sw
tri 35802 -4207 35809 -4200 ne
rect 35809 -4207 35940 -4200
tri 35940 -4207 35947 -4200 sw
tri 35809 -4219 35821 -4207 ne
rect 35821 -4219 35947 -4207
tri 35947 -4219 35959 -4207 sw
tri 35668 -4238 35687 -4219 ne
rect 35687 -4238 35742 -4219
tri 35687 -4293 35742 -4238 ne
tri 35742 -4252 35775 -4219 sw
tri 35821 -4252 35854 -4219 ne
rect 35854 -4252 35959 -4219
rect 35742 -4293 35775 -4252
tri 35775 -4293 35816 -4252 sw
tri 35918 -4281 35947 -4252 ne
rect 35947 -4281 35959 -4252
tri 35959 -4281 36021 -4219 sw
tri 35947 -4293 35959 -4281 ne
rect 35959 -4293 36021 -4281
tri 36021 -4293 36033 -4281 sw
tri 35742 -4318 35767 -4293 ne
rect 35767 -4318 35816 -4293
tri 35499 -4334 35515 -4318 se
rect 35515 -4334 35715 -4318
tri 35715 -4334 35731 -4318 sw
tri 35767 -4334 35783 -4318 ne
rect 35783 -4334 35816 -4318
tri 34122 -4391 34152 -4361 ne
rect 34152 -4367 34169 -4361
tri 34169 -4367 34202 -4334 sw
tri 35497 -4336 35499 -4334 se
rect 35499 -4336 35731 -4334
tri 35731 -4336 35733 -4334 sw
tri 35783 -4336 35785 -4334 ne
rect 35785 -4336 35816 -4334
tri 35466 -4367 35497 -4336 se
rect 35497 -4350 35733 -4336
tri 35733 -4350 35747 -4336 sw
tri 35785 -4350 35799 -4336 ne
rect 35799 -4350 35816 -4336
rect 35497 -4364 35747 -4350
rect 35497 -4367 35515 -4364
rect 34152 -4391 34202 -4367
tri 34202 -4391 34226 -4367 sw
tri 35449 -4384 35466 -4367 se
rect 35466 -4384 35515 -4367
tri 35515 -4384 35535 -4364 nw
tri 35695 -4384 35715 -4364 ne
rect 35715 -4367 35747 -4364
tri 35747 -4367 35764 -4350 sw
tri 35799 -4367 35816 -4350 ne
tri 35816 -4367 35890 -4293 sw
tri 35959 -4355 36021 -4293 ne
rect 36021 -4355 36033 -4293
tri 36033 -4355 36095 -4293 sw
tri 36021 -4367 36033 -4355 ne
rect 36033 -4367 36095 -4355
tri 36095 -4367 36107 -4355 sw
rect 35715 -4384 35764 -4367
tri 35442 -4391 35449 -4384 se
rect 35449 -4391 35497 -4384
tri 34152 -4408 34169 -4391 ne
rect 34169 -4408 34226 -4391
tri 34169 -4415 34176 -4408 ne
rect 34176 -4415 34226 -4408
tri 34226 -4415 34250 -4391 sw
tri 35431 -4402 35442 -4391 se
rect 35442 -4402 35497 -4391
tri 35497 -4402 35515 -4384 nw
tri 35715 -4402 35733 -4384 ne
rect 35733 -4391 35764 -4384
tri 35764 -4391 35788 -4367 sw
tri 35816 -4391 35840 -4367 ne
rect 35840 -4391 35890 -4367
rect 35733 -4402 35788 -4391
tri 35788 -4402 35799 -4391 sw
tri 35840 -4402 35851 -4391 ne
rect 35851 -4402 35890 -4391
tri 35425 -4408 35431 -4402 se
rect 35431 -4408 35491 -4402
tri 35491 -4408 35497 -4402 nw
tri 35733 -4408 35739 -4402 ne
rect 35739 -4408 35799 -4402
rect 35425 -4415 35484 -4408
tri 35484 -4415 35491 -4408 nw
tri 35739 -4415 35746 -4408 ne
rect 35746 -4415 35799 -4408
tri 35799 -4415 35812 -4402 sw
tri 35851 -4415 35864 -4402 ne
rect 35864 -4415 35890 -4402
tri 34094 -4421 34100 -4415 sw
tri 34176 -4421 34182 -4415 ne
rect 34182 -4421 34250 -4415
tri 34250 -4421 34256 -4415 sw
rect 35425 -4421 35478 -4415
tri 35478 -4421 35484 -4415 nw
tri 35746 -4421 35752 -4415 ne
rect 35752 -4416 35812 -4415
tri 35812 -4416 35813 -4415 sw
tri 35864 -4416 35865 -4415 ne
rect 35865 -4416 35890 -4415
rect 35752 -4421 35813 -4416
tri 35813 -4421 35818 -4416 sw
tri 35865 -4421 35870 -4416 ne
rect 35870 -4421 35890 -4416
rect 34055 -4441 34100 -4421
tri 34100 -4441 34120 -4421 sw
tri 34182 -4441 34202 -4421 ne
rect 34202 -4441 34256 -4421
tri 34256 -4441 34276 -4421 sw
rect 34055 -4450 34120 -4441
tri 34055 -4495 34100 -4450 ne
rect 34100 -4470 34120 -4450
tri 34120 -4470 34149 -4441 sw
tri 34202 -4465 34226 -4441 ne
rect 34226 -4465 34276 -4441
tri 34276 -4465 34300 -4441 sw
tri 34226 -4470 34231 -4465 ne
rect 34231 -4470 34828 -4465
rect 34100 -4495 34149 -4470
tri 34149 -4495 34174 -4470 sw
tri 34231 -4495 34256 -4470 ne
rect 34256 -4495 34828 -4470
tri 34100 -4569 34174 -4495 ne
tri 34174 -4515 34194 -4495 sw
tri 34256 -4515 34276 -4495 ne
rect 34276 -4515 34828 -4495
rect 34174 -4517 34194 -4515
tri 34194 -4517 34196 -4515 sw
tri 34276 -4517 34278 -4515 ne
rect 34278 -4517 34828 -4515
rect 34174 -4565 34196 -4517
tri 34196 -4565 34244 -4517 sw
rect 34174 -4569 34244 -4565
tri 34244 -4569 34248 -4565 sw
tri 34174 -4621 34226 -4569 ne
rect 34226 -4621 34317 -4569
rect 34369 -4621 34381 -4569
rect 34433 -4621 34439 -4569
rect 34776 -4814 34828 -4517
rect 35057 -4574 35113 -4565
rect 35109 -4637 35113 -4630
rect 35057 -4649 35113 -4637
rect 35109 -4654 35113 -4649
rect 35057 -4719 35113 -4710
rect 34776 -4866 34782 -4814
rect 34834 -4866 34846 -4814
rect 34898 -4866 34904 -4814
tri 35096 -4866 35106 -4856 se
rect 35106 -4866 35252 -4856
tri 35080 -4882 35096 -4866 se
rect 35096 -4882 35252 -4866
tri 33899 -4887 33904 -4882 sw
tri 35075 -4887 35080 -4882 se
rect 35080 -4887 35252 -4882
rect 33847 -4900 33904 -4887
tri 33904 -4900 33917 -4887 sw
tri 35062 -4900 35075 -4887 se
rect 35075 -4900 35252 -4887
rect 33847 -4904 33917 -4900
tri 33847 -4908 33851 -4904 ne
rect 33851 -4908 33917 -4904
tri 33917 -4908 33925 -4900 sw
tri 35054 -4908 35062 -4900 se
rect 35062 -4908 35252 -4900
rect 35304 -4908 35316 -4856
rect 35368 -4908 35374 -4856
tri 33851 -4924 33867 -4908 ne
rect 33867 -4924 35112 -4908
tri 35112 -4924 35128 -4908 nw
tri 33867 -4937 33880 -4924 ne
rect 33880 -4937 35099 -4924
tri 35099 -4937 35112 -4924 nw
tri 33880 -4942 33885 -4937 ne
rect 33885 -4942 35080 -4937
tri 33885 -4956 33899 -4942 ne
rect 33899 -4956 35080 -4942
tri 35080 -4956 35099 -4937 nw
tri 33899 -4960 33903 -4956 ne
rect 33903 -4960 35076 -4956
tri 35076 -4960 35080 -4956 nw
tri 33483 -5018 33494 -5007 sw
rect 33455 -5040 33494 -5018
tri 33494 -5040 33516 -5018 sw
rect 33455 -5053 33516 -5040
tri 33455 -5092 33494 -5053 ne
rect 33494 -5092 33516 -5053
tri 33516 -5092 33568 -5040 sw
tri 35373 -5092 35425 -5040 se
rect 35425 -5060 35471 -4421
tri 35471 -4428 35478 -4421 nw
tri 35752 -4428 35759 -4421 ne
rect 35759 -4428 35818 -4421
tri 35759 -4441 35772 -4428 ne
rect 35772 -4441 35818 -4428
tri 35818 -4441 35838 -4421 sw
tri 35870 -4441 35890 -4421 ne
tri 35890 -4441 35964 -4367 sw
tri 36033 -4429 36095 -4367 ne
rect 36095 -4429 36107 -4367
tri 36107 -4429 36169 -4367 sw
tri 36095 -4441 36107 -4429 ne
rect 36107 -4441 36169 -4429
tri 36169 -4441 36181 -4429 sw
tri 35772 -4465 35796 -4441 ne
rect 35796 -4465 35838 -4441
tri 35838 -4465 35862 -4441 sw
tri 35890 -4465 35914 -4441 ne
rect 35914 -4465 35964 -4441
tri 35796 -4468 35799 -4465 ne
rect 35799 -4468 35862 -4465
tri 35862 -4468 35865 -4465 sw
tri 35914 -4468 35917 -4465 ne
rect 35917 -4468 35964 -4465
tri 35799 -4534 35865 -4468 ne
tri 35865 -4470 35867 -4468 sw
tri 35917 -4470 35919 -4468 ne
rect 35919 -4470 35964 -4468
tri 35964 -4470 35993 -4441 sw
tri 36107 -4470 36136 -4441 ne
rect 36136 -4470 36181 -4441
tri 36181 -4470 36210 -4441 sw
rect 35865 -4482 35867 -4470
tri 35867 -4482 35879 -4470 sw
tri 35919 -4482 35931 -4470 ne
rect 35931 -4482 35993 -4470
rect 35865 -4515 35879 -4482
tri 35879 -4515 35912 -4482 sw
tri 35931 -4515 35964 -4482 ne
rect 35964 -4515 35993 -4482
tri 35993 -4515 36038 -4470 sw
tri 36136 -4503 36169 -4470 ne
rect 36169 -4503 36210 -4470
tri 36210 -4503 36243 -4470 sw
tri 36169 -4515 36181 -4503 ne
rect 36181 -4515 36243 -4503
tri 36243 -4515 36255 -4503 sw
rect 35865 -4534 35912 -4515
tri 35912 -4534 35931 -4515 sw
tri 35964 -4534 35983 -4515 ne
rect 35983 -4534 36038 -4515
tri 35865 -4565 35896 -4534 ne
rect 35896 -4548 35931 -4534
tri 35931 -4548 35945 -4534 sw
tri 35983 -4548 35997 -4534 ne
rect 35997 -4548 36038 -4534
rect 35896 -4565 35945 -4548
tri 35945 -4565 35962 -4548 sw
tri 35997 -4565 36014 -4548 ne
rect 36014 -4565 36038 -4548
tri 35896 -4600 35931 -4565 ne
rect 35931 -4589 35962 -4565
tri 35962 -4589 35986 -4565 sw
tri 36014 -4589 36038 -4565 ne
tri 36038 -4589 36112 -4515 sw
tri 36181 -4577 36243 -4515 ne
rect 36243 -4577 36255 -4515
tri 36255 -4577 36317 -4515 sw
tri 36243 -4589 36255 -4577 ne
rect 36255 -4589 36317 -4577
tri 36317 -4589 36329 -4577 sw
rect 35931 -4600 35986 -4589
tri 35986 -4600 35997 -4589 sw
tri 36038 -4600 36049 -4589 ne
rect 36049 -4600 36112 -4589
tri 35931 -4666 35997 -4600 ne
tri 35997 -4614 36011 -4600 sw
tri 36049 -4614 36063 -4600 ne
rect 36063 -4614 36112 -4600
rect 35997 -4663 36011 -4614
tri 36011 -4663 36060 -4614 sw
tri 36063 -4663 36112 -4614 ne
tri 36112 -4663 36186 -4589 sw
tri 36255 -4651 36317 -4589 ne
rect 36317 -4651 36329 -4589
tri 36329 -4651 36391 -4589 sw
rect 39702 -4619 39812 -4573
tri 36317 -4663 36329 -4651 ne
rect 36329 -4663 36391 -4651
tri 36391 -4663 36403 -4651 sw
rect 35997 -4666 36060 -4663
tri 36060 -4666 36063 -4663 sw
tri 35997 -4686 36017 -4666 ne
tri 36012 -4843 36017 -4838 se
rect 36017 -4843 36063 -4666
tri 36112 -4737 36186 -4663 ne
tri 36186 -4737 36260 -4663 sw
tri 36329 -4725 36391 -4663 ne
rect 36391 -4725 36403 -4663
tri 36403 -4725 36465 -4663 sw
tri 36391 -4737 36403 -4725 ne
rect 36403 -4737 36515 -4725
tri 36186 -4811 36260 -4737 ne
tri 36260 -4811 36334 -4737 sw
tri 36403 -4777 36443 -4737 ne
rect 36443 -4777 36515 -4737
tri 36260 -4843 36292 -4811 ne
rect 36292 -4843 36334 -4811
tri 35999 -4856 36012 -4843 se
rect 36012 -4856 36063 -4843
tri 36063 -4856 36076 -4843 sw
tri 36292 -4856 36305 -4843 ne
rect 36305 -4856 36334 -4843
tri 35983 -4872 35999 -4856 se
rect 35999 -4872 36076 -4856
tri 36076 -4872 36092 -4856 sw
rect 35964 -4924 35970 -4872
rect 36022 -4924 36034 -4872
rect 36086 -4924 36092 -4872
tri 36305 -4885 36334 -4856 ne
tri 36334 -4885 36408 -4811 sw
tri 36334 -4887 36336 -4885 ne
rect 36336 -4887 36526 -4885
tri 36336 -4900 36349 -4887 ne
rect 36349 -4900 36526 -4887
tri 36349 -4924 36373 -4900 ne
rect 36373 -4924 36526 -4900
tri 36373 -4937 36386 -4924 ne
rect 36386 -4937 36526 -4924
rect 35425 -5092 35439 -5060
tri 35439 -5092 35471 -5060 nw
tri 33494 -5138 33540 -5092 ne
rect 33540 -5138 35393 -5092
tri 35393 -5138 35439 -5092 nw
tri 32777 -5170 32792 -5155 se
rect 32792 -5170 32799 -5155
tri 32524 -5222 32576 -5170 se
rect 32576 -5222 32799 -5170
tri 32799 -5222 32866 -5155 nw
tri 32119 -5252 32147 -5224 ne
rect 31305 -6025 31311 -5973
rect 31363 -6025 31375 -5973
rect 31427 -6025 31433 -5973
rect 26384 -6062 26386 -6059
rect 26438 -6062 26440 -6059
rect 26384 -6068 26440 -6062
rect 30727 -6081 30733 -6029
rect 30785 -6081 30797 -6029
rect 30849 -6081 30855 -6029
rect 32147 -6268 32213 -5224
tri 32504 -5242 32524 -5222 se
rect 32524 -5230 32590 -5222
tri 32590 -5230 32598 -5222 nw
rect 32524 -5242 32559 -5230
rect 32504 -5261 32559 -5242
tri 32559 -5261 32590 -5230 nw
tri 33316 -5261 33347 -5230 sw
rect 39766 -5259 39812 -4619
tri 33634 -5261 33636 -5259 se
rect 33636 -5261 39812 -5259
rect 32244 -5402 32250 -5350
rect 32302 -5402 32314 -5350
rect 32366 -5402 32372 -5350
tri 32265 -5423 32286 -5402 ne
rect 32286 -5423 32351 -5402
tri 32351 -5423 32372 -5402 nw
tri 32286 -5436 32299 -5423 ne
rect 32299 -5827 32351 -5423
rect 32504 -5695 32556 -5261
tri 32556 -5264 32559 -5261 nw
tri 33263 -5262 33264 -5261 se
rect 33263 -5264 33264 -5262
rect 33316 -5264 33347 -5261
tri 33347 -5264 33350 -5261 sw
tri 33631 -5264 33634 -5261 se
rect 33634 -5264 39812 -5261
tri 33621 -5274 33631 -5264 se
rect 33631 -5274 39812 -5264
rect 32991 -5280 33043 -5274
tri 33603 -5292 33621 -5274 se
rect 33621 -5292 39812 -5274
rect 32991 -5344 33043 -5332
tri 33111 -5346 33165 -5292 se
tri 33573 -5322 33603 -5292 se
rect 33603 -5305 39812 -5292
rect 33603 -5322 33636 -5305
tri 33215 -5346 33239 -5322 sw
tri 33570 -5325 33573 -5322 se
rect 33573 -5325 33636 -5322
tri 33636 -5325 33656 -5305 nw
tri 33549 -5346 33570 -5325 se
tri 33504 -5391 33549 -5346 se
rect 33549 -5391 33570 -5346
tri 33570 -5391 33636 -5325 nw
rect 32991 -5402 33043 -5396
tri 33495 -5400 33504 -5391 se
rect 33504 -5400 33527 -5391
tri 33043 -5402 33045 -5400 sw
tri 33493 -5402 33495 -5400 se
rect 33495 -5402 33527 -5400
rect 32991 -5423 33045 -5402
tri 33045 -5423 33066 -5402 sw
tri 33472 -5423 33493 -5402 se
rect 33493 -5423 33527 -5402
rect 32991 -5434 33066 -5423
tri 33066 -5434 33077 -5423 sw
tri 33461 -5434 33472 -5423 se
rect 33472 -5434 33527 -5423
tri 33527 -5434 33570 -5391 nw
rect 32991 -5460 33501 -5434
tri 33501 -5460 33527 -5434 nw
tri 32991 -5469 33000 -5460 ne
rect 33000 -5469 33492 -5460
tri 33492 -5469 33501 -5460 nw
tri 32956 -5507 32990 -5473 sw
tri 32504 -5738 32547 -5695 ne
rect 32547 -5738 32556 -5695
tri 32556 -5738 32621 -5673 sw
tri 32547 -5747 32556 -5738 ne
rect 32556 -5747 32621 -5738
tri 32556 -5812 32621 -5747 ne
tri 32621 -5812 32695 -5738 sw
tri 32621 -5823 32632 -5812 ne
rect 32632 -5823 32695 -5812
rect 32299 -5891 32351 -5879
rect 32299 -5949 32351 -5943
rect 32394 -5959 32403 -5823
rect 32539 -5829 32548 -5823
rect 32540 -5881 32548 -5829
tri 32632 -5834 32643 -5823 ne
rect 32539 -5895 32548 -5881
rect 32540 -5947 32548 -5895
rect 32539 -5959 32548 -5947
rect 32643 -6099 32695 -5823
tri 34800 -5876 34824 -5852 sw
rect 38121 -5902 38173 -5896
rect 38121 -5966 38173 -5954
rect 33157 -5984 33236 -5981
tri 33236 -5984 33239 -5981 sw
rect 33157 -5987 33239 -5984
rect 33209 -5988 33239 -5987
tri 33239 -5988 33243 -5984 sw
tri 33671 -5988 33675 -5984 sw
rect 33209 -6018 33243 -5988
tri 33243 -6018 33273 -5988 sw
tri 33589 -6018 33619 -5988 se
rect 33671 -6018 33675 -5988
tri 33675 -6018 33705 -5988 sw
rect 37956 -6018 38121 -5972
rect 33209 -6019 33273 -6018
tri 33273 -6019 33274 -6018 sw
rect 33209 -6024 33274 -6019
tri 33274 -6024 33279 -6019 sw
rect 37956 -6024 38173 -6018
rect 38207 -6019 38259 -6013
rect 33209 -6039 33279 -6024
rect 33157 -6042 33279 -6039
tri 33279 -6042 33297 -6024 sw
rect 33157 -6049 33297 -6042
tri 33297 -6049 33304 -6042 sw
rect 33157 -6051 33304 -6049
rect 33209 -6053 33304 -6051
tri 33304 -6053 33308 -6049 sw
tri 37354 -6053 37358 -6049 ne
rect 33209 -6071 33308 -6053
tri 33308 -6071 33326 -6053 sw
rect 33209 -6073 33326 -6071
tri 33326 -6073 33328 -6071 sw
rect 33209 -6083 33328 -6073
tri 33328 -6083 33338 -6073 sw
rect 33209 -6103 33338 -6083
rect 33157 -6109 33338 -6103
tri 33290 -6135 33316 -6109 ne
rect 33316 -6135 33338 -6109
tri 33338 -6135 33390 -6083 sw
rect 37668 -6089 37720 -6042
tri 38191 -6071 38207 -6055 se
tri 38179 -6083 38191 -6071 se
rect 38191 -6083 38259 -6071
tri 38173 -6089 38179 -6083 se
rect 38179 -6089 38207 -6083
rect 37668 -6135 38207 -6089
tri 33316 -6147 33328 -6135 ne
rect 33328 -6141 33390 -6135
tri 33390 -6141 33396 -6135 sw
rect 37668 -6141 38259 -6135
rect 33328 -6147 33396 -6141
tri 33396 -6147 33402 -6141 sw
rect 32643 -6163 32695 -6151
rect 32643 -6221 32695 -6215
tri 33328 -6221 33402 -6147 ne
tri 33402 -6221 33476 -6147 sw
tri 33402 -6264 33445 -6221 ne
rect 33445 -6230 35113 -6221
rect 33445 -6264 35057 -6230
tri 35023 -6267 35026 -6264 ne
rect 35026 -6267 35057 -6264
tri 32213 -6268 32214 -6267 sw
tri 35026 -6268 35027 -6267 ne
rect 35027 -6268 35057 -6267
rect 32147 -6295 32214 -6268
tri 32147 -6298 32150 -6295 ne
rect 32150 -6298 32214 -6295
tri 32214 -6298 32244 -6268 sw
tri 32697 -6298 32727 -6268 se
rect 32727 -6277 32783 -6268
tri 32150 -6361 32213 -6298 ne
rect 32213 -6333 32727 -6298
tri 35027 -6298 35057 -6268 ne
rect 32213 -6357 32783 -6333
rect 32213 -6361 32727 -6357
tri 32213 -6364 32216 -6361 ne
rect 32216 -6364 32727 -6361
tri 32697 -6394 32727 -6364 ne
rect 35057 -6310 35113 -6286
rect 35057 -6375 35113 -6366
rect 32727 -6422 32783 -6413
tri 26259 -6801 26293 -6767 se
tri 26321 -6801 26355 -6767 sw
tri 41412 -8324 41444 -8292 se
tri 41195 -8404 41229 -8370 nw
tri 41410 -8404 41444 -8370 ne
<< via2 >>
rect 33819 -143 33875 -87
rect 33819 -223 33875 -167
rect 26324 -4242 26328 -4193
rect 26328 -4242 26380 -4193
rect 26324 -4249 26380 -4242
rect 26324 -4308 26328 -4273
rect 26328 -4308 26380 -4273
rect 26324 -4329 26380 -4308
rect 26384 -5946 26440 -5923
rect 26384 -5979 26386 -5946
rect 26386 -5979 26438 -5946
rect 26438 -5979 26440 -5946
rect 26384 -6010 26440 -6003
rect 26384 -6059 26386 -6010
rect 26386 -6059 26438 -6010
rect 26438 -6059 26440 -6010
rect 33819 -2179 33875 -2123
rect 33819 -2259 33875 -2203
rect 34658 -3637 34714 -3581
rect 34658 -3717 34714 -3661
rect 35057 -4585 35113 -4574
rect 35057 -4630 35109 -4585
rect 35109 -4630 35113 -4585
rect 35057 -4701 35109 -4654
rect 35109 -4701 35113 -4654
rect 35057 -4710 35113 -4701
rect 32403 -5829 32539 -5823
rect 32403 -5881 32416 -5829
rect 32416 -5881 32468 -5829
rect 32468 -5881 32488 -5829
rect 32488 -5881 32539 -5829
rect 32403 -5895 32539 -5881
rect 32403 -5947 32416 -5895
rect 32416 -5947 32468 -5895
rect 32468 -5947 32488 -5895
rect 32488 -5947 32539 -5895
rect 32403 -5959 32539 -5947
rect 32727 -6333 32783 -6277
rect 35057 -6286 35113 -6230
rect 32727 -6413 32783 -6357
rect 35057 -6366 35113 -6310
<< metal3 >>
rect 33814 -87 33880 -82
rect 33814 -143 33819 -87
rect 33875 -143 33880 -87
rect 33814 -167 33880 -143
rect 33814 -223 33819 -167
rect 33875 -223 33880 -167
rect 27216 -1234 27255 -1209
rect 33814 -2123 33880 -223
rect 33814 -2179 33819 -2123
rect 33875 -2179 33880 -2123
rect 33814 -2203 33880 -2179
rect 33814 -2259 33819 -2203
rect 33875 -2259 33880 -2203
rect 33814 -2264 33880 -2259
rect 34653 -3581 34719 -3576
rect 34653 -3637 34658 -3581
rect 34714 -3637 34719 -3581
rect 34653 -3661 34719 -3637
tri 34629 -3717 34653 -3693 se
rect 34653 -3717 34658 -3661
rect 34714 -3717 34719 -3661
tri 34559 -3787 34629 -3717 se
rect 34629 -3722 34719 -3717
rect 34629 -3787 34653 -3722
tri 34653 -3787 34718 -3722 nw
tri 34467 -3879 34559 -3787 se
rect 34559 -3879 34561 -3787
tri 34561 -3879 34653 -3787 nw
rect 26319 -4193 26385 -4188
rect 26319 -4249 26324 -4193
rect 26380 -4249 26385 -4193
rect 26319 -4273 26385 -4249
rect 26319 -4329 26324 -4273
rect 26380 -4329 26385 -4273
rect 26319 -4654 26385 -4329
tri 26385 -4654 26402 -4637 sw
rect 26319 -4665 26402 -4654
tri 26402 -4665 26413 -4654 sw
tri 26319 -4710 26364 -4665 ne
rect 26364 -4697 26413 -4665
tri 26413 -4697 26445 -4665 sw
rect 26364 -4710 26445 -4697
tri 26364 -4725 26379 -4710 ne
rect 26379 -5923 26445 -4710
rect 26379 -5979 26384 -5923
rect 26440 -5979 26445 -5923
rect 32398 -5823 32544 -5818
rect 32398 -5959 32403 -5823
rect 32539 -5959 32544 -5823
rect 32398 -5964 32544 -5959
rect 26379 -6003 26445 -5979
rect 26379 -6059 26384 -6003
rect 26440 -6059 26445 -6003
rect 26379 -6064 26445 -6059
rect 32722 -6277 32788 -6270
rect 32722 -6333 32727 -6277
rect 32783 -6333 32788 -6277
rect 32722 -6357 32788 -6333
rect 32722 -6413 32727 -6357
rect 32783 -6413 32788 -6357
rect 32722 -8303 32788 -6413
tri 34373 -7363 34467 -7269 se
rect 34467 -7297 34533 -3879
tri 34533 -3907 34561 -3879 nw
rect 35052 -4574 35118 -4569
rect 35052 -4630 35057 -4574
rect 35113 -4630 35118 -4574
rect 35052 -4654 35118 -4630
rect 35052 -4710 35057 -4654
rect 35113 -4710 35118 -4654
rect 35052 -6230 35118 -4710
rect 35052 -6286 35057 -6230
rect 35113 -6286 35118 -6230
rect 35052 -6310 35118 -6286
rect 35052 -6366 35057 -6310
rect 35113 -6366 35118 -6310
rect 35052 -6371 35118 -6366
tri 34467 -7363 34533 -7297 nw
tri 34279 -7457 34373 -7363 se
tri 34373 -7457 34467 -7363 nw
tri 34185 -7551 34279 -7457 se
tri 34279 -7551 34373 -7457 nw
tri 34091 -7645 34185 -7551 se
tri 34185 -7645 34279 -7551 nw
tri 33997 -7739 34091 -7645 se
tri 34091 -7739 34185 -7645 nw
tri 33903 -7833 33997 -7739 se
tri 33997 -7833 34091 -7739 nw
tri 33809 -7927 33903 -7833 se
tri 33903 -7927 33997 -7833 nw
tri 33715 -8021 33809 -7927 se
tri 33809 -8021 33903 -7927 nw
tri 33621 -8115 33715 -8021 se
tri 33715 -8115 33809 -8021 nw
tri 33527 -8209 33621 -8115 se
tri 33621 -8209 33715 -8115 nw
tri 33435 -8301 33527 -8209 se
tri 32788 -8303 32790 -8301 sw
tri 33433 -8303 33435 -8301 se
rect 33435 -8303 33527 -8301
tri 33527 -8303 33621 -8209 nw
rect 32722 -8329 32790 -8303
tri 32722 -8382 32775 -8329 ne
rect 32775 -8382 32790 -8329
tri 32790 -8382 32869 -8303 sw
tri 33354 -8382 33433 -8303 se
rect 33433 -8382 33448 -8303
tri 33448 -8382 33527 -8303 nw
tri 32775 -8395 32788 -8382 ne
rect 32788 -8395 33435 -8382
tri 33435 -8395 33448 -8382 nw
tri 32788 -8448 32841 -8395 ne
rect 32841 -8448 33382 -8395
tri 33382 -8448 33435 -8395 nw
use sky130_fd_io__gpiov2_amux_ls  sky130_fd_io__gpiov2_amux_ls_0
timestamp 1619729480
transform 1 0 25054 0 1 -16031
box 920 -428 17006 17121
use sky130_fd_io__gpiov2_amux_decoder  sky130_fd_io__gpiov2_amux_decoder_0
timestamp 1619729480
transform 1 0 31774 0 1 -5388
box -369 -792 8677 3339
use sky130_fd_io__gpiov2_amux_drvr  sky130_fd_io__gpiov2_amux_drvr_0
timestamp 1619729480
transform 1 0 9862 0 1 6253
box 15993 -15244 28326 -4277
<< labels >>
flabel comment s 33085 -3513 33085 -3513 0 FreeSans 440 90 0 0 LV_NET
flabel metal1 s 33752 -3713 33780 -3685 3 FreeSans 520 0 0 0 ANALOG_EN
flabel metal1 s 33086 -4668 33114 -4640 3 FreeSans 520 0 0 0 NMIDA_VCCD
flabel metal1 s 32531 -4885 32559 -4857 3 FreeSans 520 0 0 0 D_B
flabel metal1 s 28136 -4088 28164 -4060 3 FreeSans 520 0 0 0 PD_CSD_VSWITCH_H
flabel metal1 s 28983 -3582 29011 -3554 3 FreeSans 520 0 0 0 NGB_AMX_VSWITCH_H
flabel metal1 s 28637 -3170 28665 -3142 3 FreeSans 520 0 0 0 NGA_AMX_VSWITCH_H
flabel metal1 s 35982 -4887 36010 -4859 3 FreeSans 520 0 0 0 NGB_PAD_VSWITCH_H
flabel metal1 s 35326 -4887 35354 -4859 3 FreeSans 520 0 0 0 NGA_PAD_VSWITCH_H
flabel metal1 s 34851 -4893 34879 -4865 3 FreeSans 520 0 0 0 PGB_AMX_VDDA_H_N
flabel metal1 s 34402 -4670 34430 -4642 3 FreeSans 520 0 0 0 PGA_AMX_VDDA_H_N
flabel metal1 s 35044 -4676 35072 -4648 3 FreeSans 520 0 0 0 PGB_PAD_VDDIOQ_H_N
flabel metal1 s 34567 -4571 34595 -4543 3 FreeSans 520 0 0 0 PGA_PAD_VDDIOQ_H_N
flabel metal1 s 36703 -2411 36731 -2383 3 FreeSans 520 0 0 0 PU_CSD_VDDIOQ_H_N
flabel metal1 s 35760 -3734 35788 -3706 3 FreeSans 520 0 0 0 OUT
flabel metal1 s 32208 -3047 32236 -3019 3 FreeSans 520 0 0 0 ANALOG_SEL
flabel metal1 s 35760 -3047 35788 -3019 3 FreeSans 520 0 0 0 ANALOG_POL
flabel metal1 s 26770 -869 26798 -841 3 FreeSans 520 0 0 0 VSSA
flabel metal1 s 40633 -14280 40661 -14252 3 FreeSans 520 180 0 0 HLD_I_H_N
flabel metal1 s 41427 -14232 41455 -14204 3 FreeSans 520 0 0 0 HLD_I_H
flabel metal1 s 29152 -4932 29180 -4904 3 FreeSans 520 0 0 0 ENABLE_VSWITCH_H
flabel metal1 s 27432 -1093 27460 -1065 3 FreeSans 520 0 0 0 ENABLE_VDDA_H
flabel metal1 s 40244 -15218 40272 -15190 3 FreeSans 520 0 0 0 ANALOG_EN
flabel metal1 s 27142 -1090 27170 -1062 3 FreeSans 520 0 0 0 AMUX_EN_VDDIO_H_N
flabel metal1 s 26514 -819 26542 -791 3 FreeSans 520 0 0 0 AMUX_EN_VDDA_H_N
flabel metal1 s 40195 -14876 40223 -14848 3 FreeSans 520 0 0 0 VCCD
flabel metal1 s 26743 885 26771 913 3 FreeSans 520 0 0 0 VDDA
flabel metal1 s 40211 -13346 40239 -13318 3 FreeSans 520 180 0 0 VDDIO_Q
flabel metal1 s 27319 -4493 27347 -4465 3 FreeSans 520 0 0 0 VSWITCH
flabel metal1 s 40188 -15545 40216 -15517 3 FreeSans 520 0 0 0 VSSD
flabel metal1 s 36491 -6038 36519 -6010 3 FreeSans 520 0 0 0 VCCD
flabel metal1 s 32768 -4293 32796 -4265 3 FreeSans 520 0 0 0 VCCD
flabel metal1 s 28020 -2548 28048 -2520 3 FreeSans 520 0 0 0 VCCD
flabel metal1 s 27621 -6954 27649 -6926 3 FreeSans 520 0 0 0 VCCD
flabel metal1 s 26296 1600 26324 1628 3 FreeSans 520 0 0 0 VDDA
flabel metal1 s 36626 -5468 36654 -5440 3 FreeSans 520 0 0 0 VDDIO_Q
flabel metal1 s 32863 -5897 32891 -5869 3 FreeSans 520 0 0 0 VDDIO_Q
flabel metal1 s 27079 -6424 27107 -6396 3 FreeSans 520 0 0 0 VDDIO_Q
flabel metal1 s 28787 -3182 28815 -3154 3 FreeSans 520 0 0 0 VSSA
flabel metal1 s 28787 -1747 28815 -1719 3 FreeSans 520 0 0 0 VSSA
flabel metal1 s 28363 -819 28391 -791 3 FreeSans 520 0 0 0 VSSA
flabel metal1 s 38044 -6278 38072 -6250 3 FreeSans 520 0 0 0 VSSD
flabel metal1 s 32823 -5096 32851 -5068 3 FreeSans 520 0 0 0 VSSD
flabel metal1 s 26922 -7260 26950 -7232 3 FreeSans 520 0 0 0 VSSD
flabel metal1 s 28361 -4216 28389 -4188 3 FreeSans 520 0 0 0 VSWITCH
flabel metal1 s 27326 -3826 27354 -3798 3 FreeSans 520 0 0 0 VSWITCH
flabel metal1 s 40209 -14862 40209 -14862 3 FreeSans 280 180 0 0 VCCD
flabel metal1 s 41358 -13673 41386 -13645 3 FreeSans 280 0 0 0 VCCD
flabel metal1 s 26757 899 26757 899 3 FreeSans 520 0 0 0 VDDA
flabel metal1 s 40225 -13332 40225 -13332 3 FreeSans 520 180 0 0 VDDIO_Q
flabel metal1 s 26784 -855 26784 -855 3 FreeSans 520 0 0 0 VSSA
flabel metal1 s 27468 -1736 27496 -1708 3 FreeSans 520 0 0 0 VSSA
flabel metal1 s 28938 -4558 28966 -4530 3 FreeSans 520 0 0 0 VSSA
flabel metal1 s 26773 -4692 26801 -4664 3 FreeSans 520 0 0 0 VSSA
flabel metal1 s 26230 -818 26258 -790 3 FreeSans 520 0 0 0 VSSA
flabel metal1 s 40202 -15531 40202 -15531 3 FreeSans 280 180 0 0 VSSD
flabel metal1 s 41023 -14572 41051 -14544 3 FreeSans 280 0 0 0 VSSD
flabel metal1 s 27333 -4479 27333 -4479 3 FreeSans 520 0 0 0 VSWITCH
flabel metal1 s 26442 -5168 26470 -5140 3 FreeSans 520 0 0 0 VSWITCH
flabel metal1 s 35376 -3355 35404 -3327 3 FreeSans 280 0 0 0 VCCD
flabel metal1 s 37007 -4065 37035 -4037 3 FreeSans 280 0 0 0 VCCD
flabel metal1 s 35238 -4290 35266 -4262 3 FreeSans 280 0 0 0 VCCD
flabel metal1 s 35376 -2739 35404 -2711 3 FreeSans 280 0 0 0 VSSD
flabel metal1 s 35376 -4018 35404 -3990 3 FreeSans 280 0 0 0 VSSD
flabel metal1 s 35269 -5113 35297 -5085 3 FreeSans 280 0 0 0 VSSD
flabel metal1 s 37380 -2821 37408 -2793 3 FreeSans 280 0 0 0 VSSD
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 18855940
string GDS_START 18786756
<< end >>
