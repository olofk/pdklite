magic
tech sky130A
timestamp 1640697675
<< properties >>
string gencell sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_lishield
string parameter m=1
string library sky130
<< end >>
