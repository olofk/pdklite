magic
tech sky130A
magscale 1 2
timestamp 1640697980
<< nwell >>
rect -38 261 2706 582
<< pwell >>
rect 3 21 273 203
rect 293 21 735 203
rect 757 21 1195 203
rect 1473 21 1911 203
rect 1933 21 2375 203
rect 2395 21 2665 203
rect 29 -17 63 17
rect 213 -17 247 21
rect 672 -17 706 21
rect 1132 -17 1166 21
rect 1225 -17 1259 17
rect 1502 -17 1536 21
rect 1962 -17 1996 21
rect 2421 -17 2455 21
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 29 299 71 527
rect 205 299 251 527
rect 29 17 71 181
rect 563 367 629 527
rect 774 367 825 527
rect 959 367 993 527
rect 1127 299 1179 527
rect 1251 382 1317 527
rect 843 255 993 265
rect 843 221 955 255
rect 989 221 993 255
rect 843 215 993 221
rect 1027 255 1179 265
rect 1027 221 1141 255
rect 1175 221 1179 255
rect 1027 215 1179 221
rect 205 17 251 181
rect 303 17 361 111
rect 495 17 529 111
rect 663 17 718 181
rect 1043 17 1077 109
rect 1351 255 1455 493
rect 1489 299 1541 527
rect 1675 367 1709 527
rect 1843 367 1894 527
rect 2039 367 2105 527
rect 1351 221 1353 255
rect 1387 221 1455 255
rect 1351 183 1455 221
rect 1489 255 1641 265
rect 1489 221 1525 255
rect 1559 221 1641 255
rect 1489 215 1641 221
rect 1675 255 1825 265
rect 1675 221 1697 255
rect 1731 221 1825 255
rect 1675 215 1825 221
rect 2417 299 2463 527
rect 2597 299 2639 527
rect 1351 17 1419 149
rect 1591 17 1625 109
rect 1950 17 2005 181
rect 2139 17 2173 111
rect 2307 17 2365 111
rect 2417 17 2463 181
rect 2597 17 2639 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 955 221 989 255
rect 1141 221 1175 255
rect 1353 221 1387 255
rect 1525 221 1559 255
rect 1697 221 1731 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
<< obsli1 >>
rect 105 297 171 493
rect 301 459 529 493
rect 301 367 361 459
rect 395 333 461 425
rect 105 177 155 297
rect 309 289 461 333
rect 495 333 529 459
rect 663 333 718 493
rect 859 333 925 493
rect 1027 333 1093 493
rect 495 291 718 333
rect 753 299 1093 333
rect 189 215 255 265
rect 309 181 352 289
rect 386 215 540 255
rect 574 215 718 255
rect 753 181 809 299
rect 105 51 171 177
rect 309 147 629 181
rect 395 145 629 147
rect 395 51 461 145
rect 563 51 629 145
rect 753 131 925 181
rect 959 143 1179 177
rect 775 93 841 97
rect 959 93 1009 143
rect 775 51 1009 93
rect 1111 51 1179 143
rect 1213 51 1317 348
rect 1575 333 1641 493
rect 1743 333 1809 493
rect 1950 333 2005 493
rect 2139 459 2367 493
rect 2139 333 2173 459
rect 1575 299 1915 333
rect 1859 181 1915 299
rect 1950 291 2173 333
rect 2207 333 2273 425
rect 2307 367 2367 459
rect 2207 289 2359 333
rect 2497 297 2563 493
rect 1950 215 2094 255
rect 2128 215 2282 255
rect 2316 181 2359 289
rect 2413 215 2479 265
rect 1489 143 1709 177
rect 1489 51 1557 143
rect 1659 93 1709 143
rect 1743 131 1915 181
rect 1827 93 1893 97
rect 1659 51 1893 93
rect 2039 147 2359 181
rect 2039 145 2273 147
rect 2039 51 2105 145
rect 2207 51 2273 145
rect 2513 177 2563 297
rect 2497 51 2563 177
<< metal1 >>
rect 0 561 2668 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 0 496 2668 527
rect 943 255 1001 261
rect 943 221 955 255
rect 989 252 1001 255
rect 1129 255 1187 261
rect 1129 252 1141 255
rect 989 224 1141 252
rect 989 221 1001 224
rect 943 215 1001 221
rect 1129 221 1141 224
rect 1175 252 1187 255
rect 1341 255 1399 261
rect 1341 252 1353 255
rect 1175 224 1353 252
rect 1175 221 1187 224
rect 1129 215 1187 221
rect 1341 221 1353 224
rect 1387 252 1399 255
rect 1513 255 1571 261
rect 1513 252 1525 255
rect 1387 224 1525 252
rect 1387 221 1399 224
rect 1341 215 1399 221
rect 1513 221 1525 224
rect 1559 252 1571 255
rect 1685 255 1743 261
rect 1685 252 1697 255
rect 1559 224 1697 252
rect 1559 221 1571 224
rect 1513 215 1571 221
rect 1685 221 1697 224
rect 1731 221 1743 255
rect 1685 215 1743 221
rect 0 17 2668 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
rect 0 -48 2668 -17
<< obsm1 >>
rect 101 215 175 261
rect 205 252 263 261
rect 302 252 360 261
rect 205 224 360 252
rect 205 215 263 224
rect 302 215 360 224
rect 408 252 466 261
rect 580 252 638 261
rect 752 252 810 261
rect 408 224 810 252
rect 408 215 466 224
rect 580 215 638 224
rect 752 215 810 224
rect 1857 252 1915 261
rect 2029 252 2087 261
rect 2201 252 2259 261
rect 1857 224 2259 252
rect 1857 215 1915 224
rect 2029 215 2087 224
rect 2201 215 2259 224
rect 2309 252 2367 261
rect 2406 252 2464 261
rect 2309 224 2464 252
rect 2309 215 2367 224
rect 2406 215 2464 224
rect 2494 215 2567 261
<< labels >>
rlabel metal1 s 0 -48 2668 48 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 2605 -17 2639 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 2513 -17 2547 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 2421 -17 2455 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 2329 -17 2363 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 2237 -17 2271 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 2145 -17 2179 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 2053 -17 2087 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 1961 -17 1995 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 1869 -17 1903 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 1777 -17 1811 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 1685 -17 1719 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 1593 -17 1627 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 1501 -17 1535 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 1409 -17 1443 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 1317 -17 1351 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 1225 -17 1259 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 1133 -17 1167 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 1041 -17 1075 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 949 -17 983 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 857 -17 891 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 765 -17 799 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 673 -17 707 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 581 -17 615 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 489 -17 523 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 397 -17 431 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 305 -17 339 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 213 -17 247 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 121 -17 155 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 29 -17 63 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 0 -17 2668 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 2597 17 2639 181 6 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 2417 17 2463 181 6 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 2307 17 2365 111 6 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 2139 17 2173 111 6 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 1950 17 2005 181 6 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 1591 17 1625 109 6 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 1351 17 1419 149 6 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 1043 17 1077 109 6 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 663 17 718 181 6 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 495 17 529 111 6 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 303 17 361 111 6 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 205 17 251 181 6 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 29 17 71 181 6 VGND
port 1 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 2 nsew ground bidirectional
rlabel nwell s -38 261 2706 582 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 0 496 2668 592 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 2605 527 2639 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 2513 527 2547 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 2421 527 2455 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 2329 527 2363 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 2237 527 2271 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 2145 527 2179 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 2053 527 2087 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 1961 527 1995 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 1869 527 1903 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 1777 527 1811 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 1685 527 1719 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 1593 527 1627 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 1501 527 1535 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 1409 527 1443 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 1317 527 1351 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 1225 527 1259 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 1133 527 1167 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 1041 527 1075 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 949 527 983 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 857 527 891 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 765 527 799 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 673 527 707 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 581 527 615 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 489 527 523 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 397 527 431 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 305 527 339 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 213 527 247 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 121 527 155 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 29 527 63 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 2597 299 2639 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 2417 299 2463 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 2039 367 2105 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1843 367 1894 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1675 367 1709 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1489 299 1541 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1251 382 1317 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 1127 299 1179 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 959 367 993 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 774 367 825 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 563 367 629 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 205 299 251 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 29 299 71 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 2668 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 1685 215 1743 224 6 LO
port 5 nsew signal output
rlabel metal1 s 1513 215 1571 224 6 LO
port 5 nsew signal output
rlabel metal1 s 1341 215 1399 224 6 LO
port 5 nsew signal output
rlabel metal1 s 1129 215 1187 224 6 LO
port 5 nsew signal output
rlabel metal1 s 943 215 1001 224 6 LO
port 5 nsew signal output
rlabel metal1 s 943 224 1743 252 6 LO
port 5 nsew signal output
rlabel metal1 s 1685 252 1743 261 6 LO
port 5 nsew signal output
rlabel metal1 s 1513 252 1571 261 6 LO
port 5 nsew signal output
rlabel metal1 s 1341 252 1399 261 6 LO
port 5 nsew signal output
rlabel metal1 s 1129 252 1187 261 6 LO
port 5 nsew signal output
rlabel metal1 s 943 252 1001 261 6 LO
port 5 nsew signal output
rlabel viali s 1697 221 1731 255 6 LO
port 5 nsew signal output
rlabel locali s 1675 215 1825 265 6 LO
port 5 nsew signal output
rlabel viali s 1525 221 1559 255 6 LO
port 5 nsew signal output
rlabel locali s 1489 215 1641 265 6 LO
port 5 nsew signal output
rlabel viali s 1353 221 1387 255 6 LO
port 5 nsew signal output
rlabel locali s 1351 183 1455 493 6 LO
port 5 nsew signal output
rlabel viali s 1141 221 1175 255 6 LO
port 5 nsew signal output
rlabel locali s 1027 215 1179 265 6 LO
port 5 nsew signal output
rlabel viali s 955 221 989 255 6 LO
port 5 nsew signal output
rlabel locali s 843 215 993 265 6 LO
port 5 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2668 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1656842
string GDS_START 1652916
<< end >>
