magic
tech sky130A
magscale 1 2
timestamp 1640697980
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1168 157 1350 201
rect 1653 157 1930 203
rect 1 145 821 157
rect 1022 145 1930 157
rect 1 21 1930 145
rect 29 -17 63 21
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 104 427 170 527
rect 19 195 89 325
rect 103 17 169 93
rect 376 449 442 527
rect 352 167 386 337
rect 492 271 558 337
rect 746 433 785 527
rect 352 157 398 167
rect 613 157 650 219
rect 706 211 798 331
rect 352 127 650 157
rect 374 123 650 127
rect 1180 367 1214 527
rect 392 17 461 89
rect 495 61 530 123
rect 752 17 792 109
rect 1558 427 1619 527
rect 1775 325 1809 527
rect 1138 17 1212 117
rect 1846 301 1915 479
rect 1543 17 1617 123
rect 1881 164 1915 301
rect 1775 17 1809 139
rect 1846 61 1915 164
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< obsli1 >>
rect 36 393 70 493
rect 36 359 169 393
rect 123 194 169 359
rect 123 161 162 194
rect 35 127 162 161
rect 204 143 246 493
rect 35 69 69 127
rect 203 69 246 143
rect 284 415 342 489
rect 538 449 712 483
rect 284 372 644 415
rect 284 93 318 372
rect 423 226 458 372
rect 610 327 644 372
rect 678 399 712 449
rect 836 413 884 488
rect 932 438 1146 472
rect 836 399 870 413
rect 678 365 870 399
rect 610 261 654 327
rect 423 192 492 226
rect 836 177 870 365
rect 684 143 870 177
rect 904 207 952 381
rect 990 331 1078 402
rect 1112 315 1146 438
rect 1248 427 1298 493
rect 1343 433 1520 467
rect 1112 297 1214 315
rect 1054 263 1214 297
rect 904 156 1020 207
rect 284 52 358 93
rect 684 89 718 143
rect 836 123 870 143
rect 926 141 1020 156
rect 564 55 718 89
rect 836 57 892 123
rect 1054 107 1088 263
rect 1180 249 1214 263
rect 1122 213 1156 219
rect 1248 213 1282 427
rect 1316 249 1354 393
rect 1388 315 1452 381
rect 1122 153 1282 213
rect 1388 207 1426 315
rect 1486 281 1520 433
rect 1687 381 1741 491
rect 1554 315 1741 381
rect 940 73 1088 107
rect 1248 107 1282 153
rect 1316 141 1426 207
rect 1460 265 1520 281
rect 1707 265 1741 315
rect 1460 199 1673 265
rect 1707 199 1847 265
rect 1460 107 1494 199
rect 1707 165 1741 199
rect 1248 73 1340 107
rect 1386 73 1494 107
rect 1671 60 1741 165
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< obsm1 >>
rect 116 388 174 397
rect 1029 388 1087 397
rect 1306 388 1364 397
rect 116 360 1364 388
rect 116 351 174 360
rect 1029 351 1087 360
rect 1306 351 1364 360
rect 196 184 254 193
rect 937 184 995 193
rect 1314 184 1372 193
rect 196 156 1372 184
rect 196 147 254 156
rect 937 147 995 156
rect 1314 147 1372 156
<< labels >>
rlabel locali s 19 195 89 325 6 CLK
port 1 nsew clock input
rlabel locali s 492 271 558 337 6 D
port 2 nsew signal input
rlabel locali s 706 211 798 331 6 SCD
port 3 nsew signal input
rlabel locali s 495 61 530 123 6 SCE
port 4 nsew signal input
rlabel locali s 374 123 650 127 6 SCE
port 4 nsew signal input
rlabel locali s 352 127 650 157 6 SCE
port 4 nsew signal input
rlabel locali s 613 157 650 219 6 SCE
port 4 nsew signal input
rlabel locali s 352 157 398 167 6 SCE
port 4 nsew signal input
rlabel locali s 352 167 386 337 6 SCE
port 4 nsew signal input
rlabel metal1 s 0 -48 1932 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1869 -17 1903 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1777 -17 1811 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1685 -17 1719 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1593 -17 1627 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1501 -17 1535 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1409 -17 1443 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1317 -17 1351 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1225 -17 1259 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1133 -17 1167 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 1041 -17 1075 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 949 -17 983 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 857 -17 891 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 765 -17 799 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 673 -17 707 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 581 -17 615 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 489 -17 523 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 397 -17 431 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 305 -17 339 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 213 -17 247 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 121 -17 155 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel viali s 29 -17 63 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 0 -17 1932 17 8 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1775 17 1809 139 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1543 17 1617 123 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 1138 17 1212 117 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 752 17 792 109 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 392 17 461 89 6 VGND
port 5 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 1930 145 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1022 145 1930 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 145 821 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1653 157 1930 203 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1168 157 1350 201 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1970 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1869 527 1903 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1777 527 1811 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1685 527 1719 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1593 527 1627 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1501 527 1535 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1409 527 1443 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1317 527 1351 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1225 527 1259 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1133 527 1167 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 1041 527 1075 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 949 527 983 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 857 527 891 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 765 527 799 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 673 527 707 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 581 527 615 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 489 527 523 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 397 527 431 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 305 527 339 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 213 527 247 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 121 527 155 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel viali s 29 527 63 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1775 325 1809 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1558 427 1619 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1180 367 1214 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 746 433 785 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 376 449 442 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 104 427 170 527 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 0 527 1932 561 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1846 61 1915 164 6 Q
port 9 nsew signal output
rlabel locali s 1881 164 1915 301 6 Q
port 9 nsew signal output
rlabel locali s 1846 301 1915 479 6 Q
port 9 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 376304
string GDS_START 361098
<< end >>
