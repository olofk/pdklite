magic
tech sky130A
magscale 1 2
timestamp 1619729575
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 29 -17 63 17
<< locali >>
rect 17 296 85 493
rect 17 165 68 296
rect 206 199 272 265
rect 17 90 89 165
rect 442 215 556 257
rect 590 215 719 257
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 119 441 201 527
rect 350 443 416 527
rect 450 407 515 493
rect 119 373 515 407
rect 119 265 172 373
rect 215 305 340 339
rect 102 199 172 265
rect 306 165 340 305
rect 142 17 176 165
rect 232 131 340 165
rect 374 291 515 373
rect 610 307 676 527
rect 232 90 266 131
rect 374 51 408 291
rect 454 147 688 181
rect 454 51 520 147
rect 554 17 588 111
rect 622 54 688 147
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 590 215 719 257 6 A1
port 1 nsew signal input
rlabel locali s 442 215 556 257 6 A2
port 2 nsew signal input
rlabel locali s 206 199 272 265 6 B1_N
port 3 nsew signal input
rlabel locali s 17 296 85 493 6 X
port 8 nsew signal output
rlabel locali s 17 165 68 296 6 X
port 8 nsew signal output
rlabel locali s 17 90 89 165 6 X
port 8 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1709788
string GDS_START 1703684
<< end >>
