magic
tech sky130A
timestamp 1619729571
<< checkpaint >>
rect -649 -654 1201 926
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_0
timestamp 1619729571
transform 1 0 460 0 1 0
box -19 -24 111 296
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_0
timestamp 1619729571
transform 1 0 276 0 1 0
box -19 -24 203 296
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_0
timestamp 1619729571
transform 1 0 0 0 1 0
box -19 -24 295 296
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 272
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_ef_sc_hd__fill_12.gds
string LEFsymmetry X Y R90
string GDS_END 368
string GDS_START 138
<< end >>
