magic
tech sky130A
magscale 1 2
timestamp 1640697980
<< nwell >>
rect -38 261 2154 582
<< pwell >>
rect 903 157 1089 201
rect 1633 157 2075 203
rect 1 21 2075 157
rect 29 -17 63 21
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 103 427 169 527
rect 18 195 88 325
rect 103 17 169 93
rect 271 333 336 490
rect 370 435 420 527
rect 283 123 375 333
rect 798 441 864 527
rect 991 435 1065 527
rect 1388 435 1438 527
rect 761 187 919 203
rect 761 153 833 187
rect 867 153 919 187
rect 309 17 375 89
rect 895 17 961 109
rect 1542 451 1608 527
rect 1421 250 1529 281
rect 1667 315 1701 527
rect 1743 325 1801 493
rect 1835 359 1869 527
rect 1911 325 1961 493
rect 2003 359 2037 527
rect 1743 291 2088 325
rect 1455 216 1529 250
rect 1421 207 1529 216
rect 1481 187 1529 207
rect 1341 17 1379 105
rect 1515 153 1529 187
rect 1481 127 1529 153
rect 2006 181 2088 291
rect 1667 17 1701 179
rect 1735 147 2088 181
rect 1735 51 1801 147
rect 1835 17 1869 111
rect 1903 51 1969 147
rect 2003 17 2037 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 833 153 867 187
rect 1421 216 1455 250
rect 1481 153 1515 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< obsli1 >>
rect 18 393 69 493
rect 18 359 168 393
rect 122 161 168 359
rect 18 127 168 161
rect 18 69 69 127
rect 203 69 237 493
rect 454 427 504 493
rect 547 427 683 493
rect 454 401 488 427
rect 409 367 488 401
rect 409 95 443 367
rect 522 315 615 393
rect 477 153 547 277
rect 581 197 615 315
rect 649 271 683 427
rect 717 407 751 475
rect 898 407 932 475
rect 717 373 932 407
rect 1099 401 1133 493
rect 1180 425 1354 493
rect 1021 367 1133 401
rect 1021 339 1055 367
rect 755 305 1055 339
rect 1194 333 1286 391
rect 649 237 987 271
rect 581 153 652 197
rect 686 95 720 237
rect 953 201 987 237
rect 1021 167 1055 305
rect 409 61 508 95
rect 549 61 720 95
rect 1003 89 1055 167
rect 1093 331 1286 333
rect 1320 349 1354 425
rect 1472 417 1506 475
rect 1472 383 1632 417
rect 1093 299 1228 331
rect 1320 315 1564 349
rect 1093 141 1135 299
rect 1320 297 1354 315
rect 1169 141 1239 265
rect 1273 263 1354 297
rect 1273 107 1307 263
rect 1598 259 1632 383
rect 1341 173 1385 229
rect 1341 139 1447 173
rect 1003 55 1073 89
rect 1117 51 1307 107
rect 1413 93 1447 139
rect 1563 257 1632 259
rect 1563 215 1969 257
rect 1563 164 1628 215
rect 1563 93 1627 164
rect 1413 59 1627 93
<< metal1 >>
rect 0 561 2116 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 1409 250 1467 256
rect 1409 216 1421 250
rect 1455 216 1467 250
rect 1409 193 1467 216
rect 749 187 879 193
rect 749 153 833 187
rect 867 184 879 187
rect 1409 187 1527 193
rect 1409 184 1481 187
rect 867 156 1481 184
rect 867 153 879 156
rect 749 147 879 153
rect 1469 153 1481 156
rect 1515 153 1527 187
rect 1469 147 1527 153
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
<< obsm1 >>
rect 191 388 249 397
rect 569 388 627 397
rect 1193 388 1251 397
rect 191 360 1251 388
rect 191 351 249 360
rect 569 351 627 360
rect 1193 351 1251 360
rect 110 252 168 261
rect 477 252 535 261
rect 1193 252 1251 261
rect 110 224 1251 252
rect 110 215 168 224
rect 477 215 535 224
rect 1193 215 1251 224
<< labels >>
rlabel locali s 18 195 88 325 6 CLK
port 1 nsew clock input
rlabel locali s 283 123 375 333 6 D
port 2 nsew signal input
rlabel locali s 271 333 336 490 6 D
port 2 nsew signal input
rlabel metal1 s 1469 147 1527 156 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 749 147 879 156 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 749 156 1527 184 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1409 184 1527 193 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 749 184 879 193 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1409 193 1467 256 6 RESET_B
port 3 nsew signal input
rlabel viali s 1481 153 1515 187 6 RESET_B
port 3 nsew signal input
rlabel viali s 1421 216 1455 250 6 RESET_B
port 3 nsew signal input
rlabel locali s 1481 127 1529 207 6 RESET_B
port 3 nsew signal input
rlabel locali s 1421 207 1529 281 6 RESET_B
port 3 nsew signal input
rlabel viali s 833 153 867 187 6 RESET_B
port 3 nsew signal input
rlabel locali s 761 153 919 203 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 0 -48 2116 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 2053 -17 2087 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1961 -17 1995 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1869 -17 1903 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1777 -17 1811 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1685 -17 1719 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1593 -17 1627 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1501 -17 1535 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1409 -17 1443 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1317 -17 1351 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1225 -17 1259 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1133 -17 1167 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1041 -17 1075 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 949 -17 983 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 857 -17 891 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 765 -17 799 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 673 -17 707 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 581 -17 615 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 489 -17 523 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 397 -17 431 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 305 -17 339 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 213 -17 247 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 121 -17 155 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 29 -17 63 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 2116 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 2003 17 2037 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1835 17 1869 111 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1667 17 1701 179 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1341 17 1379 105 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 895 17 961 109 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 309 17 375 89 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 2075 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1633 157 2075 203 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 903 157 1089 201 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 2154 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 2116 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 2053 527 2087 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1961 527 1995 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1869 527 1903 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1777 527 1811 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1685 527 1719 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1593 527 1627 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1501 527 1535 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1409 527 1443 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1317 527 1351 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1225 527 1259 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1133 527 1167 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1041 527 1075 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 949 527 983 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 857 527 891 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 765 527 799 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 673 527 707 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 581 527 615 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 489 527 523 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 397 527 431 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 305 527 339 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 213 527 247 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 121 527 155 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 29 527 63 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 2003 359 2037 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1835 359 1869 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1667 315 1701 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1542 451 1608 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1388 435 1438 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 991 435 1065 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 798 441 864 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 370 435 420 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 2116 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1903 51 1969 147 6 Q
port 8 nsew signal output
rlabel locali s 1735 51 1801 147 6 Q
port 8 nsew signal output
rlabel locali s 1735 147 2088 181 6 Q
port 8 nsew signal output
rlabel locali s 2006 181 2088 291 6 Q
port 8 nsew signal output
rlabel locali s 1743 291 2088 325 6 Q
port 8 nsew signal output
rlabel locali s 1911 325 1961 493 6 Q
port 8 nsew signal output
rlabel locali s 1743 325 1801 493 6 Q
port 8 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2116 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2478496
string GDS_START 2460704
<< end >>
