magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -990 -1276 17293 9368
<< nwell >>
rect 270 4019 10996 5889
<< pwell >>
rect 336 7960 16032 8042
rect 336 6057 418 7960
rect 13152 6057 16032 7960
rect 336 5975 16032 6057
rect 11482 4051 11564 5975
rect 14740 4051 16032 5975
rect 11482 4017 16032 4051
rect 336 3851 10970 3933
rect 336 2247 418 3851
rect 10888 2247 10970 3851
rect 336 2165 10970 2247
rect 11482 2093 11564 4017
rect 14740 2093 16032 4017
rect 336 2011 16032 2093
rect 336 108 418 2011
rect 13152 108 16032 2011
rect 336 26 16032 108
<< pmos >>
rect 525 5512 1325 5687
rect 1381 5512 2181 5687
rect 2237 5512 3037 5687
rect 3093 5512 3893 5687
rect 3949 5512 4749 5687
rect 4805 5512 5605 5687
rect 5661 5512 6461 5687
rect 6517 5512 7317 5687
rect 7373 5512 8173 5687
rect 8229 5512 9029 5687
rect 9085 5512 9885 5687
rect 9941 5512 10741 5687
<< mvnmos >>
rect 545 2321 1345 3721
rect 1401 2321 2201 3721
rect 2257 2321 3057 3721
rect 3113 2321 3913 3721
rect 3969 2321 4769 3721
rect 4825 2321 5625 3721
rect 5681 2321 6481 3721
rect 6537 2321 7337 3721
rect 7393 2321 8193 3721
rect 8249 2321 9049 3721
rect 9105 2321 9905 3721
rect 9961 2321 10761 3721
<< mvpmos >>
rect 525 4287 1325 5512
rect 1381 4287 2181 5512
rect 2237 4287 3037 5512
rect 3093 4287 3893 5512
rect 3949 4287 4749 5512
rect 4805 4287 5605 5512
rect 5661 4287 6461 5512
rect 6517 4287 7317 5512
rect 7373 4287 8173 5512
rect 8229 4287 9029 5512
rect 9085 4287 9885 5512
rect 9941 4287 10741 5512
<< ndiff >>
rect 472 7873 582 7906
rect 472 7839 480 7873
rect 514 7839 548 7873
rect 472 7806 582 7839
rect 3382 7873 3484 7906
rect 3416 7839 3450 7873
rect 3382 7806 3484 7839
rect 12884 7873 12994 7906
rect 12918 7839 12952 7873
rect 12986 7839 12994 7873
rect 12884 7806 12994 7839
rect 472 7719 582 7752
rect 472 7685 480 7719
rect 514 7685 548 7719
rect 472 7652 582 7685
rect 3382 7719 3484 7752
rect 3416 7685 3450 7719
rect 3382 7652 3484 7685
rect 12884 7719 12994 7752
rect 12918 7685 12952 7719
rect 12986 7685 12994 7719
rect 12884 7652 12994 7685
rect 472 7565 582 7598
rect 472 7531 480 7565
rect 514 7531 548 7565
rect 472 7498 582 7531
rect 3382 7565 3484 7598
rect 3416 7531 3450 7565
rect 3382 7498 3484 7531
rect 12884 7565 12994 7598
rect 12918 7531 12952 7565
rect 12986 7531 12994 7565
rect 12884 7498 12994 7531
rect 472 7411 582 7444
rect 472 7377 480 7411
rect 514 7377 548 7411
rect 472 7344 582 7377
rect 3382 7411 3484 7444
rect 3416 7377 3450 7411
rect 3382 7344 3484 7377
rect 12884 7411 12994 7444
rect 12918 7377 12952 7411
rect 12986 7377 12994 7411
rect 12884 7344 12994 7377
rect 472 7257 582 7290
rect 472 7223 480 7257
rect 514 7223 548 7257
rect 472 7190 582 7223
rect 3382 7257 3484 7290
rect 3416 7223 3450 7257
rect 3382 7190 3484 7223
rect 12884 7257 12994 7290
rect 12918 7223 12952 7257
rect 12986 7223 12994 7257
rect 12884 7190 12994 7223
rect 472 7103 582 7136
rect 472 7069 480 7103
rect 514 7069 548 7103
rect 472 7036 582 7069
rect 3382 7103 3484 7136
rect 3416 7069 3450 7103
rect 3382 7036 3484 7069
rect 12884 7103 12994 7136
rect 12918 7069 12952 7103
rect 12986 7069 12994 7103
rect 12884 7036 12994 7069
rect 472 6949 582 6982
rect 472 6915 480 6949
rect 514 6915 548 6949
rect 472 6882 582 6915
rect 3382 6949 3484 6982
rect 3416 6915 3450 6949
rect 3382 6882 3484 6915
rect 12884 6949 12994 6982
rect 12918 6915 12952 6949
rect 12986 6915 12994 6949
rect 12884 6882 12994 6915
rect 472 6795 582 6828
rect 472 6761 480 6795
rect 514 6761 548 6795
rect 472 6728 582 6761
rect 3382 6795 3484 6828
rect 3416 6761 3450 6795
rect 3382 6728 3484 6761
rect 12884 6795 12994 6828
rect 12918 6761 12952 6795
rect 12986 6761 12994 6795
rect 12884 6728 12994 6761
rect 472 6641 582 6674
rect 472 6607 480 6641
rect 514 6607 548 6641
rect 472 6574 582 6607
rect 3382 6641 3484 6674
rect 3416 6607 3450 6641
rect 3382 6574 3484 6607
rect 12884 6641 12994 6674
rect 12918 6607 12952 6641
rect 12986 6607 12994 6641
rect 12884 6574 12994 6607
rect 472 6487 582 6520
rect 472 6453 480 6487
rect 514 6453 548 6487
rect 472 6420 582 6453
rect 3382 6487 3484 6520
rect 3416 6453 3450 6487
rect 3382 6420 3484 6453
rect 12884 6487 12994 6520
rect 12918 6453 12952 6487
rect 12986 6453 12994 6487
rect 12884 6420 12994 6453
rect 472 6333 582 6366
rect 472 6299 480 6333
rect 514 6299 548 6333
rect 472 6266 582 6299
rect 3382 6333 3484 6366
rect 3416 6299 3450 6333
rect 3382 6266 3484 6299
rect 12884 6333 12994 6366
rect 12918 6299 12952 6333
rect 12986 6299 12994 6333
rect 12884 6266 12994 6299
rect 472 6179 582 6212
rect 472 6145 480 6179
rect 514 6145 548 6179
rect 472 6112 582 6145
rect 3382 6179 3484 6212
rect 3416 6145 3450 6179
rect 3382 6112 3484 6145
rect 12884 6179 12994 6212
rect 12918 6145 12952 6179
rect 12986 6145 12994 6179
rect 12884 6112 12994 6145
rect 11618 5888 11728 5921
rect 11618 5854 11626 5888
rect 11660 5854 11694 5888
rect 11618 5821 11728 5854
rect 14528 5888 14638 5921
rect 14562 5854 14596 5888
rect 14630 5854 14638 5888
rect 14528 5821 14638 5854
rect 11618 5734 11728 5767
rect 11618 5700 11626 5734
rect 11660 5700 11694 5734
rect 11618 5667 11728 5700
rect 14528 5734 14638 5767
rect 14562 5700 14596 5734
rect 14630 5700 14638 5734
rect 14528 5667 14638 5700
rect 11618 5580 11728 5613
rect 11618 5546 11626 5580
rect 11660 5546 11694 5580
rect 11618 5513 11728 5546
rect 14528 5580 14638 5613
rect 14562 5546 14596 5580
rect 14630 5546 14638 5580
rect 14528 5513 14638 5546
rect 11618 5426 11728 5459
rect 11618 5392 11626 5426
rect 11660 5392 11694 5426
rect 11618 5359 11728 5392
rect 14528 5426 14638 5459
rect 14562 5392 14596 5426
rect 14630 5392 14638 5426
rect 14528 5359 14638 5392
rect 11618 5272 11728 5305
rect 11618 5238 11626 5272
rect 11660 5238 11694 5272
rect 11618 5205 11728 5238
rect 14528 5272 14638 5305
rect 14562 5238 14596 5272
rect 14630 5238 14638 5272
rect 14528 5205 14638 5238
rect 11618 5118 11728 5151
rect 11618 5084 11626 5118
rect 11660 5084 11694 5118
rect 11618 5051 11728 5084
rect 14528 5118 14638 5151
rect 14562 5084 14596 5118
rect 14630 5084 14638 5118
rect 14528 5051 14638 5084
rect 11618 4964 11728 4997
rect 11618 4930 11626 4964
rect 11660 4930 11694 4964
rect 11618 4897 11728 4930
rect 14528 4964 14638 4997
rect 14562 4930 14596 4964
rect 14630 4930 14638 4964
rect 14528 4897 14638 4930
rect 11618 4810 11728 4843
rect 11618 4776 11626 4810
rect 11660 4776 11694 4810
rect 11618 4743 11728 4776
rect 14528 4810 14638 4843
rect 14562 4776 14596 4810
rect 14630 4776 14638 4810
rect 14528 4743 14638 4776
rect 11618 4656 11728 4689
rect 11618 4622 11626 4656
rect 11660 4622 11694 4656
rect 11618 4589 11728 4622
rect 14528 4656 14638 4689
rect 14562 4622 14596 4656
rect 14630 4622 14638 4656
rect 14528 4589 14638 4622
rect 11618 4502 11728 4535
rect 11618 4468 11626 4502
rect 11660 4468 11694 4502
rect 11618 4435 11728 4468
rect 14528 4502 14638 4535
rect 14562 4468 14596 4502
rect 14630 4468 14638 4502
rect 14528 4435 14638 4468
rect 11618 4348 11728 4381
rect 11618 4314 11626 4348
rect 11660 4314 11694 4348
rect 11618 4281 11728 4314
rect 14528 4348 14638 4381
rect 14562 4314 14596 4348
rect 14630 4314 14638 4348
rect 14528 4281 14638 4314
rect 11618 4194 11728 4227
rect 11618 4160 11626 4194
rect 11660 4160 11694 4194
rect 11618 4127 11728 4160
rect 14528 4194 14638 4227
rect 14562 4160 14596 4194
rect 14630 4160 14638 4194
rect 14528 4127 14638 4160
rect 11618 3908 11728 3941
rect 11618 3874 11626 3908
rect 11660 3874 11694 3908
rect 11618 3841 11728 3874
rect 14528 3908 14638 3941
rect 14562 3874 14596 3908
rect 14630 3874 14638 3908
rect 14528 3841 14638 3874
rect 11618 3754 11728 3787
rect 11618 3720 11626 3754
rect 11660 3720 11694 3754
rect 11618 3687 11728 3720
rect 14528 3754 14638 3787
rect 14562 3720 14596 3754
rect 14630 3720 14638 3754
rect 14528 3687 14638 3720
rect 11618 3600 11728 3633
rect 11618 3566 11626 3600
rect 11660 3566 11694 3600
rect 11618 3533 11728 3566
rect 14528 3600 14638 3633
rect 14562 3566 14596 3600
rect 14630 3566 14638 3600
rect 14528 3533 14638 3566
rect 11618 3446 11728 3479
rect 11618 3412 11626 3446
rect 11660 3412 11694 3446
rect 11618 3379 11728 3412
rect 14528 3446 14638 3479
rect 14562 3412 14596 3446
rect 14630 3412 14638 3446
rect 14528 3379 14638 3412
rect 11618 3292 11728 3325
rect 11618 3258 11626 3292
rect 11660 3258 11694 3292
rect 11618 3225 11728 3258
rect 14528 3292 14638 3325
rect 14562 3258 14596 3292
rect 14630 3258 14638 3292
rect 14528 3225 14638 3258
rect 11618 3138 11728 3171
rect 11618 3104 11626 3138
rect 11660 3104 11694 3138
rect 11618 3071 11728 3104
rect 14528 3138 14638 3171
rect 14562 3104 14596 3138
rect 14630 3104 14638 3138
rect 14528 3071 14638 3104
rect 11618 2984 11728 3017
rect 11618 2950 11626 2984
rect 11660 2950 11694 2984
rect 11618 2917 11728 2950
rect 14528 2984 14638 3017
rect 14562 2950 14596 2984
rect 14630 2950 14638 2984
rect 14528 2917 14638 2950
rect 11618 2830 11728 2863
rect 11618 2796 11626 2830
rect 11660 2796 11694 2830
rect 11618 2763 11728 2796
rect 14528 2830 14638 2863
rect 14562 2796 14596 2830
rect 14630 2796 14638 2830
rect 14528 2763 14638 2796
rect 11618 2676 11728 2709
rect 11618 2642 11626 2676
rect 11660 2642 11694 2676
rect 11618 2609 11728 2642
rect 14528 2676 14638 2709
rect 14562 2642 14596 2676
rect 14630 2642 14638 2676
rect 14528 2609 14638 2642
rect 11618 2522 11728 2555
rect 11618 2488 11626 2522
rect 11660 2488 11694 2522
rect 11618 2455 11728 2488
rect 14528 2522 14638 2555
rect 14562 2488 14596 2522
rect 14630 2488 14638 2522
rect 14528 2455 14638 2488
rect 11618 2368 11728 2401
rect 11618 2334 11626 2368
rect 11660 2334 11694 2368
rect 11618 2301 11728 2334
rect 14528 2368 14638 2401
rect 14562 2334 14596 2368
rect 14630 2334 14638 2368
rect 14528 2301 14638 2334
rect 11618 2214 11728 2247
rect 11618 2180 11626 2214
rect 11660 2180 11694 2214
rect 11618 2147 11728 2180
rect 14528 2214 14638 2247
rect 14562 2180 14596 2214
rect 14630 2180 14638 2214
rect 14528 2147 14638 2180
rect 472 1924 582 1957
rect 472 1890 480 1924
rect 514 1890 548 1924
rect 472 1857 582 1890
rect 3382 1924 3484 1957
rect 3416 1890 3450 1924
rect 3382 1857 3484 1890
rect 12884 1924 12994 1957
rect 12918 1890 12952 1924
rect 12986 1890 12994 1924
rect 12884 1857 12994 1890
rect 472 1770 582 1803
rect 472 1736 480 1770
rect 514 1736 548 1770
rect 472 1703 582 1736
rect 3382 1770 3484 1803
rect 3416 1736 3450 1770
rect 3382 1703 3484 1736
rect 12884 1770 12994 1803
rect 12918 1736 12952 1770
rect 12986 1736 12994 1770
rect 12884 1703 12994 1736
rect 472 1616 582 1649
rect 472 1582 480 1616
rect 514 1582 548 1616
rect 472 1549 582 1582
rect 3382 1616 3484 1649
rect 3416 1582 3450 1616
rect 3382 1549 3484 1582
rect 12884 1616 12994 1649
rect 12918 1582 12952 1616
rect 12986 1582 12994 1616
rect 12884 1549 12994 1582
rect 472 1462 582 1495
rect 472 1428 480 1462
rect 514 1428 548 1462
rect 472 1395 582 1428
rect 3382 1462 3484 1495
rect 3416 1428 3450 1462
rect 3382 1395 3484 1428
rect 12884 1462 12994 1495
rect 12918 1428 12952 1462
rect 12986 1428 12994 1462
rect 12884 1395 12994 1428
rect 472 1308 582 1341
rect 472 1274 480 1308
rect 514 1274 548 1308
rect 472 1241 582 1274
rect 3382 1308 3484 1341
rect 3416 1274 3450 1308
rect 3382 1241 3484 1274
rect 12884 1308 12994 1341
rect 12918 1274 12952 1308
rect 12986 1274 12994 1308
rect 12884 1241 12994 1274
rect 472 1154 582 1187
rect 472 1120 480 1154
rect 514 1120 548 1154
rect 472 1087 582 1120
rect 3382 1154 3484 1187
rect 3416 1120 3450 1154
rect 3382 1087 3484 1120
rect 12884 1154 12994 1187
rect 12918 1120 12952 1154
rect 12986 1120 12994 1154
rect 12884 1087 12994 1120
rect 472 1000 582 1033
rect 472 966 480 1000
rect 514 966 548 1000
rect 472 933 582 966
rect 3382 1000 3484 1033
rect 3416 966 3450 1000
rect 3382 933 3484 966
rect 12884 1000 12994 1033
rect 12918 966 12952 1000
rect 12986 966 12994 1000
rect 12884 933 12994 966
rect 472 846 582 879
rect 472 812 480 846
rect 514 812 548 846
rect 472 779 582 812
rect 3382 846 3484 879
rect 3416 812 3450 846
rect 3382 779 3484 812
rect 12884 846 12994 879
rect 12918 812 12952 846
rect 12986 812 12994 846
rect 12884 779 12994 812
rect 472 692 582 725
rect 472 658 480 692
rect 514 658 548 692
rect 472 625 582 658
rect 3382 692 3484 725
rect 3416 658 3450 692
rect 3382 625 3484 658
rect 12884 692 12994 725
rect 12918 658 12952 692
rect 12986 658 12994 692
rect 12884 625 12994 658
rect 472 538 582 571
rect 472 504 480 538
rect 514 504 548 538
rect 472 471 582 504
rect 3382 538 3484 571
rect 3416 504 3450 538
rect 3382 471 3484 504
rect 12884 538 12994 571
rect 12918 504 12952 538
rect 12986 504 12994 538
rect 12884 471 12994 504
rect 472 384 582 417
rect 472 350 480 384
rect 514 350 548 384
rect 472 317 582 350
rect 3382 384 3484 417
rect 3416 350 3450 384
rect 3382 317 3484 350
rect 12884 384 12994 417
rect 12918 350 12952 384
rect 12986 350 12994 384
rect 12884 317 12994 350
rect 472 230 582 263
rect 472 196 480 230
rect 514 196 548 230
rect 472 163 582 196
rect 3382 230 3484 263
rect 3416 196 3450 230
rect 3382 163 3484 196
rect 12884 230 12994 263
rect 12918 196 12952 230
rect 12986 196 12994 230
rect 12884 163 12994 196
<< mvndiff >>
rect 492 3659 545 3721
rect 492 3625 500 3659
rect 534 3625 545 3659
rect 492 3591 545 3625
rect 492 3557 500 3591
rect 534 3557 545 3591
rect 492 3523 545 3557
rect 492 3489 500 3523
rect 534 3489 545 3523
rect 492 3455 545 3489
rect 492 3421 500 3455
rect 534 3421 545 3455
rect 492 3387 545 3421
rect 492 3353 500 3387
rect 534 3353 545 3387
rect 492 3319 545 3353
rect 492 3285 500 3319
rect 534 3285 545 3319
rect 492 3251 545 3285
rect 492 3217 500 3251
rect 534 3217 545 3251
rect 492 3183 545 3217
rect 492 3149 500 3183
rect 534 3149 545 3183
rect 492 3115 545 3149
rect 492 3081 500 3115
rect 534 3081 545 3115
rect 492 3047 545 3081
rect 492 3013 500 3047
rect 534 3013 545 3047
rect 492 2979 545 3013
rect 492 2945 500 2979
rect 534 2945 545 2979
rect 492 2911 545 2945
rect 492 2877 500 2911
rect 534 2877 545 2911
rect 492 2843 545 2877
rect 492 2809 500 2843
rect 534 2809 545 2843
rect 492 2775 545 2809
rect 492 2741 500 2775
rect 534 2741 545 2775
rect 492 2707 545 2741
rect 492 2673 500 2707
rect 534 2673 545 2707
rect 492 2639 545 2673
rect 492 2605 500 2639
rect 534 2605 545 2639
rect 492 2571 545 2605
rect 492 2537 500 2571
rect 534 2537 545 2571
rect 492 2503 545 2537
rect 492 2469 500 2503
rect 534 2469 545 2503
rect 492 2435 545 2469
rect 492 2401 500 2435
rect 534 2401 545 2435
rect 492 2367 545 2401
rect 492 2333 500 2367
rect 534 2333 545 2367
rect 492 2321 545 2333
rect 1345 3659 1401 3721
rect 1345 3625 1356 3659
rect 1390 3625 1401 3659
rect 1345 3591 1401 3625
rect 1345 3557 1356 3591
rect 1390 3557 1401 3591
rect 1345 3523 1401 3557
rect 1345 3489 1356 3523
rect 1390 3489 1401 3523
rect 1345 3455 1401 3489
rect 1345 3421 1356 3455
rect 1390 3421 1401 3455
rect 1345 3387 1401 3421
rect 1345 3353 1356 3387
rect 1390 3353 1401 3387
rect 1345 3319 1401 3353
rect 1345 3285 1356 3319
rect 1390 3285 1401 3319
rect 1345 3251 1401 3285
rect 1345 3217 1356 3251
rect 1390 3217 1401 3251
rect 1345 3183 1401 3217
rect 1345 3149 1356 3183
rect 1390 3149 1401 3183
rect 1345 3115 1401 3149
rect 1345 3081 1356 3115
rect 1390 3081 1401 3115
rect 1345 3047 1401 3081
rect 1345 3013 1356 3047
rect 1390 3013 1401 3047
rect 1345 2979 1401 3013
rect 1345 2945 1356 2979
rect 1390 2945 1401 2979
rect 1345 2911 1401 2945
rect 1345 2877 1356 2911
rect 1390 2877 1401 2911
rect 1345 2843 1401 2877
rect 1345 2809 1356 2843
rect 1390 2809 1401 2843
rect 1345 2775 1401 2809
rect 1345 2741 1356 2775
rect 1390 2741 1401 2775
rect 1345 2707 1401 2741
rect 1345 2673 1356 2707
rect 1390 2673 1401 2707
rect 1345 2639 1401 2673
rect 1345 2605 1356 2639
rect 1390 2605 1401 2639
rect 1345 2571 1401 2605
rect 1345 2537 1356 2571
rect 1390 2537 1401 2571
rect 1345 2503 1401 2537
rect 1345 2469 1356 2503
rect 1390 2469 1401 2503
rect 1345 2435 1401 2469
rect 1345 2401 1356 2435
rect 1390 2401 1401 2435
rect 1345 2367 1401 2401
rect 1345 2333 1356 2367
rect 1390 2333 1401 2367
rect 1345 2321 1401 2333
rect 2201 3659 2257 3721
rect 2201 3625 2212 3659
rect 2246 3625 2257 3659
rect 2201 3591 2257 3625
rect 2201 3557 2212 3591
rect 2246 3557 2257 3591
rect 2201 3523 2257 3557
rect 2201 3489 2212 3523
rect 2246 3489 2257 3523
rect 2201 3455 2257 3489
rect 2201 3421 2212 3455
rect 2246 3421 2257 3455
rect 2201 3387 2257 3421
rect 2201 3353 2212 3387
rect 2246 3353 2257 3387
rect 2201 3319 2257 3353
rect 2201 3285 2212 3319
rect 2246 3285 2257 3319
rect 2201 3251 2257 3285
rect 2201 3217 2212 3251
rect 2246 3217 2257 3251
rect 2201 3183 2257 3217
rect 2201 3149 2212 3183
rect 2246 3149 2257 3183
rect 2201 3115 2257 3149
rect 2201 3081 2212 3115
rect 2246 3081 2257 3115
rect 2201 3047 2257 3081
rect 2201 3013 2212 3047
rect 2246 3013 2257 3047
rect 2201 2979 2257 3013
rect 2201 2945 2212 2979
rect 2246 2945 2257 2979
rect 2201 2911 2257 2945
rect 2201 2877 2212 2911
rect 2246 2877 2257 2911
rect 2201 2843 2257 2877
rect 2201 2809 2212 2843
rect 2246 2809 2257 2843
rect 2201 2775 2257 2809
rect 2201 2741 2212 2775
rect 2246 2741 2257 2775
rect 2201 2707 2257 2741
rect 2201 2673 2212 2707
rect 2246 2673 2257 2707
rect 2201 2639 2257 2673
rect 2201 2605 2212 2639
rect 2246 2605 2257 2639
rect 2201 2571 2257 2605
rect 2201 2537 2212 2571
rect 2246 2537 2257 2571
rect 2201 2503 2257 2537
rect 2201 2469 2212 2503
rect 2246 2469 2257 2503
rect 2201 2435 2257 2469
rect 2201 2401 2212 2435
rect 2246 2401 2257 2435
rect 2201 2367 2257 2401
rect 2201 2333 2212 2367
rect 2246 2333 2257 2367
rect 2201 2321 2257 2333
rect 3057 3659 3113 3721
rect 3057 3625 3068 3659
rect 3102 3625 3113 3659
rect 3057 3591 3113 3625
rect 3057 3557 3068 3591
rect 3102 3557 3113 3591
rect 3057 3523 3113 3557
rect 3057 3489 3068 3523
rect 3102 3489 3113 3523
rect 3057 3455 3113 3489
rect 3057 3421 3068 3455
rect 3102 3421 3113 3455
rect 3057 3387 3113 3421
rect 3057 3353 3068 3387
rect 3102 3353 3113 3387
rect 3057 3319 3113 3353
rect 3057 3285 3068 3319
rect 3102 3285 3113 3319
rect 3057 3251 3113 3285
rect 3057 3217 3068 3251
rect 3102 3217 3113 3251
rect 3057 3183 3113 3217
rect 3057 3149 3068 3183
rect 3102 3149 3113 3183
rect 3057 3115 3113 3149
rect 3057 3081 3068 3115
rect 3102 3081 3113 3115
rect 3057 3047 3113 3081
rect 3057 3013 3068 3047
rect 3102 3013 3113 3047
rect 3057 2979 3113 3013
rect 3057 2945 3068 2979
rect 3102 2945 3113 2979
rect 3057 2911 3113 2945
rect 3057 2877 3068 2911
rect 3102 2877 3113 2911
rect 3057 2843 3113 2877
rect 3057 2809 3068 2843
rect 3102 2809 3113 2843
rect 3057 2775 3113 2809
rect 3057 2741 3068 2775
rect 3102 2741 3113 2775
rect 3057 2707 3113 2741
rect 3057 2673 3068 2707
rect 3102 2673 3113 2707
rect 3057 2639 3113 2673
rect 3057 2605 3068 2639
rect 3102 2605 3113 2639
rect 3057 2571 3113 2605
rect 3057 2537 3068 2571
rect 3102 2537 3113 2571
rect 3057 2503 3113 2537
rect 3057 2469 3068 2503
rect 3102 2469 3113 2503
rect 3057 2435 3113 2469
rect 3057 2401 3068 2435
rect 3102 2401 3113 2435
rect 3057 2367 3113 2401
rect 3057 2333 3068 2367
rect 3102 2333 3113 2367
rect 3057 2321 3113 2333
rect 3913 3659 3969 3721
rect 3913 3625 3924 3659
rect 3958 3625 3969 3659
rect 3913 3591 3969 3625
rect 3913 3557 3924 3591
rect 3958 3557 3969 3591
rect 3913 3523 3969 3557
rect 3913 3489 3924 3523
rect 3958 3489 3969 3523
rect 3913 3455 3969 3489
rect 3913 3421 3924 3455
rect 3958 3421 3969 3455
rect 3913 3387 3969 3421
rect 3913 3353 3924 3387
rect 3958 3353 3969 3387
rect 3913 3319 3969 3353
rect 3913 3285 3924 3319
rect 3958 3285 3969 3319
rect 3913 3251 3969 3285
rect 3913 3217 3924 3251
rect 3958 3217 3969 3251
rect 3913 3183 3969 3217
rect 3913 3149 3924 3183
rect 3958 3149 3969 3183
rect 3913 3115 3969 3149
rect 3913 3081 3924 3115
rect 3958 3081 3969 3115
rect 3913 3047 3969 3081
rect 3913 3013 3924 3047
rect 3958 3013 3969 3047
rect 3913 2979 3969 3013
rect 3913 2945 3924 2979
rect 3958 2945 3969 2979
rect 3913 2911 3969 2945
rect 3913 2877 3924 2911
rect 3958 2877 3969 2911
rect 3913 2843 3969 2877
rect 3913 2809 3924 2843
rect 3958 2809 3969 2843
rect 3913 2775 3969 2809
rect 3913 2741 3924 2775
rect 3958 2741 3969 2775
rect 3913 2707 3969 2741
rect 3913 2673 3924 2707
rect 3958 2673 3969 2707
rect 3913 2639 3969 2673
rect 3913 2605 3924 2639
rect 3958 2605 3969 2639
rect 3913 2571 3969 2605
rect 3913 2537 3924 2571
rect 3958 2537 3969 2571
rect 3913 2503 3969 2537
rect 3913 2469 3924 2503
rect 3958 2469 3969 2503
rect 3913 2435 3969 2469
rect 3913 2401 3924 2435
rect 3958 2401 3969 2435
rect 3913 2367 3969 2401
rect 3913 2333 3924 2367
rect 3958 2333 3969 2367
rect 3913 2321 3969 2333
rect 4769 3659 4825 3721
rect 4769 3625 4780 3659
rect 4814 3625 4825 3659
rect 4769 3591 4825 3625
rect 4769 3557 4780 3591
rect 4814 3557 4825 3591
rect 4769 3523 4825 3557
rect 4769 3489 4780 3523
rect 4814 3489 4825 3523
rect 4769 3455 4825 3489
rect 4769 3421 4780 3455
rect 4814 3421 4825 3455
rect 4769 3387 4825 3421
rect 4769 3353 4780 3387
rect 4814 3353 4825 3387
rect 4769 3319 4825 3353
rect 4769 3285 4780 3319
rect 4814 3285 4825 3319
rect 4769 3251 4825 3285
rect 4769 3217 4780 3251
rect 4814 3217 4825 3251
rect 4769 3183 4825 3217
rect 4769 3149 4780 3183
rect 4814 3149 4825 3183
rect 4769 3115 4825 3149
rect 4769 3081 4780 3115
rect 4814 3081 4825 3115
rect 4769 3047 4825 3081
rect 4769 3013 4780 3047
rect 4814 3013 4825 3047
rect 4769 2979 4825 3013
rect 4769 2945 4780 2979
rect 4814 2945 4825 2979
rect 4769 2911 4825 2945
rect 4769 2877 4780 2911
rect 4814 2877 4825 2911
rect 4769 2843 4825 2877
rect 4769 2809 4780 2843
rect 4814 2809 4825 2843
rect 4769 2775 4825 2809
rect 4769 2741 4780 2775
rect 4814 2741 4825 2775
rect 4769 2707 4825 2741
rect 4769 2673 4780 2707
rect 4814 2673 4825 2707
rect 4769 2639 4825 2673
rect 4769 2605 4780 2639
rect 4814 2605 4825 2639
rect 4769 2571 4825 2605
rect 4769 2537 4780 2571
rect 4814 2537 4825 2571
rect 4769 2503 4825 2537
rect 4769 2469 4780 2503
rect 4814 2469 4825 2503
rect 4769 2435 4825 2469
rect 4769 2401 4780 2435
rect 4814 2401 4825 2435
rect 4769 2367 4825 2401
rect 4769 2333 4780 2367
rect 4814 2333 4825 2367
rect 4769 2321 4825 2333
rect 5625 3659 5681 3721
rect 5625 3625 5636 3659
rect 5670 3625 5681 3659
rect 5625 3591 5681 3625
rect 5625 3557 5636 3591
rect 5670 3557 5681 3591
rect 5625 3523 5681 3557
rect 5625 3489 5636 3523
rect 5670 3489 5681 3523
rect 5625 3455 5681 3489
rect 5625 3421 5636 3455
rect 5670 3421 5681 3455
rect 5625 3387 5681 3421
rect 5625 3353 5636 3387
rect 5670 3353 5681 3387
rect 5625 3319 5681 3353
rect 5625 3285 5636 3319
rect 5670 3285 5681 3319
rect 5625 3251 5681 3285
rect 5625 3217 5636 3251
rect 5670 3217 5681 3251
rect 5625 3183 5681 3217
rect 5625 3149 5636 3183
rect 5670 3149 5681 3183
rect 5625 3115 5681 3149
rect 5625 3081 5636 3115
rect 5670 3081 5681 3115
rect 5625 3047 5681 3081
rect 5625 3013 5636 3047
rect 5670 3013 5681 3047
rect 5625 2979 5681 3013
rect 5625 2945 5636 2979
rect 5670 2945 5681 2979
rect 5625 2911 5681 2945
rect 5625 2877 5636 2911
rect 5670 2877 5681 2911
rect 5625 2843 5681 2877
rect 5625 2809 5636 2843
rect 5670 2809 5681 2843
rect 5625 2775 5681 2809
rect 5625 2741 5636 2775
rect 5670 2741 5681 2775
rect 5625 2707 5681 2741
rect 5625 2673 5636 2707
rect 5670 2673 5681 2707
rect 5625 2639 5681 2673
rect 5625 2605 5636 2639
rect 5670 2605 5681 2639
rect 5625 2571 5681 2605
rect 5625 2537 5636 2571
rect 5670 2537 5681 2571
rect 5625 2503 5681 2537
rect 5625 2469 5636 2503
rect 5670 2469 5681 2503
rect 5625 2435 5681 2469
rect 5625 2401 5636 2435
rect 5670 2401 5681 2435
rect 5625 2367 5681 2401
rect 5625 2333 5636 2367
rect 5670 2333 5681 2367
rect 5625 2321 5681 2333
rect 6481 3659 6537 3721
rect 6481 3625 6492 3659
rect 6526 3625 6537 3659
rect 6481 3591 6537 3625
rect 6481 3557 6492 3591
rect 6526 3557 6537 3591
rect 6481 3523 6537 3557
rect 6481 3489 6492 3523
rect 6526 3489 6537 3523
rect 6481 3455 6537 3489
rect 6481 3421 6492 3455
rect 6526 3421 6537 3455
rect 6481 3387 6537 3421
rect 6481 3353 6492 3387
rect 6526 3353 6537 3387
rect 6481 3319 6537 3353
rect 6481 3285 6492 3319
rect 6526 3285 6537 3319
rect 6481 3251 6537 3285
rect 6481 3217 6492 3251
rect 6526 3217 6537 3251
rect 6481 3183 6537 3217
rect 6481 3149 6492 3183
rect 6526 3149 6537 3183
rect 6481 3115 6537 3149
rect 6481 3081 6492 3115
rect 6526 3081 6537 3115
rect 6481 3047 6537 3081
rect 6481 3013 6492 3047
rect 6526 3013 6537 3047
rect 6481 2979 6537 3013
rect 6481 2945 6492 2979
rect 6526 2945 6537 2979
rect 6481 2911 6537 2945
rect 6481 2877 6492 2911
rect 6526 2877 6537 2911
rect 6481 2843 6537 2877
rect 6481 2809 6492 2843
rect 6526 2809 6537 2843
rect 6481 2775 6537 2809
rect 6481 2741 6492 2775
rect 6526 2741 6537 2775
rect 6481 2707 6537 2741
rect 6481 2673 6492 2707
rect 6526 2673 6537 2707
rect 6481 2639 6537 2673
rect 6481 2605 6492 2639
rect 6526 2605 6537 2639
rect 6481 2571 6537 2605
rect 6481 2537 6492 2571
rect 6526 2537 6537 2571
rect 6481 2503 6537 2537
rect 6481 2469 6492 2503
rect 6526 2469 6537 2503
rect 6481 2435 6537 2469
rect 6481 2401 6492 2435
rect 6526 2401 6537 2435
rect 6481 2367 6537 2401
rect 6481 2333 6492 2367
rect 6526 2333 6537 2367
rect 6481 2321 6537 2333
rect 7337 3659 7393 3721
rect 7337 3625 7348 3659
rect 7382 3625 7393 3659
rect 7337 3591 7393 3625
rect 7337 3557 7348 3591
rect 7382 3557 7393 3591
rect 7337 3523 7393 3557
rect 7337 3489 7348 3523
rect 7382 3489 7393 3523
rect 7337 3455 7393 3489
rect 7337 3421 7348 3455
rect 7382 3421 7393 3455
rect 7337 3387 7393 3421
rect 7337 3353 7348 3387
rect 7382 3353 7393 3387
rect 7337 3319 7393 3353
rect 7337 3285 7348 3319
rect 7382 3285 7393 3319
rect 7337 3251 7393 3285
rect 7337 3217 7348 3251
rect 7382 3217 7393 3251
rect 7337 3183 7393 3217
rect 7337 3149 7348 3183
rect 7382 3149 7393 3183
rect 7337 3115 7393 3149
rect 7337 3081 7348 3115
rect 7382 3081 7393 3115
rect 7337 3047 7393 3081
rect 7337 3013 7348 3047
rect 7382 3013 7393 3047
rect 7337 2979 7393 3013
rect 7337 2945 7348 2979
rect 7382 2945 7393 2979
rect 7337 2911 7393 2945
rect 7337 2877 7348 2911
rect 7382 2877 7393 2911
rect 7337 2843 7393 2877
rect 7337 2809 7348 2843
rect 7382 2809 7393 2843
rect 7337 2775 7393 2809
rect 7337 2741 7348 2775
rect 7382 2741 7393 2775
rect 7337 2707 7393 2741
rect 7337 2673 7348 2707
rect 7382 2673 7393 2707
rect 7337 2639 7393 2673
rect 7337 2605 7348 2639
rect 7382 2605 7393 2639
rect 7337 2571 7393 2605
rect 7337 2537 7348 2571
rect 7382 2537 7393 2571
rect 7337 2503 7393 2537
rect 7337 2469 7348 2503
rect 7382 2469 7393 2503
rect 7337 2435 7393 2469
rect 7337 2401 7348 2435
rect 7382 2401 7393 2435
rect 7337 2367 7393 2401
rect 7337 2333 7348 2367
rect 7382 2333 7393 2367
rect 7337 2321 7393 2333
rect 8193 3659 8249 3721
rect 8193 3625 8204 3659
rect 8238 3625 8249 3659
rect 8193 3591 8249 3625
rect 8193 3557 8204 3591
rect 8238 3557 8249 3591
rect 8193 3523 8249 3557
rect 8193 3489 8204 3523
rect 8238 3489 8249 3523
rect 8193 3455 8249 3489
rect 8193 3421 8204 3455
rect 8238 3421 8249 3455
rect 8193 3387 8249 3421
rect 8193 3353 8204 3387
rect 8238 3353 8249 3387
rect 8193 3319 8249 3353
rect 8193 3285 8204 3319
rect 8238 3285 8249 3319
rect 8193 3251 8249 3285
rect 8193 3217 8204 3251
rect 8238 3217 8249 3251
rect 8193 3183 8249 3217
rect 8193 3149 8204 3183
rect 8238 3149 8249 3183
rect 8193 3115 8249 3149
rect 8193 3081 8204 3115
rect 8238 3081 8249 3115
rect 8193 3047 8249 3081
rect 8193 3013 8204 3047
rect 8238 3013 8249 3047
rect 8193 2979 8249 3013
rect 8193 2945 8204 2979
rect 8238 2945 8249 2979
rect 8193 2911 8249 2945
rect 8193 2877 8204 2911
rect 8238 2877 8249 2911
rect 8193 2843 8249 2877
rect 8193 2809 8204 2843
rect 8238 2809 8249 2843
rect 8193 2775 8249 2809
rect 8193 2741 8204 2775
rect 8238 2741 8249 2775
rect 8193 2707 8249 2741
rect 8193 2673 8204 2707
rect 8238 2673 8249 2707
rect 8193 2639 8249 2673
rect 8193 2605 8204 2639
rect 8238 2605 8249 2639
rect 8193 2571 8249 2605
rect 8193 2537 8204 2571
rect 8238 2537 8249 2571
rect 8193 2503 8249 2537
rect 8193 2469 8204 2503
rect 8238 2469 8249 2503
rect 8193 2435 8249 2469
rect 8193 2401 8204 2435
rect 8238 2401 8249 2435
rect 8193 2367 8249 2401
rect 8193 2333 8204 2367
rect 8238 2333 8249 2367
rect 8193 2321 8249 2333
rect 9049 3659 9105 3721
rect 9049 3625 9060 3659
rect 9094 3625 9105 3659
rect 9049 3591 9105 3625
rect 9049 3557 9060 3591
rect 9094 3557 9105 3591
rect 9049 3523 9105 3557
rect 9049 3489 9060 3523
rect 9094 3489 9105 3523
rect 9049 3455 9105 3489
rect 9049 3421 9060 3455
rect 9094 3421 9105 3455
rect 9049 3387 9105 3421
rect 9049 3353 9060 3387
rect 9094 3353 9105 3387
rect 9049 3319 9105 3353
rect 9049 3285 9060 3319
rect 9094 3285 9105 3319
rect 9049 3251 9105 3285
rect 9049 3217 9060 3251
rect 9094 3217 9105 3251
rect 9049 3183 9105 3217
rect 9049 3149 9060 3183
rect 9094 3149 9105 3183
rect 9049 3115 9105 3149
rect 9049 3081 9060 3115
rect 9094 3081 9105 3115
rect 9049 3047 9105 3081
rect 9049 3013 9060 3047
rect 9094 3013 9105 3047
rect 9049 2979 9105 3013
rect 9049 2945 9060 2979
rect 9094 2945 9105 2979
rect 9049 2911 9105 2945
rect 9049 2877 9060 2911
rect 9094 2877 9105 2911
rect 9049 2843 9105 2877
rect 9049 2809 9060 2843
rect 9094 2809 9105 2843
rect 9049 2775 9105 2809
rect 9049 2741 9060 2775
rect 9094 2741 9105 2775
rect 9049 2707 9105 2741
rect 9049 2673 9060 2707
rect 9094 2673 9105 2707
rect 9049 2639 9105 2673
rect 9049 2605 9060 2639
rect 9094 2605 9105 2639
rect 9049 2571 9105 2605
rect 9049 2537 9060 2571
rect 9094 2537 9105 2571
rect 9049 2503 9105 2537
rect 9049 2469 9060 2503
rect 9094 2469 9105 2503
rect 9049 2435 9105 2469
rect 9049 2401 9060 2435
rect 9094 2401 9105 2435
rect 9049 2367 9105 2401
rect 9049 2333 9060 2367
rect 9094 2333 9105 2367
rect 9049 2321 9105 2333
rect 9905 3659 9961 3721
rect 9905 3625 9916 3659
rect 9950 3625 9961 3659
rect 9905 3591 9961 3625
rect 9905 3557 9916 3591
rect 9950 3557 9961 3591
rect 9905 3523 9961 3557
rect 9905 3489 9916 3523
rect 9950 3489 9961 3523
rect 9905 3455 9961 3489
rect 9905 3421 9916 3455
rect 9950 3421 9961 3455
rect 9905 3387 9961 3421
rect 9905 3353 9916 3387
rect 9950 3353 9961 3387
rect 9905 3319 9961 3353
rect 9905 3285 9916 3319
rect 9950 3285 9961 3319
rect 9905 3251 9961 3285
rect 9905 3217 9916 3251
rect 9950 3217 9961 3251
rect 9905 3183 9961 3217
rect 9905 3149 9916 3183
rect 9950 3149 9961 3183
rect 9905 3115 9961 3149
rect 9905 3081 9916 3115
rect 9950 3081 9961 3115
rect 9905 3047 9961 3081
rect 9905 3013 9916 3047
rect 9950 3013 9961 3047
rect 9905 2979 9961 3013
rect 9905 2945 9916 2979
rect 9950 2945 9961 2979
rect 9905 2911 9961 2945
rect 9905 2877 9916 2911
rect 9950 2877 9961 2911
rect 9905 2843 9961 2877
rect 9905 2809 9916 2843
rect 9950 2809 9961 2843
rect 9905 2775 9961 2809
rect 9905 2741 9916 2775
rect 9950 2741 9961 2775
rect 9905 2707 9961 2741
rect 9905 2673 9916 2707
rect 9950 2673 9961 2707
rect 9905 2639 9961 2673
rect 9905 2605 9916 2639
rect 9950 2605 9961 2639
rect 9905 2571 9961 2605
rect 9905 2537 9916 2571
rect 9950 2537 9961 2571
rect 9905 2503 9961 2537
rect 9905 2469 9916 2503
rect 9950 2469 9961 2503
rect 9905 2435 9961 2469
rect 9905 2401 9916 2435
rect 9950 2401 9961 2435
rect 9905 2367 9961 2401
rect 9905 2333 9916 2367
rect 9950 2333 9961 2367
rect 9905 2321 9961 2333
rect 10761 3659 10814 3721
rect 10761 3625 10772 3659
rect 10806 3625 10814 3659
rect 10761 3591 10814 3625
rect 10761 3557 10772 3591
rect 10806 3557 10814 3591
rect 10761 3523 10814 3557
rect 10761 3489 10772 3523
rect 10806 3489 10814 3523
rect 10761 3455 10814 3489
rect 10761 3421 10772 3455
rect 10806 3421 10814 3455
rect 10761 3387 10814 3421
rect 10761 3353 10772 3387
rect 10806 3353 10814 3387
rect 10761 3319 10814 3353
rect 10761 3285 10772 3319
rect 10806 3285 10814 3319
rect 10761 3251 10814 3285
rect 10761 3217 10772 3251
rect 10806 3217 10814 3251
rect 10761 3183 10814 3217
rect 10761 3149 10772 3183
rect 10806 3149 10814 3183
rect 10761 3115 10814 3149
rect 10761 3081 10772 3115
rect 10806 3081 10814 3115
rect 10761 3047 10814 3081
rect 10761 3013 10772 3047
rect 10806 3013 10814 3047
rect 10761 2979 10814 3013
rect 10761 2945 10772 2979
rect 10806 2945 10814 2979
rect 10761 2911 10814 2945
rect 10761 2877 10772 2911
rect 10806 2877 10814 2911
rect 10761 2843 10814 2877
rect 10761 2809 10772 2843
rect 10806 2809 10814 2843
rect 10761 2775 10814 2809
rect 10761 2741 10772 2775
rect 10806 2741 10814 2775
rect 10761 2707 10814 2741
rect 10761 2673 10772 2707
rect 10806 2673 10814 2707
rect 10761 2639 10814 2673
rect 10761 2605 10772 2639
rect 10806 2605 10814 2639
rect 10761 2571 10814 2605
rect 10761 2537 10772 2571
rect 10806 2537 10814 2571
rect 10761 2503 10814 2537
rect 10761 2469 10772 2503
rect 10806 2469 10814 2503
rect 10761 2435 10814 2469
rect 10761 2401 10772 2435
rect 10806 2401 10814 2435
rect 10761 2367 10814 2401
rect 10761 2333 10772 2367
rect 10806 2333 10814 2367
rect 10761 2321 10814 2333
<< mvpdiff >>
rect 472 5625 525 5687
rect 472 5591 480 5625
rect 514 5591 525 5625
rect 472 5557 525 5591
rect 472 5523 480 5557
rect 514 5523 525 5557
rect 472 5489 525 5523
rect 1325 5625 1381 5687
rect 1325 5591 1336 5625
rect 1370 5591 1381 5625
rect 1325 5557 1381 5591
rect 1325 5523 1336 5557
rect 1370 5523 1381 5557
rect 472 5455 480 5489
rect 514 5455 525 5489
rect 472 5421 525 5455
rect 472 5387 480 5421
rect 514 5387 525 5421
rect 472 5353 525 5387
rect 472 5319 480 5353
rect 514 5319 525 5353
rect 472 5285 525 5319
rect 472 5251 480 5285
rect 514 5251 525 5285
rect 472 5217 525 5251
rect 472 5183 480 5217
rect 514 5183 525 5217
rect 472 5149 525 5183
rect 472 5115 480 5149
rect 514 5115 525 5149
rect 472 5081 525 5115
rect 472 5047 480 5081
rect 514 5047 525 5081
rect 472 5013 525 5047
rect 472 4979 480 5013
rect 514 4979 525 5013
rect 472 4945 525 4979
rect 472 4911 480 4945
rect 514 4911 525 4945
rect 472 4877 525 4911
rect 472 4843 480 4877
rect 514 4843 525 4877
rect 472 4809 525 4843
rect 472 4775 480 4809
rect 514 4775 525 4809
rect 472 4741 525 4775
rect 472 4707 480 4741
rect 514 4707 525 4741
rect 472 4673 525 4707
rect 472 4639 480 4673
rect 514 4639 525 4673
rect 472 4605 525 4639
rect 472 4571 480 4605
rect 514 4571 525 4605
rect 472 4537 525 4571
rect 472 4503 480 4537
rect 514 4503 525 4537
rect 472 4469 525 4503
rect 472 4435 480 4469
rect 514 4435 525 4469
rect 472 4401 525 4435
rect 472 4367 480 4401
rect 514 4367 525 4401
rect 472 4333 525 4367
rect 472 4299 480 4333
rect 514 4299 525 4333
rect 472 4287 525 4299
rect 1325 5489 1381 5523
rect 2181 5625 2237 5687
rect 2181 5591 2192 5625
rect 2226 5591 2237 5625
rect 2181 5557 2237 5591
rect 2181 5523 2192 5557
rect 2226 5523 2237 5557
rect 1325 5455 1336 5489
rect 1370 5455 1381 5489
rect 1325 5421 1381 5455
rect 1325 5387 1336 5421
rect 1370 5387 1381 5421
rect 1325 5353 1381 5387
rect 1325 5319 1336 5353
rect 1370 5319 1381 5353
rect 1325 5285 1381 5319
rect 1325 5251 1336 5285
rect 1370 5251 1381 5285
rect 1325 5217 1381 5251
rect 1325 5183 1336 5217
rect 1370 5183 1381 5217
rect 1325 5149 1381 5183
rect 1325 5115 1336 5149
rect 1370 5115 1381 5149
rect 1325 5081 1381 5115
rect 1325 5047 1336 5081
rect 1370 5047 1381 5081
rect 1325 5013 1381 5047
rect 1325 4979 1336 5013
rect 1370 4979 1381 5013
rect 1325 4945 1381 4979
rect 1325 4911 1336 4945
rect 1370 4911 1381 4945
rect 1325 4877 1381 4911
rect 1325 4843 1336 4877
rect 1370 4843 1381 4877
rect 1325 4809 1381 4843
rect 1325 4775 1336 4809
rect 1370 4775 1381 4809
rect 1325 4741 1381 4775
rect 1325 4707 1336 4741
rect 1370 4707 1381 4741
rect 1325 4673 1381 4707
rect 1325 4639 1336 4673
rect 1370 4639 1381 4673
rect 1325 4605 1381 4639
rect 1325 4571 1336 4605
rect 1370 4571 1381 4605
rect 1325 4537 1381 4571
rect 1325 4503 1336 4537
rect 1370 4503 1381 4537
rect 1325 4469 1381 4503
rect 1325 4435 1336 4469
rect 1370 4435 1381 4469
rect 1325 4401 1381 4435
rect 1325 4367 1336 4401
rect 1370 4367 1381 4401
rect 1325 4333 1381 4367
rect 1325 4299 1336 4333
rect 1370 4299 1381 4333
rect 1325 4287 1381 4299
rect 2181 5489 2237 5523
rect 3037 5625 3093 5687
rect 3037 5591 3048 5625
rect 3082 5591 3093 5625
rect 3037 5557 3093 5591
rect 3037 5523 3048 5557
rect 3082 5523 3093 5557
rect 2181 5455 2192 5489
rect 2226 5455 2237 5489
rect 2181 5421 2237 5455
rect 2181 5387 2192 5421
rect 2226 5387 2237 5421
rect 2181 5353 2237 5387
rect 2181 5319 2192 5353
rect 2226 5319 2237 5353
rect 2181 5285 2237 5319
rect 2181 5251 2192 5285
rect 2226 5251 2237 5285
rect 2181 5217 2237 5251
rect 2181 5183 2192 5217
rect 2226 5183 2237 5217
rect 2181 5149 2237 5183
rect 2181 5115 2192 5149
rect 2226 5115 2237 5149
rect 2181 5081 2237 5115
rect 2181 5047 2192 5081
rect 2226 5047 2237 5081
rect 2181 5013 2237 5047
rect 2181 4979 2192 5013
rect 2226 4979 2237 5013
rect 2181 4945 2237 4979
rect 2181 4911 2192 4945
rect 2226 4911 2237 4945
rect 2181 4877 2237 4911
rect 2181 4843 2192 4877
rect 2226 4843 2237 4877
rect 2181 4809 2237 4843
rect 2181 4775 2192 4809
rect 2226 4775 2237 4809
rect 2181 4741 2237 4775
rect 2181 4707 2192 4741
rect 2226 4707 2237 4741
rect 2181 4673 2237 4707
rect 2181 4639 2192 4673
rect 2226 4639 2237 4673
rect 2181 4605 2237 4639
rect 2181 4571 2192 4605
rect 2226 4571 2237 4605
rect 2181 4537 2237 4571
rect 2181 4503 2192 4537
rect 2226 4503 2237 4537
rect 2181 4469 2237 4503
rect 2181 4435 2192 4469
rect 2226 4435 2237 4469
rect 2181 4401 2237 4435
rect 2181 4367 2192 4401
rect 2226 4367 2237 4401
rect 2181 4333 2237 4367
rect 2181 4299 2192 4333
rect 2226 4299 2237 4333
rect 2181 4287 2237 4299
rect 3037 5489 3093 5523
rect 3893 5625 3949 5687
rect 3893 5591 3904 5625
rect 3938 5591 3949 5625
rect 3893 5557 3949 5591
rect 3893 5523 3904 5557
rect 3938 5523 3949 5557
rect 3037 5455 3048 5489
rect 3082 5455 3093 5489
rect 3037 5421 3093 5455
rect 3037 5387 3048 5421
rect 3082 5387 3093 5421
rect 3037 5353 3093 5387
rect 3037 5319 3048 5353
rect 3082 5319 3093 5353
rect 3037 5285 3093 5319
rect 3037 5251 3048 5285
rect 3082 5251 3093 5285
rect 3037 5217 3093 5251
rect 3037 5183 3048 5217
rect 3082 5183 3093 5217
rect 3037 5149 3093 5183
rect 3037 5115 3048 5149
rect 3082 5115 3093 5149
rect 3037 5081 3093 5115
rect 3037 5047 3048 5081
rect 3082 5047 3093 5081
rect 3037 5013 3093 5047
rect 3037 4979 3048 5013
rect 3082 4979 3093 5013
rect 3037 4945 3093 4979
rect 3037 4911 3048 4945
rect 3082 4911 3093 4945
rect 3037 4877 3093 4911
rect 3037 4843 3048 4877
rect 3082 4843 3093 4877
rect 3037 4809 3093 4843
rect 3037 4775 3048 4809
rect 3082 4775 3093 4809
rect 3037 4741 3093 4775
rect 3037 4707 3048 4741
rect 3082 4707 3093 4741
rect 3037 4673 3093 4707
rect 3037 4639 3048 4673
rect 3082 4639 3093 4673
rect 3037 4605 3093 4639
rect 3037 4571 3048 4605
rect 3082 4571 3093 4605
rect 3037 4537 3093 4571
rect 3037 4503 3048 4537
rect 3082 4503 3093 4537
rect 3037 4469 3093 4503
rect 3037 4435 3048 4469
rect 3082 4435 3093 4469
rect 3037 4401 3093 4435
rect 3037 4367 3048 4401
rect 3082 4367 3093 4401
rect 3037 4333 3093 4367
rect 3037 4299 3048 4333
rect 3082 4299 3093 4333
rect 3037 4287 3093 4299
rect 3893 5489 3949 5523
rect 4749 5625 4805 5687
rect 4749 5591 4760 5625
rect 4794 5591 4805 5625
rect 4749 5557 4805 5591
rect 4749 5523 4760 5557
rect 4794 5523 4805 5557
rect 3893 5455 3904 5489
rect 3938 5455 3949 5489
rect 3893 5421 3949 5455
rect 3893 5387 3904 5421
rect 3938 5387 3949 5421
rect 3893 5353 3949 5387
rect 3893 5319 3904 5353
rect 3938 5319 3949 5353
rect 3893 5285 3949 5319
rect 3893 5251 3904 5285
rect 3938 5251 3949 5285
rect 3893 5217 3949 5251
rect 3893 5183 3904 5217
rect 3938 5183 3949 5217
rect 3893 5149 3949 5183
rect 3893 5115 3904 5149
rect 3938 5115 3949 5149
rect 3893 5081 3949 5115
rect 3893 5047 3904 5081
rect 3938 5047 3949 5081
rect 3893 5013 3949 5047
rect 3893 4979 3904 5013
rect 3938 4979 3949 5013
rect 3893 4945 3949 4979
rect 3893 4911 3904 4945
rect 3938 4911 3949 4945
rect 3893 4877 3949 4911
rect 3893 4843 3904 4877
rect 3938 4843 3949 4877
rect 3893 4809 3949 4843
rect 3893 4775 3904 4809
rect 3938 4775 3949 4809
rect 3893 4741 3949 4775
rect 3893 4707 3904 4741
rect 3938 4707 3949 4741
rect 3893 4673 3949 4707
rect 3893 4639 3904 4673
rect 3938 4639 3949 4673
rect 3893 4605 3949 4639
rect 3893 4571 3904 4605
rect 3938 4571 3949 4605
rect 3893 4537 3949 4571
rect 3893 4503 3904 4537
rect 3938 4503 3949 4537
rect 3893 4469 3949 4503
rect 3893 4435 3904 4469
rect 3938 4435 3949 4469
rect 3893 4401 3949 4435
rect 3893 4367 3904 4401
rect 3938 4367 3949 4401
rect 3893 4333 3949 4367
rect 3893 4299 3904 4333
rect 3938 4299 3949 4333
rect 3893 4287 3949 4299
rect 4749 5489 4805 5523
rect 5605 5625 5661 5687
rect 5605 5591 5616 5625
rect 5650 5591 5661 5625
rect 5605 5557 5661 5591
rect 5605 5523 5616 5557
rect 5650 5523 5661 5557
rect 4749 5455 4760 5489
rect 4794 5455 4805 5489
rect 4749 5421 4805 5455
rect 4749 5387 4760 5421
rect 4794 5387 4805 5421
rect 4749 5353 4805 5387
rect 4749 5319 4760 5353
rect 4794 5319 4805 5353
rect 4749 5285 4805 5319
rect 4749 5251 4760 5285
rect 4794 5251 4805 5285
rect 4749 5217 4805 5251
rect 4749 5183 4760 5217
rect 4794 5183 4805 5217
rect 4749 5149 4805 5183
rect 4749 5115 4760 5149
rect 4794 5115 4805 5149
rect 4749 5081 4805 5115
rect 4749 5047 4760 5081
rect 4794 5047 4805 5081
rect 4749 5013 4805 5047
rect 4749 4979 4760 5013
rect 4794 4979 4805 5013
rect 4749 4945 4805 4979
rect 4749 4911 4760 4945
rect 4794 4911 4805 4945
rect 4749 4877 4805 4911
rect 4749 4843 4760 4877
rect 4794 4843 4805 4877
rect 4749 4809 4805 4843
rect 4749 4775 4760 4809
rect 4794 4775 4805 4809
rect 4749 4741 4805 4775
rect 4749 4707 4760 4741
rect 4794 4707 4805 4741
rect 4749 4673 4805 4707
rect 4749 4639 4760 4673
rect 4794 4639 4805 4673
rect 4749 4605 4805 4639
rect 4749 4571 4760 4605
rect 4794 4571 4805 4605
rect 4749 4537 4805 4571
rect 4749 4503 4760 4537
rect 4794 4503 4805 4537
rect 4749 4469 4805 4503
rect 4749 4435 4760 4469
rect 4794 4435 4805 4469
rect 4749 4401 4805 4435
rect 4749 4367 4760 4401
rect 4794 4367 4805 4401
rect 4749 4333 4805 4367
rect 4749 4299 4760 4333
rect 4794 4299 4805 4333
rect 4749 4287 4805 4299
rect 5605 5489 5661 5523
rect 6461 5625 6517 5687
rect 6461 5591 6472 5625
rect 6506 5591 6517 5625
rect 6461 5557 6517 5591
rect 6461 5523 6472 5557
rect 6506 5523 6517 5557
rect 5605 5455 5616 5489
rect 5650 5455 5661 5489
rect 5605 5421 5661 5455
rect 5605 5387 5616 5421
rect 5650 5387 5661 5421
rect 5605 5353 5661 5387
rect 5605 5319 5616 5353
rect 5650 5319 5661 5353
rect 5605 5285 5661 5319
rect 5605 5251 5616 5285
rect 5650 5251 5661 5285
rect 5605 5217 5661 5251
rect 5605 5183 5616 5217
rect 5650 5183 5661 5217
rect 5605 5149 5661 5183
rect 5605 5115 5616 5149
rect 5650 5115 5661 5149
rect 5605 5081 5661 5115
rect 5605 5047 5616 5081
rect 5650 5047 5661 5081
rect 5605 5013 5661 5047
rect 5605 4979 5616 5013
rect 5650 4979 5661 5013
rect 5605 4945 5661 4979
rect 5605 4911 5616 4945
rect 5650 4911 5661 4945
rect 5605 4877 5661 4911
rect 5605 4843 5616 4877
rect 5650 4843 5661 4877
rect 5605 4809 5661 4843
rect 5605 4775 5616 4809
rect 5650 4775 5661 4809
rect 5605 4741 5661 4775
rect 5605 4707 5616 4741
rect 5650 4707 5661 4741
rect 5605 4673 5661 4707
rect 5605 4639 5616 4673
rect 5650 4639 5661 4673
rect 5605 4605 5661 4639
rect 5605 4571 5616 4605
rect 5650 4571 5661 4605
rect 5605 4537 5661 4571
rect 5605 4503 5616 4537
rect 5650 4503 5661 4537
rect 5605 4469 5661 4503
rect 5605 4435 5616 4469
rect 5650 4435 5661 4469
rect 5605 4401 5661 4435
rect 5605 4367 5616 4401
rect 5650 4367 5661 4401
rect 5605 4333 5661 4367
rect 5605 4299 5616 4333
rect 5650 4299 5661 4333
rect 5605 4287 5661 4299
rect 6461 5489 6517 5523
rect 7317 5625 7373 5687
rect 7317 5591 7328 5625
rect 7362 5591 7373 5625
rect 7317 5557 7373 5591
rect 7317 5523 7328 5557
rect 7362 5523 7373 5557
rect 6461 5455 6472 5489
rect 6506 5455 6517 5489
rect 6461 5421 6517 5455
rect 6461 5387 6472 5421
rect 6506 5387 6517 5421
rect 6461 5353 6517 5387
rect 6461 5319 6472 5353
rect 6506 5319 6517 5353
rect 6461 5285 6517 5319
rect 6461 5251 6472 5285
rect 6506 5251 6517 5285
rect 6461 5217 6517 5251
rect 6461 5183 6472 5217
rect 6506 5183 6517 5217
rect 6461 5149 6517 5183
rect 6461 5115 6472 5149
rect 6506 5115 6517 5149
rect 6461 5081 6517 5115
rect 6461 5047 6472 5081
rect 6506 5047 6517 5081
rect 6461 5013 6517 5047
rect 6461 4979 6472 5013
rect 6506 4979 6517 5013
rect 6461 4945 6517 4979
rect 6461 4911 6472 4945
rect 6506 4911 6517 4945
rect 6461 4877 6517 4911
rect 6461 4843 6472 4877
rect 6506 4843 6517 4877
rect 6461 4809 6517 4843
rect 6461 4775 6472 4809
rect 6506 4775 6517 4809
rect 6461 4741 6517 4775
rect 6461 4707 6472 4741
rect 6506 4707 6517 4741
rect 6461 4673 6517 4707
rect 6461 4639 6472 4673
rect 6506 4639 6517 4673
rect 6461 4605 6517 4639
rect 6461 4571 6472 4605
rect 6506 4571 6517 4605
rect 6461 4537 6517 4571
rect 6461 4503 6472 4537
rect 6506 4503 6517 4537
rect 6461 4469 6517 4503
rect 6461 4435 6472 4469
rect 6506 4435 6517 4469
rect 6461 4401 6517 4435
rect 6461 4367 6472 4401
rect 6506 4367 6517 4401
rect 6461 4333 6517 4367
rect 6461 4299 6472 4333
rect 6506 4299 6517 4333
rect 6461 4287 6517 4299
rect 7317 5489 7373 5523
rect 8173 5625 8229 5687
rect 8173 5591 8184 5625
rect 8218 5591 8229 5625
rect 8173 5557 8229 5591
rect 8173 5523 8184 5557
rect 8218 5523 8229 5557
rect 7317 5455 7328 5489
rect 7362 5455 7373 5489
rect 7317 5421 7373 5455
rect 7317 5387 7328 5421
rect 7362 5387 7373 5421
rect 7317 5353 7373 5387
rect 7317 5319 7328 5353
rect 7362 5319 7373 5353
rect 7317 5285 7373 5319
rect 7317 5251 7328 5285
rect 7362 5251 7373 5285
rect 7317 5217 7373 5251
rect 7317 5183 7328 5217
rect 7362 5183 7373 5217
rect 7317 5149 7373 5183
rect 7317 5115 7328 5149
rect 7362 5115 7373 5149
rect 7317 5081 7373 5115
rect 7317 5047 7328 5081
rect 7362 5047 7373 5081
rect 7317 5013 7373 5047
rect 7317 4979 7328 5013
rect 7362 4979 7373 5013
rect 7317 4945 7373 4979
rect 7317 4911 7328 4945
rect 7362 4911 7373 4945
rect 7317 4877 7373 4911
rect 7317 4843 7328 4877
rect 7362 4843 7373 4877
rect 7317 4809 7373 4843
rect 7317 4775 7328 4809
rect 7362 4775 7373 4809
rect 7317 4741 7373 4775
rect 7317 4707 7328 4741
rect 7362 4707 7373 4741
rect 7317 4673 7373 4707
rect 7317 4639 7328 4673
rect 7362 4639 7373 4673
rect 7317 4605 7373 4639
rect 7317 4571 7328 4605
rect 7362 4571 7373 4605
rect 7317 4537 7373 4571
rect 7317 4503 7328 4537
rect 7362 4503 7373 4537
rect 7317 4469 7373 4503
rect 7317 4435 7328 4469
rect 7362 4435 7373 4469
rect 7317 4401 7373 4435
rect 7317 4367 7328 4401
rect 7362 4367 7373 4401
rect 7317 4333 7373 4367
rect 7317 4299 7328 4333
rect 7362 4299 7373 4333
rect 7317 4287 7373 4299
rect 8173 5489 8229 5523
rect 9029 5625 9085 5687
rect 9029 5591 9040 5625
rect 9074 5591 9085 5625
rect 9029 5557 9085 5591
rect 9029 5523 9040 5557
rect 9074 5523 9085 5557
rect 8173 5455 8184 5489
rect 8218 5455 8229 5489
rect 8173 5421 8229 5455
rect 8173 5387 8184 5421
rect 8218 5387 8229 5421
rect 8173 5353 8229 5387
rect 8173 5319 8184 5353
rect 8218 5319 8229 5353
rect 8173 5285 8229 5319
rect 8173 5251 8184 5285
rect 8218 5251 8229 5285
rect 8173 5217 8229 5251
rect 8173 5183 8184 5217
rect 8218 5183 8229 5217
rect 8173 5149 8229 5183
rect 8173 5115 8184 5149
rect 8218 5115 8229 5149
rect 8173 5081 8229 5115
rect 8173 5047 8184 5081
rect 8218 5047 8229 5081
rect 8173 5013 8229 5047
rect 8173 4979 8184 5013
rect 8218 4979 8229 5013
rect 8173 4945 8229 4979
rect 8173 4911 8184 4945
rect 8218 4911 8229 4945
rect 8173 4877 8229 4911
rect 8173 4843 8184 4877
rect 8218 4843 8229 4877
rect 8173 4809 8229 4843
rect 8173 4775 8184 4809
rect 8218 4775 8229 4809
rect 8173 4741 8229 4775
rect 8173 4707 8184 4741
rect 8218 4707 8229 4741
rect 8173 4673 8229 4707
rect 8173 4639 8184 4673
rect 8218 4639 8229 4673
rect 8173 4605 8229 4639
rect 8173 4571 8184 4605
rect 8218 4571 8229 4605
rect 8173 4537 8229 4571
rect 8173 4503 8184 4537
rect 8218 4503 8229 4537
rect 8173 4469 8229 4503
rect 8173 4435 8184 4469
rect 8218 4435 8229 4469
rect 8173 4401 8229 4435
rect 8173 4367 8184 4401
rect 8218 4367 8229 4401
rect 8173 4333 8229 4367
rect 8173 4299 8184 4333
rect 8218 4299 8229 4333
rect 8173 4287 8229 4299
rect 9029 5489 9085 5523
rect 9885 5625 9941 5687
rect 9885 5591 9896 5625
rect 9930 5591 9941 5625
rect 9885 5557 9941 5591
rect 9885 5523 9896 5557
rect 9930 5523 9941 5557
rect 9029 5455 9040 5489
rect 9074 5455 9085 5489
rect 9029 5421 9085 5455
rect 9029 5387 9040 5421
rect 9074 5387 9085 5421
rect 9029 5353 9085 5387
rect 9029 5319 9040 5353
rect 9074 5319 9085 5353
rect 9029 5285 9085 5319
rect 9029 5251 9040 5285
rect 9074 5251 9085 5285
rect 9029 5217 9085 5251
rect 9029 5183 9040 5217
rect 9074 5183 9085 5217
rect 9029 5149 9085 5183
rect 9029 5115 9040 5149
rect 9074 5115 9085 5149
rect 9029 5081 9085 5115
rect 9029 5047 9040 5081
rect 9074 5047 9085 5081
rect 9029 5013 9085 5047
rect 9029 4979 9040 5013
rect 9074 4979 9085 5013
rect 9029 4945 9085 4979
rect 9029 4911 9040 4945
rect 9074 4911 9085 4945
rect 9029 4877 9085 4911
rect 9029 4843 9040 4877
rect 9074 4843 9085 4877
rect 9029 4809 9085 4843
rect 9029 4775 9040 4809
rect 9074 4775 9085 4809
rect 9029 4741 9085 4775
rect 9029 4707 9040 4741
rect 9074 4707 9085 4741
rect 9029 4673 9085 4707
rect 9029 4639 9040 4673
rect 9074 4639 9085 4673
rect 9029 4605 9085 4639
rect 9029 4571 9040 4605
rect 9074 4571 9085 4605
rect 9029 4537 9085 4571
rect 9029 4503 9040 4537
rect 9074 4503 9085 4537
rect 9029 4469 9085 4503
rect 9029 4435 9040 4469
rect 9074 4435 9085 4469
rect 9029 4401 9085 4435
rect 9029 4367 9040 4401
rect 9074 4367 9085 4401
rect 9029 4333 9085 4367
rect 9029 4299 9040 4333
rect 9074 4299 9085 4333
rect 9029 4287 9085 4299
rect 9885 5489 9941 5523
rect 10741 5625 10794 5687
rect 10741 5591 10752 5625
rect 10786 5591 10794 5625
rect 10741 5557 10794 5591
rect 10741 5523 10752 5557
rect 10786 5523 10794 5557
rect 9885 5455 9896 5489
rect 9930 5455 9941 5489
rect 9885 5421 9941 5455
rect 9885 5387 9896 5421
rect 9930 5387 9941 5421
rect 9885 5353 9941 5387
rect 9885 5319 9896 5353
rect 9930 5319 9941 5353
rect 9885 5285 9941 5319
rect 9885 5251 9896 5285
rect 9930 5251 9941 5285
rect 9885 5217 9941 5251
rect 9885 5183 9896 5217
rect 9930 5183 9941 5217
rect 9885 5149 9941 5183
rect 9885 5115 9896 5149
rect 9930 5115 9941 5149
rect 9885 5081 9941 5115
rect 9885 5047 9896 5081
rect 9930 5047 9941 5081
rect 9885 5013 9941 5047
rect 9885 4979 9896 5013
rect 9930 4979 9941 5013
rect 9885 4945 9941 4979
rect 9885 4911 9896 4945
rect 9930 4911 9941 4945
rect 9885 4877 9941 4911
rect 9885 4843 9896 4877
rect 9930 4843 9941 4877
rect 9885 4809 9941 4843
rect 9885 4775 9896 4809
rect 9930 4775 9941 4809
rect 9885 4741 9941 4775
rect 9885 4707 9896 4741
rect 9930 4707 9941 4741
rect 9885 4673 9941 4707
rect 9885 4639 9896 4673
rect 9930 4639 9941 4673
rect 9885 4605 9941 4639
rect 9885 4571 9896 4605
rect 9930 4571 9941 4605
rect 9885 4537 9941 4571
rect 9885 4503 9896 4537
rect 9930 4503 9941 4537
rect 9885 4469 9941 4503
rect 9885 4435 9896 4469
rect 9930 4435 9941 4469
rect 9885 4401 9941 4435
rect 9885 4367 9896 4401
rect 9930 4367 9941 4401
rect 9885 4333 9941 4367
rect 9885 4299 9896 4333
rect 9930 4299 9941 4333
rect 9885 4287 9941 4299
rect 10741 5489 10794 5523
rect 10741 5455 10752 5489
rect 10786 5455 10794 5489
rect 10741 5421 10794 5455
rect 10741 5387 10752 5421
rect 10786 5387 10794 5421
rect 10741 5353 10794 5387
rect 10741 5319 10752 5353
rect 10786 5319 10794 5353
rect 10741 5285 10794 5319
rect 10741 5251 10752 5285
rect 10786 5251 10794 5285
rect 10741 5217 10794 5251
rect 10741 5183 10752 5217
rect 10786 5183 10794 5217
rect 10741 5149 10794 5183
rect 10741 5115 10752 5149
rect 10786 5115 10794 5149
rect 10741 5081 10794 5115
rect 10741 5047 10752 5081
rect 10786 5047 10794 5081
rect 10741 5013 10794 5047
rect 10741 4979 10752 5013
rect 10786 4979 10794 5013
rect 10741 4945 10794 4979
rect 10741 4911 10752 4945
rect 10786 4911 10794 4945
rect 10741 4877 10794 4911
rect 10741 4843 10752 4877
rect 10786 4843 10794 4877
rect 10741 4809 10794 4843
rect 10741 4775 10752 4809
rect 10786 4775 10794 4809
rect 10741 4741 10794 4775
rect 10741 4707 10752 4741
rect 10786 4707 10794 4741
rect 10741 4673 10794 4707
rect 10741 4639 10752 4673
rect 10786 4639 10794 4673
rect 10741 4605 10794 4639
rect 10741 4571 10752 4605
rect 10786 4571 10794 4605
rect 10741 4537 10794 4571
rect 10741 4503 10752 4537
rect 10786 4503 10794 4537
rect 10741 4469 10794 4503
rect 10741 4435 10752 4469
rect 10786 4435 10794 4469
rect 10741 4401 10794 4435
rect 10741 4367 10752 4401
rect 10786 4367 10794 4401
rect 10741 4333 10794 4367
rect 10741 4299 10752 4333
rect 10786 4299 10794 4333
rect 10741 4287 10794 4299
<< ndiffc >>
rect 480 7839 514 7873
rect 548 7839 582 7873
rect 3382 7839 3416 7873
rect 3450 7839 3484 7873
rect 12884 7839 12918 7873
rect 12952 7839 12986 7873
rect 480 7685 514 7719
rect 548 7685 582 7719
rect 3382 7685 3416 7719
rect 3450 7685 3484 7719
rect 12884 7685 12918 7719
rect 12952 7685 12986 7719
rect 480 7531 514 7565
rect 548 7531 582 7565
rect 3382 7531 3416 7565
rect 3450 7531 3484 7565
rect 12884 7531 12918 7565
rect 12952 7531 12986 7565
rect 480 7377 514 7411
rect 548 7377 582 7411
rect 3382 7377 3416 7411
rect 3450 7377 3484 7411
rect 12884 7377 12918 7411
rect 12952 7377 12986 7411
rect 480 7223 514 7257
rect 548 7223 582 7257
rect 3382 7223 3416 7257
rect 3450 7223 3484 7257
rect 12884 7223 12918 7257
rect 12952 7223 12986 7257
rect 480 7069 514 7103
rect 548 7069 582 7103
rect 3382 7069 3416 7103
rect 3450 7069 3484 7103
rect 12884 7069 12918 7103
rect 12952 7069 12986 7103
rect 480 6915 514 6949
rect 548 6915 582 6949
rect 3382 6915 3416 6949
rect 3450 6915 3484 6949
rect 12884 6915 12918 6949
rect 12952 6915 12986 6949
rect 480 6761 514 6795
rect 548 6761 582 6795
rect 3382 6761 3416 6795
rect 3450 6761 3484 6795
rect 12884 6761 12918 6795
rect 12952 6761 12986 6795
rect 480 6607 514 6641
rect 548 6607 582 6641
rect 3382 6607 3416 6641
rect 3450 6607 3484 6641
rect 12884 6607 12918 6641
rect 12952 6607 12986 6641
rect 480 6453 514 6487
rect 548 6453 582 6487
rect 3382 6453 3416 6487
rect 3450 6453 3484 6487
rect 12884 6453 12918 6487
rect 12952 6453 12986 6487
rect 480 6299 514 6333
rect 548 6299 582 6333
rect 3382 6299 3416 6333
rect 3450 6299 3484 6333
rect 12884 6299 12918 6333
rect 12952 6299 12986 6333
rect 480 6145 514 6179
rect 548 6145 582 6179
rect 3382 6145 3416 6179
rect 3450 6145 3484 6179
rect 12884 6145 12918 6179
rect 12952 6145 12986 6179
rect 11626 5854 11660 5888
rect 11694 5854 11728 5888
rect 14528 5854 14562 5888
rect 14596 5854 14630 5888
rect 11626 5700 11660 5734
rect 11694 5700 11728 5734
rect 14528 5700 14562 5734
rect 14596 5700 14630 5734
rect 11626 5546 11660 5580
rect 11694 5546 11728 5580
rect 14528 5546 14562 5580
rect 14596 5546 14630 5580
rect 11626 5392 11660 5426
rect 11694 5392 11728 5426
rect 14528 5392 14562 5426
rect 14596 5392 14630 5426
rect 11626 5238 11660 5272
rect 11694 5238 11728 5272
rect 14528 5238 14562 5272
rect 14596 5238 14630 5272
rect 11626 5084 11660 5118
rect 11694 5084 11728 5118
rect 14528 5084 14562 5118
rect 14596 5084 14630 5118
rect 11626 4930 11660 4964
rect 11694 4930 11728 4964
rect 14528 4930 14562 4964
rect 14596 4930 14630 4964
rect 11626 4776 11660 4810
rect 11694 4776 11728 4810
rect 14528 4776 14562 4810
rect 14596 4776 14630 4810
rect 11626 4622 11660 4656
rect 11694 4622 11728 4656
rect 14528 4622 14562 4656
rect 14596 4622 14630 4656
rect 11626 4468 11660 4502
rect 11694 4468 11728 4502
rect 14528 4468 14562 4502
rect 14596 4468 14630 4502
rect 11626 4314 11660 4348
rect 11694 4314 11728 4348
rect 14528 4314 14562 4348
rect 14596 4314 14630 4348
rect 11626 4160 11660 4194
rect 11694 4160 11728 4194
rect 14528 4160 14562 4194
rect 14596 4160 14630 4194
rect 11626 3874 11660 3908
rect 11694 3874 11728 3908
rect 14528 3874 14562 3908
rect 14596 3874 14630 3908
rect 11626 3720 11660 3754
rect 11694 3720 11728 3754
rect 14528 3720 14562 3754
rect 14596 3720 14630 3754
rect 11626 3566 11660 3600
rect 11694 3566 11728 3600
rect 14528 3566 14562 3600
rect 14596 3566 14630 3600
rect 11626 3412 11660 3446
rect 11694 3412 11728 3446
rect 14528 3412 14562 3446
rect 14596 3412 14630 3446
rect 11626 3258 11660 3292
rect 11694 3258 11728 3292
rect 14528 3258 14562 3292
rect 14596 3258 14630 3292
rect 11626 3104 11660 3138
rect 11694 3104 11728 3138
rect 14528 3104 14562 3138
rect 14596 3104 14630 3138
rect 11626 2950 11660 2984
rect 11694 2950 11728 2984
rect 14528 2950 14562 2984
rect 14596 2950 14630 2984
rect 11626 2796 11660 2830
rect 11694 2796 11728 2830
rect 14528 2796 14562 2830
rect 14596 2796 14630 2830
rect 11626 2642 11660 2676
rect 11694 2642 11728 2676
rect 14528 2642 14562 2676
rect 14596 2642 14630 2676
rect 11626 2488 11660 2522
rect 11694 2488 11728 2522
rect 14528 2488 14562 2522
rect 14596 2488 14630 2522
rect 11626 2334 11660 2368
rect 11694 2334 11728 2368
rect 14528 2334 14562 2368
rect 14596 2334 14630 2368
rect 11626 2180 11660 2214
rect 11694 2180 11728 2214
rect 14528 2180 14562 2214
rect 14596 2180 14630 2214
rect 480 1890 514 1924
rect 548 1890 582 1924
rect 3382 1890 3416 1924
rect 3450 1890 3484 1924
rect 12884 1890 12918 1924
rect 12952 1890 12986 1924
rect 480 1736 514 1770
rect 548 1736 582 1770
rect 3382 1736 3416 1770
rect 3450 1736 3484 1770
rect 12884 1736 12918 1770
rect 12952 1736 12986 1770
rect 480 1582 514 1616
rect 548 1582 582 1616
rect 3382 1582 3416 1616
rect 3450 1582 3484 1616
rect 12884 1582 12918 1616
rect 12952 1582 12986 1616
rect 480 1428 514 1462
rect 548 1428 582 1462
rect 3382 1428 3416 1462
rect 3450 1428 3484 1462
rect 12884 1428 12918 1462
rect 12952 1428 12986 1462
rect 480 1274 514 1308
rect 548 1274 582 1308
rect 3382 1274 3416 1308
rect 3450 1274 3484 1308
rect 12884 1274 12918 1308
rect 12952 1274 12986 1308
rect 480 1120 514 1154
rect 548 1120 582 1154
rect 3382 1120 3416 1154
rect 3450 1120 3484 1154
rect 12884 1120 12918 1154
rect 12952 1120 12986 1154
rect 480 966 514 1000
rect 548 966 582 1000
rect 3382 966 3416 1000
rect 3450 966 3484 1000
rect 12884 966 12918 1000
rect 12952 966 12986 1000
rect 480 812 514 846
rect 548 812 582 846
rect 3382 812 3416 846
rect 3450 812 3484 846
rect 12884 812 12918 846
rect 12952 812 12986 846
rect 480 658 514 692
rect 548 658 582 692
rect 3382 658 3416 692
rect 3450 658 3484 692
rect 12884 658 12918 692
rect 12952 658 12986 692
rect 480 504 514 538
rect 548 504 582 538
rect 3382 504 3416 538
rect 3450 504 3484 538
rect 12884 504 12918 538
rect 12952 504 12986 538
rect 480 350 514 384
rect 548 350 582 384
rect 3382 350 3416 384
rect 3450 350 3484 384
rect 12884 350 12918 384
rect 12952 350 12986 384
rect 480 196 514 230
rect 548 196 582 230
rect 3382 196 3416 230
rect 3450 196 3484 230
rect 12884 196 12918 230
rect 12952 196 12986 230
<< mvndiffc >>
rect 500 3625 534 3659
rect 500 3557 534 3591
rect 500 3489 534 3523
rect 500 3421 534 3455
rect 500 3353 534 3387
rect 500 3285 534 3319
rect 500 3217 534 3251
rect 500 3149 534 3183
rect 500 3081 534 3115
rect 500 3013 534 3047
rect 500 2945 534 2979
rect 500 2877 534 2911
rect 500 2809 534 2843
rect 500 2741 534 2775
rect 500 2673 534 2707
rect 500 2605 534 2639
rect 500 2537 534 2571
rect 500 2469 534 2503
rect 500 2401 534 2435
rect 500 2333 534 2367
rect 1356 3625 1390 3659
rect 1356 3557 1390 3591
rect 1356 3489 1390 3523
rect 1356 3421 1390 3455
rect 1356 3353 1390 3387
rect 1356 3285 1390 3319
rect 1356 3217 1390 3251
rect 1356 3149 1390 3183
rect 1356 3081 1390 3115
rect 1356 3013 1390 3047
rect 1356 2945 1390 2979
rect 1356 2877 1390 2911
rect 1356 2809 1390 2843
rect 1356 2741 1390 2775
rect 1356 2673 1390 2707
rect 1356 2605 1390 2639
rect 1356 2537 1390 2571
rect 1356 2469 1390 2503
rect 1356 2401 1390 2435
rect 1356 2333 1390 2367
rect 2212 3625 2246 3659
rect 2212 3557 2246 3591
rect 2212 3489 2246 3523
rect 2212 3421 2246 3455
rect 2212 3353 2246 3387
rect 2212 3285 2246 3319
rect 2212 3217 2246 3251
rect 2212 3149 2246 3183
rect 2212 3081 2246 3115
rect 2212 3013 2246 3047
rect 2212 2945 2246 2979
rect 2212 2877 2246 2911
rect 2212 2809 2246 2843
rect 2212 2741 2246 2775
rect 2212 2673 2246 2707
rect 2212 2605 2246 2639
rect 2212 2537 2246 2571
rect 2212 2469 2246 2503
rect 2212 2401 2246 2435
rect 2212 2333 2246 2367
rect 3068 3625 3102 3659
rect 3068 3557 3102 3591
rect 3068 3489 3102 3523
rect 3068 3421 3102 3455
rect 3068 3353 3102 3387
rect 3068 3285 3102 3319
rect 3068 3217 3102 3251
rect 3068 3149 3102 3183
rect 3068 3081 3102 3115
rect 3068 3013 3102 3047
rect 3068 2945 3102 2979
rect 3068 2877 3102 2911
rect 3068 2809 3102 2843
rect 3068 2741 3102 2775
rect 3068 2673 3102 2707
rect 3068 2605 3102 2639
rect 3068 2537 3102 2571
rect 3068 2469 3102 2503
rect 3068 2401 3102 2435
rect 3068 2333 3102 2367
rect 3924 3625 3958 3659
rect 3924 3557 3958 3591
rect 3924 3489 3958 3523
rect 3924 3421 3958 3455
rect 3924 3353 3958 3387
rect 3924 3285 3958 3319
rect 3924 3217 3958 3251
rect 3924 3149 3958 3183
rect 3924 3081 3958 3115
rect 3924 3013 3958 3047
rect 3924 2945 3958 2979
rect 3924 2877 3958 2911
rect 3924 2809 3958 2843
rect 3924 2741 3958 2775
rect 3924 2673 3958 2707
rect 3924 2605 3958 2639
rect 3924 2537 3958 2571
rect 3924 2469 3958 2503
rect 3924 2401 3958 2435
rect 3924 2333 3958 2367
rect 4780 3625 4814 3659
rect 4780 3557 4814 3591
rect 4780 3489 4814 3523
rect 4780 3421 4814 3455
rect 4780 3353 4814 3387
rect 4780 3285 4814 3319
rect 4780 3217 4814 3251
rect 4780 3149 4814 3183
rect 4780 3081 4814 3115
rect 4780 3013 4814 3047
rect 4780 2945 4814 2979
rect 4780 2877 4814 2911
rect 4780 2809 4814 2843
rect 4780 2741 4814 2775
rect 4780 2673 4814 2707
rect 4780 2605 4814 2639
rect 4780 2537 4814 2571
rect 4780 2469 4814 2503
rect 4780 2401 4814 2435
rect 4780 2333 4814 2367
rect 5636 3625 5670 3659
rect 5636 3557 5670 3591
rect 5636 3489 5670 3523
rect 5636 3421 5670 3455
rect 5636 3353 5670 3387
rect 5636 3285 5670 3319
rect 5636 3217 5670 3251
rect 5636 3149 5670 3183
rect 5636 3081 5670 3115
rect 5636 3013 5670 3047
rect 5636 2945 5670 2979
rect 5636 2877 5670 2911
rect 5636 2809 5670 2843
rect 5636 2741 5670 2775
rect 5636 2673 5670 2707
rect 5636 2605 5670 2639
rect 5636 2537 5670 2571
rect 5636 2469 5670 2503
rect 5636 2401 5670 2435
rect 5636 2333 5670 2367
rect 6492 3625 6526 3659
rect 6492 3557 6526 3591
rect 6492 3489 6526 3523
rect 6492 3421 6526 3455
rect 6492 3353 6526 3387
rect 6492 3285 6526 3319
rect 6492 3217 6526 3251
rect 6492 3149 6526 3183
rect 6492 3081 6526 3115
rect 6492 3013 6526 3047
rect 6492 2945 6526 2979
rect 6492 2877 6526 2911
rect 6492 2809 6526 2843
rect 6492 2741 6526 2775
rect 6492 2673 6526 2707
rect 6492 2605 6526 2639
rect 6492 2537 6526 2571
rect 6492 2469 6526 2503
rect 6492 2401 6526 2435
rect 6492 2333 6526 2367
rect 7348 3625 7382 3659
rect 7348 3557 7382 3591
rect 7348 3489 7382 3523
rect 7348 3421 7382 3455
rect 7348 3353 7382 3387
rect 7348 3285 7382 3319
rect 7348 3217 7382 3251
rect 7348 3149 7382 3183
rect 7348 3081 7382 3115
rect 7348 3013 7382 3047
rect 7348 2945 7382 2979
rect 7348 2877 7382 2911
rect 7348 2809 7382 2843
rect 7348 2741 7382 2775
rect 7348 2673 7382 2707
rect 7348 2605 7382 2639
rect 7348 2537 7382 2571
rect 7348 2469 7382 2503
rect 7348 2401 7382 2435
rect 7348 2333 7382 2367
rect 8204 3625 8238 3659
rect 8204 3557 8238 3591
rect 8204 3489 8238 3523
rect 8204 3421 8238 3455
rect 8204 3353 8238 3387
rect 8204 3285 8238 3319
rect 8204 3217 8238 3251
rect 8204 3149 8238 3183
rect 8204 3081 8238 3115
rect 8204 3013 8238 3047
rect 8204 2945 8238 2979
rect 8204 2877 8238 2911
rect 8204 2809 8238 2843
rect 8204 2741 8238 2775
rect 8204 2673 8238 2707
rect 8204 2605 8238 2639
rect 8204 2537 8238 2571
rect 8204 2469 8238 2503
rect 8204 2401 8238 2435
rect 8204 2333 8238 2367
rect 9060 3625 9094 3659
rect 9060 3557 9094 3591
rect 9060 3489 9094 3523
rect 9060 3421 9094 3455
rect 9060 3353 9094 3387
rect 9060 3285 9094 3319
rect 9060 3217 9094 3251
rect 9060 3149 9094 3183
rect 9060 3081 9094 3115
rect 9060 3013 9094 3047
rect 9060 2945 9094 2979
rect 9060 2877 9094 2911
rect 9060 2809 9094 2843
rect 9060 2741 9094 2775
rect 9060 2673 9094 2707
rect 9060 2605 9094 2639
rect 9060 2537 9094 2571
rect 9060 2469 9094 2503
rect 9060 2401 9094 2435
rect 9060 2333 9094 2367
rect 9916 3625 9950 3659
rect 9916 3557 9950 3591
rect 9916 3489 9950 3523
rect 9916 3421 9950 3455
rect 9916 3353 9950 3387
rect 9916 3285 9950 3319
rect 9916 3217 9950 3251
rect 9916 3149 9950 3183
rect 9916 3081 9950 3115
rect 9916 3013 9950 3047
rect 9916 2945 9950 2979
rect 9916 2877 9950 2911
rect 9916 2809 9950 2843
rect 9916 2741 9950 2775
rect 9916 2673 9950 2707
rect 9916 2605 9950 2639
rect 9916 2537 9950 2571
rect 9916 2469 9950 2503
rect 9916 2401 9950 2435
rect 9916 2333 9950 2367
rect 10772 3625 10806 3659
rect 10772 3557 10806 3591
rect 10772 3489 10806 3523
rect 10772 3421 10806 3455
rect 10772 3353 10806 3387
rect 10772 3285 10806 3319
rect 10772 3217 10806 3251
rect 10772 3149 10806 3183
rect 10772 3081 10806 3115
rect 10772 3013 10806 3047
rect 10772 2945 10806 2979
rect 10772 2877 10806 2911
rect 10772 2809 10806 2843
rect 10772 2741 10806 2775
rect 10772 2673 10806 2707
rect 10772 2605 10806 2639
rect 10772 2537 10806 2571
rect 10772 2469 10806 2503
rect 10772 2401 10806 2435
rect 10772 2333 10806 2367
<< mvpdiffc >>
rect 480 5591 514 5625
rect 480 5523 514 5557
rect 1336 5591 1370 5625
rect 1336 5523 1370 5557
rect 480 5455 514 5489
rect 480 5387 514 5421
rect 480 5319 514 5353
rect 480 5251 514 5285
rect 480 5183 514 5217
rect 480 5115 514 5149
rect 480 5047 514 5081
rect 480 4979 514 5013
rect 480 4911 514 4945
rect 480 4843 514 4877
rect 480 4775 514 4809
rect 480 4707 514 4741
rect 480 4639 514 4673
rect 480 4571 514 4605
rect 480 4503 514 4537
rect 480 4435 514 4469
rect 480 4367 514 4401
rect 480 4299 514 4333
rect 2192 5591 2226 5625
rect 2192 5523 2226 5557
rect 1336 5455 1370 5489
rect 1336 5387 1370 5421
rect 1336 5319 1370 5353
rect 1336 5251 1370 5285
rect 1336 5183 1370 5217
rect 1336 5115 1370 5149
rect 1336 5047 1370 5081
rect 1336 4979 1370 5013
rect 1336 4911 1370 4945
rect 1336 4843 1370 4877
rect 1336 4775 1370 4809
rect 1336 4707 1370 4741
rect 1336 4639 1370 4673
rect 1336 4571 1370 4605
rect 1336 4503 1370 4537
rect 1336 4435 1370 4469
rect 1336 4367 1370 4401
rect 1336 4299 1370 4333
rect 3048 5591 3082 5625
rect 3048 5523 3082 5557
rect 2192 5455 2226 5489
rect 2192 5387 2226 5421
rect 2192 5319 2226 5353
rect 2192 5251 2226 5285
rect 2192 5183 2226 5217
rect 2192 5115 2226 5149
rect 2192 5047 2226 5081
rect 2192 4979 2226 5013
rect 2192 4911 2226 4945
rect 2192 4843 2226 4877
rect 2192 4775 2226 4809
rect 2192 4707 2226 4741
rect 2192 4639 2226 4673
rect 2192 4571 2226 4605
rect 2192 4503 2226 4537
rect 2192 4435 2226 4469
rect 2192 4367 2226 4401
rect 2192 4299 2226 4333
rect 3904 5591 3938 5625
rect 3904 5523 3938 5557
rect 3048 5455 3082 5489
rect 3048 5387 3082 5421
rect 3048 5319 3082 5353
rect 3048 5251 3082 5285
rect 3048 5183 3082 5217
rect 3048 5115 3082 5149
rect 3048 5047 3082 5081
rect 3048 4979 3082 5013
rect 3048 4911 3082 4945
rect 3048 4843 3082 4877
rect 3048 4775 3082 4809
rect 3048 4707 3082 4741
rect 3048 4639 3082 4673
rect 3048 4571 3082 4605
rect 3048 4503 3082 4537
rect 3048 4435 3082 4469
rect 3048 4367 3082 4401
rect 3048 4299 3082 4333
rect 4760 5591 4794 5625
rect 4760 5523 4794 5557
rect 3904 5455 3938 5489
rect 3904 5387 3938 5421
rect 3904 5319 3938 5353
rect 3904 5251 3938 5285
rect 3904 5183 3938 5217
rect 3904 5115 3938 5149
rect 3904 5047 3938 5081
rect 3904 4979 3938 5013
rect 3904 4911 3938 4945
rect 3904 4843 3938 4877
rect 3904 4775 3938 4809
rect 3904 4707 3938 4741
rect 3904 4639 3938 4673
rect 3904 4571 3938 4605
rect 3904 4503 3938 4537
rect 3904 4435 3938 4469
rect 3904 4367 3938 4401
rect 3904 4299 3938 4333
rect 5616 5591 5650 5625
rect 5616 5523 5650 5557
rect 4760 5455 4794 5489
rect 4760 5387 4794 5421
rect 4760 5319 4794 5353
rect 4760 5251 4794 5285
rect 4760 5183 4794 5217
rect 4760 5115 4794 5149
rect 4760 5047 4794 5081
rect 4760 4979 4794 5013
rect 4760 4911 4794 4945
rect 4760 4843 4794 4877
rect 4760 4775 4794 4809
rect 4760 4707 4794 4741
rect 4760 4639 4794 4673
rect 4760 4571 4794 4605
rect 4760 4503 4794 4537
rect 4760 4435 4794 4469
rect 4760 4367 4794 4401
rect 4760 4299 4794 4333
rect 6472 5591 6506 5625
rect 6472 5523 6506 5557
rect 5616 5455 5650 5489
rect 5616 5387 5650 5421
rect 5616 5319 5650 5353
rect 5616 5251 5650 5285
rect 5616 5183 5650 5217
rect 5616 5115 5650 5149
rect 5616 5047 5650 5081
rect 5616 4979 5650 5013
rect 5616 4911 5650 4945
rect 5616 4843 5650 4877
rect 5616 4775 5650 4809
rect 5616 4707 5650 4741
rect 5616 4639 5650 4673
rect 5616 4571 5650 4605
rect 5616 4503 5650 4537
rect 5616 4435 5650 4469
rect 5616 4367 5650 4401
rect 5616 4299 5650 4333
rect 7328 5591 7362 5625
rect 7328 5523 7362 5557
rect 6472 5455 6506 5489
rect 6472 5387 6506 5421
rect 6472 5319 6506 5353
rect 6472 5251 6506 5285
rect 6472 5183 6506 5217
rect 6472 5115 6506 5149
rect 6472 5047 6506 5081
rect 6472 4979 6506 5013
rect 6472 4911 6506 4945
rect 6472 4843 6506 4877
rect 6472 4775 6506 4809
rect 6472 4707 6506 4741
rect 6472 4639 6506 4673
rect 6472 4571 6506 4605
rect 6472 4503 6506 4537
rect 6472 4435 6506 4469
rect 6472 4367 6506 4401
rect 6472 4299 6506 4333
rect 8184 5591 8218 5625
rect 8184 5523 8218 5557
rect 7328 5455 7362 5489
rect 7328 5387 7362 5421
rect 7328 5319 7362 5353
rect 7328 5251 7362 5285
rect 7328 5183 7362 5217
rect 7328 5115 7362 5149
rect 7328 5047 7362 5081
rect 7328 4979 7362 5013
rect 7328 4911 7362 4945
rect 7328 4843 7362 4877
rect 7328 4775 7362 4809
rect 7328 4707 7362 4741
rect 7328 4639 7362 4673
rect 7328 4571 7362 4605
rect 7328 4503 7362 4537
rect 7328 4435 7362 4469
rect 7328 4367 7362 4401
rect 7328 4299 7362 4333
rect 9040 5591 9074 5625
rect 9040 5523 9074 5557
rect 8184 5455 8218 5489
rect 8184 5387 8218 5421
rect 8184 5319 8218 5353
rect 8184 5251 8218 5285
rect 8184 5183 8218 5217
rect 8184 5115 8218 5149
rect 8184 5047 8218 5081
rect 8184 4979 8218 5013
rect 8184 4911 8218 4945
rect 8184 4843 8218 4877
rect 8184 4775 8218 4809
rect 8184 4707 8218 4741
rect 8184 4639 8218 4673
rect 8184 4571 8218 4605
rect 8184 4503 8218 4537
rect 8184 4435 8218 4469
rect 8184 4367 8218 4401
rect 8184 4299 8218 4333
rect 9896 5591 9930 5625
rect 9896 5523 9930 5557
rect 9040 5455 9074 5489
rect 9040 5387 9074 5421
rect 9040 5319 9074 5353
rect 9040 5251 9074 5285
rect 9040 5183 9074 5217
rect 9040 5115 9074 5149
rect 9040 5047 9074 5081
rect 9040 4979 9074 5013
rect 9040 4911 9074 4945
rect 9040 4843 9074 4877
rect 9040 4775 9074 4809
rect 9040 4707 9074 4741
rect 9040 4639 9074 4673
rect 9040 4571 9074 4605
rect 9040 4503 9074 4537
rect 9040 4435 9074 4469
rect 9040 4367 9074 4401
rect 9040 4299 9074 4333
rect 10752 5591 10786 5625
rect 10752 5523 10786 5557
rect 9896 5455 9930 5489
rect 9896 5387 9930 5421
rect 9896 5319 9930 5353
rect 9896 5251 9930 5285
rect 9896 5183 9930 5217
rect 9896 5115 9930 5149
rect 9896 5047 9930 5081
rect 9896 4979 9930 5013
rect 9896 4911 9930 4945
rect 9896 4843 9930 4877
rect 9896 4775 9930 4809
rect 9896 4707 9930 4741
rect 9896 4639 9930 4673
rect 9896 4571 9930 4605
rect 9896 4503 9930 4537
rect 9896 4435 9930 4469
rect 9896 4367 9930 4401
rect 9896 4299 9930 4333
rect 10752 5455 10786 5489
rect 10752 5387 10786 5421
rect 10752 5319 10786 5353
rect 10752 5251 10786 5285
rect 10752 5183 10786 5217
rect 10752 5115 10786 5149
rect 10752 5047 10786 5081
rect 10752 4979 10786 5013
rect 10752 4911 10786 4945
rect 10752 4843 10786 4877
rect 10752 4775 10786 4809
rect 10752 4707 10786 4741
rect 10752 4639 10786 4673
rect 10752 4571 10786 4605
rect 10752 4503 10786 4537
rect 10752 4435 10786 4469
rect 10752 4367 10786 4401
rect 10752 4299 10786 4333
<< psubdiff >>
rect 336 8018 16032 8042
rect 370 7984 405 8018
rect 439 7984 474 8018
rect 508 7984 543 8018
rect 577 7984 612 8018
rect 646 7984 681 8018
rect 715 7984 750 8018
rect 784 7984 819 8018
rect 853 7984 888 8018
rect 922 7984 957 8018
rect 991 7984 1026 8018
rect 1060 7984 1095 8018
rect 1129 7984 1164 8018
rect 1198 7984 1233 8018
rect 1267 7984 1302 8018
rect 1336 7984 1371 8018
rect 1405 7984 1440 8018
rect 1474 7984 1509 8018
rect 1543 7984 1578 8018
rect 1612 7984 1647 8018
rect 1681 7984 1716 8018
rect 1750 7984 1784 8018
rect 1818 7984 1852 8018
rect 1886 7984 1920 8018
rect 1954 7984 1988 8018
rect 2022 7984 2056 8018
rect 2090 7984 2124 8018
rect 2158 7984 2192 8018
rect 2226 7984 2260 8018
rect 2294 7984 2328 8018
rect 2362 7984 2396 8018
rect 2430 7984 2464 8018
rect 2498 7984 2532 8018
rect 2566 7984 2600 8018
rect 2634 7984 2668 8018
rect 2702 7984 2736 8018
rect 2770 7984 2804 8018
rect 2838 7984 2872 8018
rect 2906 7984 2940 8018
rect 2974 7984 3008 8018
rect 3042 7984 3076 8018
rect 3110 7984 3144 8018
rect 3178 7984 3212 8018
rect 3246 7984 3280 8018
rect 3314 7984 3348 8018
rect 3382 7984 3416 8018
rect 3450 7984 3484 8018
rect 3518 7984 3552 8018
rect 3586 7984 3620 8018
rect 3654 7984 3688 8018
rect 3722 7984 3756 8018
rect 3790 7984 3824 8018
rect 3858 7984 3892 8018
rect 3926 7984 3960 8018
rect 3994 7984 4028 8018
rect 4062 7984 4096 8018
rect 4130 7984 4164 8018
rect 4198 7984 4232 8018
rect 4266 7984 4300 8018
rect 4334 7984 4368 8018
rect 4402 7984 4436 8018
rect 4470 7984 4504 8018
rect 4538 7984 4572 8018
rect 4606 7984 4640 8018
rect 4674 7984 4708 8018
rect 4742 7984 4776 8018
rect 4810 7984 4844 8018
rect 4878 7984 4912 8018
rect 4946 7984 4980 8018
rect 5014 7984 5048 8018
rect 5082 7984 5116 8018
rect 5150 7984 5184 8018
rect 5218 7984 5252 8018
rect 5286 7984 5320 8018
rect 5354 7984 5388 8018
rect 5422 7984 5456 8018
rect 5490 7984 5524 8018
rect 5558 7984 5592 8018
rect 5626 7984 5660 8018
rect 5694 7984 5728 8018
rect 5762 7984 5796 8018
rect 5830 7984 5864 8018
rect 5898 7984 5932 8018
rect 5966 7984 6000 8018
rect 6034 7984 6068 8018
rect 6102 7984 6136 8018
rect 6170 7984 6204 8018
rect 6238 7984 6272 8018
rect 6306 7984 6340 8018
rect 6374 7984 6408 8018
rect 6442 7984 6476 8018
rect 6510 7984 6544 8018
rect 6578 7984 6612 8018
rect 6646 7984 6680 8018
rect 6714 7984 6748 8018
rect 6782 7984 6816 8018
rect 6850 7984 6884 8018
rect 6918 7984 6952 8018
rect 6986 7984 7020 8018
rect 7054 7984 7088 8018
rect 7122 7984 7156 8018
rect 7190 7984 7224 8018
rect 7258 7984 7292 8018
rect 7326 7984 7360 8018
rect 7394 7984 7428 8018
rect 7462 7984 7496 8018
rect 7530 7984 7564 8018
rect 7598 7984 7632 8018
rect 7666 7984 7700 8018
rect 7734 7984 7768 8018
rect 7802 7984 7836 8018
rect 7870 7984 7904 8018
rect 7938 7984 7972 8018
rect 8006 7984 8040 8018
rect 8074 7984 8108 8018
rect 8142 7984 8176 8018
rect 8210 7984 8244 8018
rect 8278 7984 8312 8018
rect 8346 7984 8380 8018
rect 8414 7984 8448 8018
rect 8482 7984 8516 8018
rect 8550 7984 8584 8018
rect 8618 7984 8652 8018
rect 8686 7984 8720 8018
rect 8754 7984 8788 8018
rect 8822 7984 8856 8018
rect 8890 7984 8924 8018
rect 8958 7984 8992 8018
rect 9026 7984 9060 8018
rect 9094 7984 9128 8018
rect 9162 7984 9196 8018
rect 9230 7984 9264 8018
rect 9298 7984 9332 8018
rect 9366 7984 9400 8018
rect 9434 7984 9468 8018
rect 9502 7984 9536 8018
rect 9570 7984 9604 8018
rect 9638 7984 9672 8018
rect 9706 7984 9740 8018
rect 9774 7984 9808 8018
rect 9842 7984 9876 8018
rect 9910 7984 9944 8018
rect 9978 7984 10012 8018
rect 10046 7984 10080 8018
rect 10114 7984 10148 8018
rect 10182 7984 10216 8018
rect 10250 7984 10284 8018
rect 10318 7984 10352 8018
rect 10386 7984 10420 8018
rect 10454 7984 10488 8018
rect 10522 7984 10556 8018
rect 10590 7984 10624 8018
rect 10658 7984 10692 8018
rect 10726 7984 10760 8018
rect 10794 7984 10828 8018
rect 10862 7984 10896 8018
rect 10930 7984 10964 8018
rect 10998 7984 11032 8018
rect 11066 7984 11100 8018
rect 11134 7984 11168 8018
rect 11202 7984 11236 8018
rect 11270 7984 11304 8018
rect 11338 7984 11372 8018
rect 11406 7984 11440 8018
rect 11474 7984 11508 8018
rect 11542 7984 11576 8018
rect 11610 7984 11644 8018
rect 11678 7984 11712 8018
rect 11746 7984 11780 8018
rect 11814 7984 11848 8018
rect 11882 7984 11916 8018
rect 11950 7984 11984 8018
rect 12018 7984 12052 8018
rect 12086 7984 12120 8018
rect 12154 7984 12188 8018
rect 12222 7984 12256 8018
rect 12290 7984 12324 8018
rect 12358 7984 12392 8018
rect 12426 7984 12460 8018
rect 12494 7984 12528 8018
rect 12562 7984 12596 8018
rect 12630 7984 12664 8018
rect 12698 7984 12732 8018
rect 12766 7984 12800 8018
rect 12834 7984 12868 8018
rect 12902 7984 12936 8018
rect 12970 7984 13004 8018
rect 13038 7984 13072 8018
rect 13106 7984 13140 8018
rect 13174 7984 13208 8018
rect 13242 7984 13276 8018
rect 13310 7984 13344 8018
rect 13378 7984 13412 8018
rect 13446 7984 13480 8018
rect 13514 7984 13548 8018
rect 13582 7984 13616 8018
rect 13650 7984 13684 8018
rect 13718 7984 13752 8018
rect 13786 7984 13820 8018
rect 13854 7984 13888 8018
rect 13922 7984 13956 8018
rect 13990 7984 14024 8018
rect 14058 7984 14092 8018
rect 14126 7984 14160 8018
rect 14194 7984 14228 8018
rect 14262 7984 14296 8018
rect 14330 7984 14364 8018
rect 14398 7984 14432 8018
rect 14466 7984 14500 8018
rect 14534 7984 14568 8018
rect 14602 7984 14636 8018
rect 14670 7984 14774 8018
rect 14808 7984 14844 8018
rect 14878 7984 14914 8018
rect 14948 7984 14984 8018
rect 15018 7984 15054 8018
rect 15088 7984 15124 8018
rect 15158 7984 15194 8018
rect 15228 7984 15264 8018
rect 15298 7984 15334 8018
rect 15368 7984 15404 8018
rect 15438 7984 15474 8018
rect 15508 7984 15544 8018
rect 15578 7984 15614 8018
rect 15648 7984 15684 8018
rect 15718 7984 15754 8018
rect 15788 7984 15824 8018
rect 15858 7984 15894 8018
rect 15928 7984 15964 8018
rect 15998 7984 16032 8018
rect 336 7960 16032 7984
rect 336 7908 418 7960
rect 336 7874 360 7908
rect 394 7874 418 7908
rect 13152 7949 16032 7960
rect 13152 7928 14774 7949
rect 336 7838 418 7874
rect 336 7804 360 7838
rect 394 7804 418 7838
rect 13152 7894 13194 7928
rect 13228 7894 13264 7928
rect 13298 7894 13334 7928
rect 13368 7894 13404 7928
rect 13438 7894 13474 7928
rect 13508 7894 13544 7928
rect 13578 7894 13614 7928
rect 13648 7894 13684 7928
rect 13718 7894 13754 7928
rect 13788 7894 13824 7928
rect 13858 7894 13894 7928
rect 13928 7894 13964 7928
rect 13998 7894 14034 7928
rect 14068 7894 14104 7928
rect 14138 7894 14174 7928
rect 14208 7894 14244 7928
rect 14278 7894 14314 7928
rect 14348 7894 14384 7928
rect 14418 7894 14454 7928
rect 14488 7894 14524 7928
rect 14558 7894 14594 7928
rect 14628 7894 14664 7928
rect 14698 7915 14774 7928
rect 14808 7915 14844 7949
rect 14878 7915 14914 7949
rect 14948 7915 14984 7949
rect 15018 7915 15054 7949
rect 15088 7915 15124 7949
rect 15158 7915 15194 7949
rect 15228 7915 15264 7949
rect 15298 7915 15334 7949
rect 15368 7915 15404 7949
rect 15438 7915 15474 7949
rect 15508 7915 15544 7949
rect 15578 7915 15614 7949
rect 15648 7915 15684 7949
rect 15718 7915 15754 7949
rect 15788 7915 15824 7949
rect 15858 7915 15894 7949
rect 15928 7915 15964 7949
rect 15998 7915 16032 7949
rect 14698 7894 16032 7915
rect 13152 7880 16032 7894
rect 13152 7858 14774 7880
rect 13152 7824 13194 7858
rect 13228 7824 13264 7858
rect 13298 7824 13334 7858
rect 13368 7824 13404 7858
rect 13438 7824 13474 7858
rect 13508 7824 13544 7858
rect 13578 7824 13614 7858
rect 13648 7824 13684 7858
rect 13718 7824 13754 7858
rect 13788 7824 13824 7858
rect 13858 7824 13894 7858
rect 13928 7824 13964 7858
rect 13998 7824 14034 7858
rect 14068 7824 14104 7858
rect 14138 7824 14174 7858
rect 14208 7824 14244 7858
rect 14278 7824 14314 7858
rect 14348 7824 14384 7858
rect 14418 7824 14454 7858
rect 14488 7824 14524 7858
rect 14558 7824 14594 7858
rect 14628 7824 14664 7858
rect 14698 7846 14774 7858
rect 14808 7846 14844 7880
rect 14878 7846 14914 7880
rect 14948 7846 14984 7880
rect 15018 7846 15054 7880
rect 15088 7846 15124 7880
rect 15158 7846 15194 7880
rect 15228 7846 15264 7880
rect 15298 7846 15334 7880
rect 15368 7846 15404 7880
rect 15438 7846 15474 7880
rect 15508 7846 15544 7880
rect 15578 7846 15614 7880
rect 15648 7846 15684 7880
rect 15718 7846 15754 7880
rect 15788 7846 15824 7880
rect 15858 7846 15894 7880
rect 15928 7846 15964 7880
rect 15998 7846 16032 7880
rect 14698 7824 16032 7846
rect 13152 7811 16032 7824
rect 336 7768 418 7804
rect 336 7734 360 7768
rect 394 7734 418 7768
rect 13152 7788 14774 7811
rect 13152 7754 13194 7788
rect 13228 7754 13264 7788
rect 13298 7754 13334 7788
rect 13368 7754 13404 7788
rect 13438 7754 13474 7788
rect 13508 7754 13544 7788
rect 13578 7754 13614 7788
rect 13648 7754 13684 7788
rect 13718 7754 13754 7788
rect 13788 7754 13824 7788
rect 13858 7754 13894 7788
rect 13928 7754 13964 7788
rect 13998 7754 14034 7788
rect 14068 7754 14104 7788
rect 14138 7754 14174 7788
rect 14208 7754 14244 7788
rect 14278 7754 14314 7788
rect 14348 7754 14384 7788
rect 14418 7754 14454 7788
rect 14488 7754 14524 7788
rect 14558 7754 14594 7788
rect 14628 7754 14664 7788
rect 14698 7777 14774 7788
rect 14808 7777 14844 7811
rect 14878 7777 14914 7811
rect 14948 7777 14984 7811
rect 15018 7777 15054 7811
rect 15088 7777 15124 7811
rect 15158 7777 15194 7811
rect 15228 7777 15264 7811
rect 15298 7777 15334 7811
rect 15368 7777 15404 7811
rect 15438 7777 15474 7811
rect 15508 7777 15544 7811
rect 15578 7777 15614 7811
rect 15648 7777 15684 7811
rect 15718 7777 15754 7811
rect 15788 7777 15824 7811
rect 15858 7777 15894 7811
rect 15928 7777 15964 7811
rect 15998 7777 16032 7811
rect 14698 7754 16032 7777
rect 336 7698 418 7734
rect 336 7664 360 7698
rect 394 7664 418 7698
rect 336 7628 418 7664
rect 13152 7742 16032 7754
rect 13152 7718 14774 7742
rect 13152 7684 13194 7718
rect 13228 7684 13264 7718
rect 13298 7684 13334 7718
rect 13368 7684 13404 7718
rect 13438 7684 13474 7718
rect 13508 7684 13544 7718
rect 13578 7684 13614 7718
rect 13648 7684 13684 7718
rect 13718 7684 13754 7718
rect 13788 7684 13824 7718
rect 13858 7684 13894 7718
rect 13928 7684 13964 7718
rect 13998 7684 14034 7718
rect 14068 7684 14104 7718
rect 14138 7684 14174 7718
rect 14208 7684 14244 7718
rect 14278 7684 14314 7718
rect 14348 7684 14384 7718
rect 14418 7684 14454 7718
rect 14488 7684 14524 7718
rect 14558 7684 14594 7718
rect 14628 7684 14664 7718
rect 14698 7708 14774 7718
rect 14808 7708 14844 7742
rect 14878 7708 14914 7742
rect 14948 7708 14984 7742
rect 15018 7708 15054 7742
rect 15088 7708 15124 7742
rect 15158 7708 15194 7742
rect 15228 7708 15264 7742
rect 15298 7708 15334 7742
rect 15368 7708 15404 7742
rect 15438 7708 15474 7742
rect 15508 7708 15544 7742
rect 15578 7708 15614 7742
rect 15648 7708 15684 7742
rect 15718 7708 15754 7742
rect 15788 7708 15824 7742
rect 15858 7708 15894 7742
rect 15928 7708 15964 7742
rect 15998 7708 16032 7742
rect 14698 7684 16032 7708
rect 13152 7673 16032 7684
rect 336 7594 360 7628
rect 394 7594 418 7628
rect 13152 7648 14774 7673
rect 13152 7614 13194 7648
rect 13228 7614 13264 7648
rect 13298 7614 13334 7648
rect 13368 7614 13404 7648
rect 13438 7614 13474 7648
rect 13508 7614 13544 7648
rect 13578 7614 13614 7648
rect 13648 7614 13684 7648
rect 13718 7614 13754 7648
rect 13788 7614 13824 7648
rect 13858 7614 13894 7648
rect 13928 7614 13964 7648
rect 13998 7614 14034 7648
rect 14068 7614 14104 7648
rect 14138 7614 14174 7648
rect 14208 7614 14244 7648
rect 14278 7614 14314 7648
rect 14348 7614 14384 7648
rect 14418 7614 14454 7648
rect 14488 7614 14524 7648
rect 14558 7614 14594 7648
rect 14628 7614 14664 7648
rect 14698 7639 14774 7648
rect 14808 7639 14844 7673
rect 14878 7639 14914 7673
rect 14948 7639 14984 7673
rect 15018 7639 15054 7673
rect 15088 7639 15124 7673
rect 15158 7639 15194 7673
rect 15228 7639 15264 7673
rect 15298 7639 15334 7673
rect 15368 7639 15404 7673
rect 15438 7639 15474 7673
rect 15508 7639 15544 7673
rect 15578 7639 15614 7673
rect 15648 7639 15684 7673
rect 15718 7639 15754 7673
rect 15788 7639 15824 7673
rect 15858 7639 15894 7673
rect 15928 7639 15964 7673
rect 15998 7639 16032 7673
rect 14698 7614 16032 7639
rect 13152 7604 16032 7614
rect 336 7558 418 7594
rect 336 7524 360 7558
rect 394 7524 418 7558
rect 336 7488 418 7524
rect 13152 7578 14774 7604
rect 13152 7544 13194 7578
rect 13228 7544 13264 7578
rect 13298 7544 13334 7578
rect 13368 7544 13404 7578
rect 13438 7544 13474 7578
rect 13508 7544 13544 7578
rect 13578 7544 13614 7578
rect 13648 7544 13684 7578
rect 13718 7544 13754 7578
rect 13788 7544 13824 7578
rect 13858 7544 13894 7578
rect 13928 7544 13964 7578
rect 13998 7544 14034 7578
rect 14068 7544 14104 7578
rect 14138 7544 14174 7578
rect 14208 7544 14244 7578
rect 14278 7544 14314 7578
rect 14348 7544 14384 7578
rect 14418 7544 14454 7578
rect 14488 7544 14524 7578
rect 14558 7544 14594 7578
rect 14628 7544 14664 7578
rect 14698 7570 14774 7578
rect 14808 7570 14844 7604
rect 14878 7570 14914 7604
rect 14948 7570 14984 7604
rect 15018 7570 15054 7604
rect 15088 7570 15124 7604
rect 15158 7570 15194 7604
rect 15228 7570 15264 7604
rect 15298 7570 15334 7604
rect 15368 7570 15404 7604
rect 15438 7570 15474 7604
rect 15508 7570 15544 7604
rect 15578 7570 15614 7604
rect 15648 7570 15684 7604
rect 15718 7570 15754 7604
rect 15788 7570 15824 7604
rect 15858 7570 15894 7604
rect 15928 7570 15964 7604
rect 15998 7570 16032 7604
rect 14698 7544 16032 7570
rect 13152 7535 16032 7544
rect 13152 7508 14774 7535
rect 336 7454 360 7488
rect 394 7454 418 7488
rect 336 7418 418 7454
rect 13152 7474 13194 7508
rect 13228 7474 13264 7508
rect 13298 7474 13334 7508
rect 13368 7474 13404 7508
rect 13438 7474 13474 7508
rect 13508 7474 13544 7508
rect 13578 7474 13614 7508
rect 13648 7474 13684 7508
rect 13718 7474 13754 7508
rect 13788 7474 13824 7508
rect 13858 7474 13894 7508
rect 13928 7474 13964 7508
rect 13998 7474 14034 7508
rect 14068 7474 14104 7508
rect 14138 7474 14174 7508
rect 14208 7474 14244 7508
rect 14278 7474 14314 7508
rect 14348 7474 14384 7508
rect 14418 7474 14454 7508
rect 14488 7474 14524 7508
rect 14558 7474 14594 7508
rect 14628 7474 14664 7508
rect 14698 7501 14774 7508
rect 14808 7501 14844 7535
rect 14878 7501 14914 7535
rect 14948 7501 14984 7535
rect 15018 7501 15054 7535
rect 15088 7501 15124 7535
rect 15158 7501 15194 7535
rect 15228 7501 15264 7535
rect 15298 7501 15334 7535
rect 15368 7501 15404 7535
rect 15438 7501 15474 7535
rect 15508 7501 15544 7535
rect 15578 7501 15614 7535
rect 15648 7501 15684 7535
rect 15718 7501 15754 7535
rect 15788 7501 15824 7535
rect 15858 7501 15894 7535
rect 15928 7501 15964 7535
rect 15998 7501 16032 7535
rect 14698 7474 16032 7501
rect 13152 7466 16032 7474
rect 336 7384 360 7418
rect 394 7384 418 7418
rect 336 7348 418 7384
rect 336 7314 360 7348
rect 394 7314 418 7348
rect 13152 7438 14774 7466
rect 13152 7404 13194 7438
rect 13228 7404 13264 7438
rect 13298 7404 13334 7438
rect 13368 7404 13404 7438
rect 13438 7404 13474 7438
rect 13508 7404 13544 7438
rect 13578 7404 13614 7438
rect 13648 7404 13684 7438
rect 13718 7404 13754 7438
rect 13788 7404 13824 7438
rect 13858 7404 13894 7438
rect 13928 7404 13964 7438
rect 13998 7404 14034 7438
rect 14068 7404 14104 7438
rect 14138 7404 14174 7438
rect 14208 7404 14244 7438
rect 14278 7404 14314 7438
rect 14348 7404 14384 7438
rect 14418 7404 14454 7438
rect 14488 7404 14524 7438
rect 14558 7404 14594 7438
rect 14628 7404 14664 7438
rect 14698 7432 14774 7438
rect 14808 7432 14844 7466
rect 14878 7432 14914 7466
rect 14948 7432 14984 7466
rect 15018 7432 15054 7466
rect 15088 7432 15124 7466
rect 15158 7432 15194 7466
rect 15228 7432 15264 7466
rect 15298 7432 15334 7466
rect 15368 7432 15404 7466
rect 15438 7432 15474 7466
rect 15508 7432 15544 7466
rect 15578 7432 15614 7466
rect 15648 7432 15684 7466
rect 15718 7432 15754 7466
rect 15788 7432 15824 7466
rect 15858 7432 15894 7466
rect 15928 7432 15964 7466
rect 15998 7432 16032 7466
rect 14698 7404 16032 7432
rect 13152 7397 16032 7404
rect 13152 7368 14774 7397
rect 336 7278 418 7314
rect 13152 7334 13194 7368
rect 13228 7334 13264 7368
rect 13298 7334 13334 7368
rect 13368 7334 13404 7368
rect 13438 7334 13474 7368
rect 13508 7334 13544 7368
rect 13578 7334 13614 7368
rect 13648 7334 13684 7368
rect 13718 7334 13754 7368
rect 13788 7334 13824 7368
rect 13858 7334 13894 7368
rect 13928 7334 13964 7368
rect 13998 7334 14034 7368
rect 14068 7334 14104 7368
rect 14138 7334 14174 7368
rect 14208 7334 14244 7368
rect 14278 7334 14314 7368
rect 14348 7334 14384 7368
rect 14418 7334 14454 7368
rect 14488 7334 14524 7368
rect 14558 7334 14594 7368
rect 14628 7334 14664 7368
rect 14698 7363 14774 7368
rect 14808 7363 14844 7397
rect 14878 7363 14914 7397
rect 14948 7363 14984 7397
rect 15018 7363 15054 7397
rect 15088 7363 15124 7397
rect 15158 7363 15194 7397
rect 15228 7363 15264 7397
rect 15298 7363 15334 7397
rect 15368 7363 15404 7397
rect 15438 7363 15474 7397
rect 15508 7363 15544 7397
rect 15578 7363 15614 7397
rect 15648 7363 15684 7397
rect 15718 7363 15754 7397
rect 15788 7363 15824 7397
rect 15858 7363 15894 7397
rect 15928 7363 15964 7397
rect 15998 7363 16032 7397
rect 14698 7334 16032 7363
rect 13152 7328 16032 7334
rect 13152 7298 14774 7328
rect 336 7244 360 7278
rect 394 7244 418 7278
rect 336 7208 418 7244
rect 336 7174 360 7208
rect 394 7174 418 7208
rect 13152 7264 13194 7298
rect 13228 7264 13264 7298
rect 13298 7264 13334 7298
rect 13368 7264 13404 7298
rect 13438 7264 13474 7298
rect 13508 7264 13544 7298
rect 13578 7264 13614 7298
rect 13648 7264 13684 7298
rect 13718 7264 13754 7298
rect 13788 7264 13824 7298
rect 13858 7264 13894 7298
rect 13928 7264 13964 7298
rect 13998 7264 14034 7298
rect 14068 7264 14104 7298
rect 14138 7264 14174 7298
rect 14208 7264 14244 7298
rect 14278 7264 14314 7298
rect 14348 7264 14384 7298
rect 14418 7264 14454 7298
rect 14488 7264 14524 7298
rect 14558 7264 14594 7298
rect 14628 7264 14664 7298
rect 14698 7294 14774 7298
rect 14808 7294 14844 7328
rect 14878 7294 14914 7328
rect 14948 7294 14984 7328
rect 15018 7294 15054 7328
rect 15088 7294 15124 7328
rect 15158 7294 15194 7328
rect 15228 7294 15264 7328
rect 15298 7294 15334 7328
rect 15368 7294 15404 7328
rect 15438 7294 15474 7328
rect 15508 7294 15544 7328
rect 15578 7294 15614 7328
rect 15648 7294 15684 7328
rect 15718 7294 15754 7328
rect 15788 7294 15824 7328
rect 15858 7294 15894 7328
rect 15928 7294 15964 7328
rect 15998 7294 16032 7328
rect 14698 7264 16032 7294
rect 13152 7259 16032 7264
rect 13152 7228 14774 7259
rect 13152 7194 13194 7228
rect 13228 7194 13264 7228
rect 13298 7194 13334 7228
rect 13368 7194 13404 7228
rect 13438 7194 13474 7228
rect 13508 7194 13544 7228
rect 13578 7194 13614 7228
rect 13648 7194 13684 7228
rect 13718 7194 13754 7228
rect 13788 7194 13824 7228
rect 13858 7194 13894 7228
rect 13928 7194 13964 7228
rect 13998 7194 14034 7228
rect 14068 7194 14104 7228
rect 14138 7194 14174 7228
rect 14208 7194 14244 7228
rect 14278 7194 14314 7228
rect 14348 7194 14384 7228
rect 14418 7194 14454 7228
rect 14488 7194 14524 7228
rect 14558 7194 14594 7228
rect 14628 7194 14664 7228
rect 14698 7225 14774 7228
rect 14808 7225 14844 7259
rect 14878 7225 14914 7259
rect 14948 7225 14984 7259
rect 15018 7225 15054 7259
rect 15088 7225 15124 7259
rect 15158 7225 15194 7259
rect 15228 7225 15264 7259
rect 15298 7225 15334 7259
rect 15368 7225 15404 7259
rect 15438 7225 15474 7259
rect 15508 7225 15544 7259
rect 15578 7225 15614 7259
rect 15648 7225 15684 7259
rect 15718 7225 15754 7259
rect 15788 7225 15824 7259
rect 15858 7225 15894 7259
rect 15928 7225 15964 7259
rect 15998 7225 16032 7259
rect 14698 7194 16032 7225
rect 13152 7190 16032 7194
rect 336 7138 418 7174
rect 336 7104 360 7138
rect 394 7104 418 7138
rect 13152 7158 14774 7190
rect 336 7068 418 7104
rect 336 7034 360 7068
rect 394 7034 418 7068
rect 13152 7124 13194 7158
rect 13228 7124 13264 7158
rect 13298 7124 13334 7158
rect 13368 7124 13404 7158
rect 13438 7124 13474 7158
rect 13508 7124 13544 7158
rect 13578 7124 13614 7158
rect 13648 7124 13684 7158
rect 13718 7124 13754 7158
rect 13788 7124 13824 7158
rect 13858 7124 13894 7158
rect 13928 7124 13964 7158
rect 13998 7124 14034 7158
rect 14068 7124 14104 7158
rect 14138 7124 14174 7158
rect 14208 7124 14244 7158
rect 14278 7124 14314 7158
rect 14348 7124 14384 7158
rect 14418 7124 14454 7158
rect 14488 7124 14524 7158
rect 14558 7124 14594 7158
rect 14628 7124 14664 7158
rect 14698 7156 14774 7158
rect 14808 7156 14844 7190
rect 14878 7156 14914 7190
rect 14948 7156 14984 7190
rect 15018 7156 15054 7190
rect 15088 7156 15124 7190
rect 15158 7156 15194 7190
rect 15228 7156 15264 7190
rect 15298 7156 15334 7190
rect 15368 7156 15404 7190
rect 15438 7156 15474 7190
rect 15508 7156 15544 7190
rect 15578 7156 15614 7190
rect 15648 7156 15684 7190
rect 15718 7156 15754 7190
rect 15788 7156 15824 7190
rect 15858 7156 15894 7190
rect 15928 7156 15964 7190
rect 15998 7156 16032 7190
rect 14698 7124 16032 7156
rect 13152 7121 16032 7124
rect 13152 7088 14774 7121
rect 13152 7054 13194 7088
rect 13228 7054 13264 7088
rect 13298 7054 13334 7088
rect 13368 7054 13404 7088
rect 13438 7054 13474 7088
rect 13508 7054 13544 7088
rect 13578 7054 13614 7088
rect 13648 7054 13684 7088
rect 13718 7054 13754 7088
rect 13788 7054 13824 7088
rect 13858 7054 13894 7088
rect 13928 7054 13964 7088
rect 13998 7054 14034 7088
rect 14068 7054 14104 7088
rect 14138 7054 14174 7088
rect 14208 7054 14244 7088
rect 14278 7054 14314 7088
rect 14348 7054 14384 7088
rect 14418 7054 14454 7088
rect 14488 7054 14524 7088
rect 14558 7054 14594 7088
rect 14628 7054 14664 7088
rect 14698 7087 14774 7088
rect 14808 7087 14844 7121
rect 14878 7087 14914 7121
rect 14948 7087 14984 7121
rect 15018 7087 15054 7121
rect 15088 7087 15124 7121
rect 15158 7087 15194 7121
rect 15228 7087 15264 7121
rect 15298 7087 15334 7121
rect 15368 7087 15404 7121
rect 15438 7087 15474 7121
rect 15508 7087 15544 7121
rect 15578 7087 15614 7121
rect 15648 7087 15684 7121
rect 15718 7087 15754 7121
rect 15788 7087 15824 7121
rect 15858 7087 15894 7121
rect 15928 7087 15964 7121
rect 15998 7087 16032 7121
rect 14698 7054 16032 7087
rect 13152 7052 16032 7054
rect 336 6999 418 7034
rect 336 6965 360 6999
rect 394 6965 418 6999
rect 13152 7018 14774 7052
rect 14808 7018 14844 7052
rect 14878 7018 14914 7052
rect 14948 7018 14984 7052
rect 15018 7018 15054 7052
rect 15088 7018 15124 7052
rect 15158 7018 15194 7052
rect 15228 7018 15264 7052
rect 15298 7018 15334 7052
rect 15368 7018 15404 7052
rect 15438 7018 15474 7052
rect 15508 7018 15544 7052
rect 15578 7018 15614 7052
rect 15648 7018 15684 7052
rect 15718 7018 15754 7052
rect 15788 7018 15824 7052
rect 15858 7018 15894 7052
rect 15928 7018 15964 7052
rect 15998 7018 16032 7052
rect 13152 6984 13194 7018
rect 13228 6984 13264 7018
rect 13298 6984 13334 7018
rect 13368 6984 13404 7018
rect 13438 6984 13474 7018
rect 13508 6984 13544 7018
rect 13578 6984 13614 7018
rect 13648 6984 13684 7018
rect 13718 6984 13754 7018
rect 13788 6984 13824 7018
rect 13858 6984 13894 7018
rect 13928 6984 13964 7018
rect 13998 6984 14034 7018
rect 14068 6984 14104 7018
rect 14138 6984 14174 7018
rect 14208 6984 14244 7018
rect 14278 6984 14314 7018
rect 14348 6984 14384 7018
rect 14418 6984 14454 7018
rect 14488 6984 14524 7018
rect 14558 6984 14594 7018
rect 14628 6984 14664 7018
rect 14698 6984 16032 7018
rect 13152 6983 16032 6984
rect 336 6930 418 6965
rect 336 6896 360 6930
rect 394 6896 418 6930
rect 336 6861 418 6896
rect 13152 6949 14774 6983
rect 14808 6949 14844 6983
rect 14878 6949 14914 6983
rect 14948 6949 14984 6983
rect 15018 6949 15054 6983
rect 15088 6949 15124 6983
rect 15158 6949 15194 6983
rect 15228 6949 15264 6983
rect 15298 6949 15334 6983
rect 15368 6949 15404 6983
rect 15438 6949 15474 6983
rect 15508 6949 15544 6983
rect 15578 6949 15614 6983
rect 15648 6949 15684 6983
rect 15718 6949 15754 6983
rect 15788 6949 15824 6983
rect 15858 6949 15894 6983
rect 15928 6949 15964 6983
rect 15998 6949 16032 6983
rect 13152 6948 16032 6949
rect 13152 6914 13194 6948
rect 13228 6914 13264 6948
rect 13298 6914 13334 6948
rect 13368 6914 13404 6948
rect 13438 6914 13474 6948
rect 13508 6914 13544 6948
rect 13578 6914 13614 6948
rect 13648 6914 13684 6948
rect 13718 6914 13754 6948
rect 13788 6914 13824 6948
rect 13858 6914 13894 6948
rect 13928 6914 13964 6948
rect 13998 6914 14034 6948
rect 14068 6914 14104 6948
rect 14138 6914 14174 6948
rect 14208 6914 14244 6948
rect 14278 6914 14314 6948
rect 14348 6914 14384 6948
rect 14418 6914 14454 6948
rect 14488 6914 14524 6948
rect 14558 6914 14594 6948
rect 14628 6914 14664 6948
rect 14698 6914 16032 6948
rect 336 6827 360 6861
rect 394 6827 418 6861
rect 13152 6880 14774 6914
rect 14808 6880 14844 6914
rect 14878 6880 14914 6914
rect 14948 6880 14984 6914
rect 15018 6880 15054 6914
rect 15088 6880 15124 6914
rect 15158 6880 15194 6914
rect 15228 6880 15264 6914
rect 15298 6880 15334 6914
rect 15368 6880 15404 6914
rect 15438 6880 15474 6914
rect 15508 6880 15544 6914
rect 15578 6880 15614 6914
rect 15648 6880 15684 6914
rect 15718 6880 15754 6914
rect 15788 6880 15824 6914
rect 15858 6880 15894 6914
rect 15928 6880 15964 6914
rect 15998 6880 16032 6914
rect 13152 6878 16032 6880
rect 13152 6844 13194 6878
rect 13228 6844 13264 6878
rect 13298 6844 13334 6878
rect 13368 6844 13404 6878
rect 13438 6844 13474 6878
rect 13508 6844 13544 6878
rect 13578 6844 13614 6878
rect 13648 6844 13684 6878
rect 13718 6844 13754 6878
rect 13788 6844 13824 6878
rect 13858 6844 13894 6878
rect 13928 6844 13964 6878
rect 13998 6844 14034 6878
rect 14068 6844 14104 6878
rect 14138 6844 14174 6878
rect 14208 6844 14244 6878
rect 14278 6844 14314 6878
rect 14348 6844 14384 6878
rect 14418 6844 14454 6878
rect 14488 6844 14524 6878
rect 14558 6844 14594 6878
rect 14628 6844 14664 6878
rect 14698 6845 16032 6878
rect 14698 6844 14774 6845
rect 336 6792 418 6827
rect 336 6758 360 6792
rect 394 6758 418 6792
rect 336 6723 418 6758
rect 13152 6811 14774 6844
rect 14808 6811 14844 6845
rect 14878 6811 14914 6845
rect 14948 6811 14984 6845
rect 15018 6811 15054 6845
rect 15088 6811 15124 6845
rect 15158 6811 15194 6845
rect 15228 6811 15264 6845
rect 15298 6811 15334 6845
rect 15368 6811 15404 6845
rect 15438 6811 15474 6845
rect 15508 6811 15544 6845
rect 15578 6811 15614 6845
rect 15648 6811 15684 6845
rect 15718 6811 15754 6845
rect 15788 6811 15824 6845
rect 15858 6811 15894 6845
rect 15928 6811 15964 6845
rect 15998 6811 16032 6845
rect 13152 6808 16032 6811
rect 13152 6774 13194 6808
rect 13228 6774 13264 6808
rect 13298 6774 13334 6808
rect 13368 6774 13404 6808
rect 13438 6774 13474 6808
rect 13508 6774 13544 6808
rect 13578 6774 13614 6808
rect 13648 6774 13684 6808
rect 13718 6774 13754 6808
rect 13788 6774 13824 6808
rect 13858 6774 13894 6808
rect 13928 6774 13964 6808
rect 13998 6774 14034 6808
rect 14068 6774 14104 6808
rect 14138 6774 14174 6808
rect 14208 6774 14244 6808
rect 14278 6774 14314 6808
rect 14348 6774 14384 6808
rect 14418 6774 14454 6808
rect 14488 6774 14524 6808
rect 14558 6774 14594 6808
rect 14628 6774 14664 6808
rect 14698 6776 16032 6808
rect 14698 6774 14774 6776
rect 13152 6742 14774 6774
rect 14808 6742 14844 6776
rect 14878 6742 14914 6776
rect 14948 6742 14984 6776
rect 15018 6742 15054 6776
rect 15088 6742 15124 6776
rect 15158 6742 15194 6776
rect 15228 6742 15264 6776
rect 15298 6742 15334 6776
rect 15368 6742 15404 6776
rect 15438 6742 15474 6776
rect 15508 6742 15544 6776
rect 15578 6742 15614 6776
rect 15648 6742 15684 6776
rect 15718 6742 15754 6776
rect 15788 6742 15824 6776
rect 15858 6742 15894 6776
rect 15928 6742 15964 6776
rect 15998 6742 16032 6776
rect 13152 6738 16032 6742
rect 336 6689 360 6723
rect 394 6689 418 6723
rect 336 6654 418 6689
rect 13152 6704 13194 6738
rect 13228 6704 13264 6738
rect 13298 6704 13334 6738
rect 13368 6704 13404 6738
rect 13438 6704 13474 6738
rect 13508 6704 13544 6738
rect 13578 6704 13614 6738
rect 13648 6704 13684 6738
rect 13718 6704 13754 6738
rect 13788 6704 13824 6738
rect 13858 6704 13894 6738
rect 13928 6704 13964 6738
rect 13998 6704 14034 6738
rect 14068 6704 14104 6738
rect 14138 6704 14174 6738
rect 14208 6704 14244 6738
rect 14278 6704 14314 6738
rect 14348 6704 14384 6738
rect 14418 6704 14454 6738
rect 14488 6704 14524 6738
rect 14558 6704 14594 6738
rect 14628 6704 14664 6738
rect 14698 6707 16032 6738
rect 14698 6704 14774 6707
rect 336 6620 360 6654
rect 394 6620 418 6654
rect 336 6585 418 6620
rect 336 6551 360 6585
rect 394 6551 418 6585
rect 13152 6673 14774 6704
rect 14808 6673 14844 6707
rect 14878 6673 14914 6707
rect 14948 6673 14984 6707
rect 15018 6673 15054 6707
rect 15088 6673 15124 6707
rect 15158 6673 15194 6707
rect 15228 6673 15264 6707
rect 15298 6673 15334 6707
rect 15368 6673 15404 6707
rect 15438 6673 15474 6707
rect 15508 6673 15544 6707
rect 15578 6673 15614 6707
rect 15648 6673 15684 6707
rect 15718 6673 15754 6707
rect 15788 6673 15824 6707
rect 15858 6673 15894 6707
rect 15928 6673 15964 6707
rect 15998 6673 16032 6707
rect 13152 6668 16032 6673
rect 13152 6634 13194 6668
rect 13228 6634 13264 6668
rect 13298 6634 13334 6668
rect 13368 6634 13404 6668
rect 13438 6634 13474 6668
rect 13508 6634 13544 6668
rect 13578 6634 13614 6668
rect 13648 6634 13684 6668
rect 13718 6634 13754 6668
rect 13788 6634 13824 6668
rect 13858 6634 13894 6668
rect 13928 6634 13964 6668
rect 13998 6634 14034 6668
rect 14068 6634 14104 6668
rect 14138 6634 14174 6668
rect 14208 6634 14244 6668
rect 14278 6634 14314 6668
rect 14348 6634 14384 6668
rect 14418 6634 14454 6668
rect 14488 6634 14524 6668
rect 14558 6634 14594 6668
rect 14628 6634 14664 6668
rect 14698 6638 16032 6668
rect 14698 6634 14774 6638
rect 13152 6604 14774 6634
rect 14808 6604 14844 6638
rect 14878 6604 14914 6638
rect 14948 6604 14984 6638
rect 15018 6604 15054 6638
rect 15088 6604 15124 6638
rect 15158 6604 15194 6638
rect 15228 6604 15264 6638
rect 15298 6604 15334 6638
rect 15368 6604 15404 6638
rect 15438 6604 15474 6638
rect 15508 6604 15544 6638
rect 15578 6604 15614 6638
rect 15648 6604 15684 6638
rect 15718 6604 15754 6638
rect 15788 6604 15824 6638
rect 15858 6604 15894 6638
rect 15928 6604 15964 6638
rect 15998 6604 16032 6638
rect 13152 6598 16032 6604
rect 336 6516 418 6551
rect 13152 6564 13194 6598
rect 13228 6564 13264 6598
rect 13298 6564 13334 6598
rect 13368 6564 13404 6598
rect 13438 6564 13474 6598
rect 13508 6564 13544 6598
rect 13578 6564 13614 6598
rect 13648 6564 13684 6598
rect 13718 6564 13754 6598
rect 13788 6564 13824 6598
rect 13858 6564 13894 6598
rect 13928 6564 13964 6598
rect 13998 6564 14034 6598
rect 14068 6564 14104 6598
rect 14138 6564 14174 6598
rect 14208 6564 14244 6598
rect 14278 6564 14314 6598
rect 14348 6564 14384 6598
rect 14418 6564 14454 6598
rect 14488 6564 14524 6598
rect 14558 6564 14594 6598
rect 14628 6564 14664 6598
rect 14698 6569 16032 6598
rect 14698 6564 14774 6569
rect 13152 6535 14774 6564
rect 14808 6535 14844 6569
rect 14878 6535 14914 6569
rect 14948 6535 14984 6569
rect 15018 6535 15054 6569
rect 15088 6535 15124 6569
rect 15158 6535 15194 6569
rect 15228 6535 15264 6569
rect 15298 6535 15334 6569
rect 15368 6535 15404 6569
rect 15438 6535 15474 6569
rect 15508 6535 15544 6569
rect 15578 6535 15614 6569
rect 15648 6535 15684 6569
rect 15718 6535 15754 6569
rect 15788 6535 15824 6569
rect 15858 6535 15894 6569
rect 15928 6535 15964 6569
rect 15998 6535 16032 6569
rect 13152 6528 16032 6535
rect 336 6482 360 6516
rect 394 6482 418 6516
rect 336 6447 418 6482
rect 336 6413 360 6447
rect 394 6413 418 6447
rect 13152 6494 13194 6528
rect 13228 6494 13264 6528
rect 13298 6494 13334 6528
rect 13368 6494 13404 6528
rect 13438 6494 13474 6528
rect 13508 6494 13544 6528
rect 13578 6494 13614 6528
rect 13648 6494 13684 6528
rect 13718 6494 13754 6528
rect 13788 6494 13824 6528
rect 13858 6494 13894 6528
rect 13928 6494 13964 6528
rect 13998 6494 14034 6528
rect 14068 6494 14104 6528
rect 14138 6494 14174 6528
rect 14208 6494 14244 6528
rect 14278 6494 14314 6528
rect 14348 6494 14384 6528
rect 14418 6494 14454 6528
rect 14488 6494 14524 6528
rect 14558 6494 14594 6528
rect 14628 6494 14664 6528
rect 14698 6500 16032 6528
rect 14698 6494 14774 6500
rect 13152 6466 14774 6494
rect 14808 6466 14844 6500
rect 14878 6466 14914 6500
rect 14948 6466 14984 6500
rect 15018 6466 15054 6500
rect 15088 6466 15124 6500
rect 15158 6466 15194 6500
rect 15228 6466 15264 6500
rect 15298 6466 15334 6500
rect 15368 6466 15404 6500
rect 15438 6466 15474 6500
rect 15508 6466 15544 6500
rect 15578 6466 15614 6500
rect 15648 6466 15684 6500
rect 15718 6466 15754 6500
rect 15788 6466 15824 6500
rect 15858 6466 15894 6500
rect 15928 6466 15964 6500
rect 15998 6466 16032 6500
rect 13152 6458 16032 6466
rect 13152 6424 13194 6458
rect 13228 6424 13264 6458
rect 13298 6424 13334 6458
rect 13368 6424 13404 6458
rect 13438 6424 13474 6458
rect 13508 6424 13544 6458
rect 13578 6424 13614 6458
rect 13648 6424 13684 6458
rect 13718 6424 13754 6458
rect 13788 6424 13824 6458
rect 13858 6424 13894 6458
rect 13928 6424 13964 6458
rect 13998 6424 14034 6458
rect 14068 6424 14104 6458
rect 14138 6424 14174 6458
rect 14208 6424 14244 6458
rect 14278 6424 14314 6458
rect 14348 6424 14384 6458
rect 14418 6424 14454 6458
rect 14488 6424 14524 6458
rect 14558 6424 14594 6458
rect 14628 6424 14664 6458
rect 14698 6431 16032 6458
rect 14698 6424 14774 6431
rect 336 6378 418 6413
rect 336 6344 360 6378
rect 394 6344 418 6378
rect 13152 6397 14774 6424
rect 14808 6397 14844 6431
rect 14878 6397 14914 6431
rect 14948 6397 14984 6431
rect 15018 6397 15054 6431
rect 15088 6397 15124 6431
rect 15158 6397 15194 6431
rect 15228 6397 15264 6431
rect 15298 6397 15334 6431
rect 15368 6397 15404 6431
rect 15438 6397 15474 6431
rect 15508 6397 15544 6431
rect 15578 6397 15614 6431
rect 15648 6397 15684 6431
rect 15718 6397 15754 6431
rect 15788 6397 15824 6431
rect 15858 6397 15894 6431
rect 15928 6397 15964 6431
rect 15998 6397 16032 6431
rect 13152 6388 16032 6397
rect 336 6309 418 6344
rect 336 6275 360 6309
rect 394 6275 418 6309
rect 336 6240 418 6275
rect 13152 6354 13194 6388
rect 13228 6354 13264 6388
rect 13298 6354 13334 6388
rect 13368 6354 13404 6388
rect 13438 6354 13474 6388
rect 13508 6354 13544 6388
rect 13578 6354 13614 6388
rect 13648 6354 13684 6388
rect 13718 6354 13754 6388
rect 13788 6354 13824 6388
rect 13858 6354 13894 6388
rect 13928 6354 13964 6388
rect 13998 6354 14034 6388
rect 14068 6354 14104 6388
rect 14138 6354 14174 6388
rect 14208 6354 14244 6388
rect 14278 6354 14314 6388
rect 14348 6354 14384 6388
rect 14418 6354 14454 6388
rect 14488 6354 14524 6388
rect 14558 6354 14594 6388
rect 14628 6354 14664 6388
rect 14698 6362 16032 6388
rect 14698 6354 14774 6362
rect 13152 6328 14774 6354
rect 14808 6328 14844 6362
rect 14878 6328 14914 6362
rect 14948 6328 14984 6362
rect 15018 6328 15054 6362
rect 15088 6328 15124 6362
rect 15158 6328 15194 6362
rect 15228 6328 15264 6362
rect 15298 6328 15334 6362
rect 15368 6328 15404 6362
rect 15438 6328 15474 6362
rect 15508 6328 15544 6362
rect 15578 6328 15614 6362
rect 15648 6328 15684 6362
rect 15718 6328 15754 6362
rect 15788 6328 15824 6362
rect 15858 6328 15894 6362
rect 15928 6328 15964 6362
rect 15998 6328 16032 6362
rect 13152 6318 16032 6328
rect 13152 6284 13194 6318
rect 13228 6284 13264 6318
rect 13298 6284 13334 6318
rect 13368 6284 13404 6318
rect 13438 6284 13474 6318
rect 13508 6284 13544 6318
rect 13578 6284 13614 6318
rect 13648 6284 13684 6318
rect 13718 6284 13754 6318
rect 13788 6284 13824 6318
rect 13858 6284 13894 6318
rect 13928 6284 13964 6318
rect 13998 6284 14034 6318
rect 14068 6284 14104 6318
rect 14138 6284 14174 6318
rect 14208 6284 14244 6318
rect 14278 6284 14314 6318
rect 14348 6284 14384 6318
rect 14418 6284 14454 6318
rect 14488 6284 14524 6318
rect 14558 6284 14594 6318
rect 14628 6284 14664 6318
rect 14698 6293 16032 6318
rect 14698 6284 14774 6293
rect 336 6206 360 6240
rect 394 6206 418 6240
rect 13152 6259 14774 6284
rect 14808 6259 14844 6293
rect 14878 6259 14914 6293
rect 14948 6259 14984 6293
rect 15018 6259 15054 6293
rect 15088 6259 15124 6293
rect 15158 6259 15194 6293
rect 15228 6259 15264 6293
rect 15298 6259 15334 6293
rect 15368 6259 15404 6293
rect 15438 6259 15474 6293
rect 15508 6259 15544 6293
rect 15578 6259 15614 6293
rect 15648 6259 15684 6293
rect 15718 6259 15754 6293
rect 15788 6259 15824 6293
rect 15858 6259 15894 6293
rect 15928 6259 15964 6293
rect 15998 6259 16032 6293
rect 13152 6248 16032 6259
rect 13152 6214 13194 6248
rect 13228 6214 13264 6248
rect 13298 6214 13334 6248
rect 13368 6214 13404 6248
rect 13438 6214 13474 6248
rect 13508 6214 13544 6248
rect 13578 6214 13614 6248
rect 13648 6214 13684 6248
rect 13718 6214 13754 6248
rect 13788 6214 13824 6248
rect 13858 6214 13894 6248
rect 13928 6214 13964 6248
rect 13998 6214 14034 6248
rect 14068 6214 14104 6248
rect 14138 6214 14174 6248
rect 14208 6214 14244 6248
rect 14278 6214 14314 6248
rect 14348 6214 14384 6248
rect 14418 6214 14454 6248
rect 14488 6214 14524 6248
rect 14558 6214 14594 6248
rect 14628 6214 14664 6248
rect 14698 6224 16032 6248
rect 14698 6214 14774 6224
rect 336 6171 418 6206
rect 336 6137 360 6171
rect 394 6137 418 6171
rect 336 6102 418 6137
rect 13152 6190 14774 6214
rect 14808 6190 14844 6224
rect 14878 6190 14914 6224
rect 14948 6190 14984 6224
rect 15018 6190 15054 6224
rect 15088 6190 15124 6224
rect 15158 6190 15194 6224
rect 15228 6190 15264 6224
rect 15298 6190 15334 6224
rect 15368 6190 15404 6224
rect 15438 6190 15474 6224
rect 15508 6190 15544 6224
rect 15578 6190 15614 6224
rect 15648 6190 15684 6224
rect 15718 6190 15754 6224
rect 15788 6190 15824 6224
rect 15858 6190 15894 6224
rect 15928 6190 15964 6224
rect 15998 6190 16032 6224
rect 13152 6178 16032 6190
rect 13152 6144 13194 6178
rect 13228 6144 13264 6178
rect 13298 6144 13334 6178
rect 13368 6144 13404 6178
rect 13438 6144 13474 6178
rect 13508 6144 13544 6178
rect 13578 6144 13614 6178
rect 13648 6144 13684 6178
rect 13718 6144 13754 6178
rect 13788 6144 13824 6178
rect 13858 6144 13894 6178
rect 13928 6144 13964 6178
rect 13998 6144 14034 6178
rect 14068 6144 14104 6178
rect 14138 6144 14174 6178
rect 14208 6144 14244 6178
rect 14278 6144 14314 6178
rect 14348 6144 14384 6178
rect 14418 6144 14454 6178
rect 14488 6144 14524 6178
rect 14558 6144 14594 6178
rect 14628 6144 14664 6178
rect 14698 6155 16032 6178
rect 14698 6144 14774 6155
rect 13152 6121 14774 6144
rect 14808 6121 14844 6155
rect 14878 6121 14914 6155
rect 14948 6121 14984 6155
rect 15018 6121 15054 6155
rect 15088 6121 15124 6155
rect 15158 6121 15194 6155
rect 15228 6121 15264 6155
rect 15298 6121 15334 6155
rect 15368 6121 15404 6155
rect 15438 6121 15474 6155
rect 15508 6121 15544 6155
rect 15578 6121 15614 6155
rect 15648 6121 15684 6155
rect 15718 6121 15754 6155
rect 15788 6121 15824 6155
rect 15858 6121 15894 6155
rect 15928 6121 15964 6155
rect 15998 6121 16032 6155
rect 336 6068 360 6102
rect 394 6068 418 6102
rect 336 6057 418 6068
rect 13152 6108 16032 6121
rect 13152 6074 13194 6108
rect 13228 6074 13264 6108
rect 13298 6074 13334 6108
rect 13368 6074 13404 6108
rect 13438 6074 13474 6108
rect 13508 6074 13544 6108
rect 13578 6074 13614 6108
rect 13648 6074 13684 6108
rect 13718 6074 13754 6108
rect 13788 6074 13824 6108
rect 13858 6074 13894 6108
rect 13928 6074 13964 6108
rect 13998 6074 14034 6108
rect 14068 6074 14104 6108
rect 14138 6074 14174 6108
rect 14208 6074 14244 6108
rect 14278 6074 14314 6108
rect 14348 6074 14384 6108
rect 14418 6074 14454 6108
rect 14488 6074 14524 6108
rect 14558 6074 14594 6108
rect 14628 6074 14664 6108
rect 14698 6086 16032 6108
rect 14698 6074 14774 6086
rect 13152 6057 14774 6074
rect 336 6052 14774 6057
rect 14808 6052 14844 6086
rect 14878 6052 14914 6086
rect 14948 6052 14984 6086
rect 15018 6052 15054 6086
rect 15088 6052 15124 6086
rect 15158 6052 15194 6086
rect 15228 6052 15264 6086
rect 15298 6052 15334 6086
rect 15368 6052 15404 6086
rect 15438 6052 15474 6086
rect 15508 6052 15544 6086
rect 15578 6052 15614 6086
rect 15648 6052 15684 6086
rect 15718 6052 15754 6086
rect 15788 6052 15824 6086
rect 15858 6052 15894 6086
rect 15928 6052 15964 6086
rect 15998 6052 16032 6086
rect 336 6033 16032 6052
rect 336 5999 360 6033
rect 394 5999 429 6033
rect 463 5999 498 6033
rect 532 5999 567 6033
rect 601 5999 636 6033
rect 670 5999 705 6033
rect 739 5999 774 6033
rect 808 5999 843 6033
rect 877 5999 912 6033
rect 946 5999 981 6033
rect 1015 5999 1050 6033
rect 1084 5999 1119 6033
rect 1153 5999 1188 6033
rect 1222 5999 1257 6033
rect 1291 5999 1326 6033
rect 1360 5999 1395 6033
rect 1429 5999 1464 6033
rect 1498 5999 1533 6033
rect 1567 5999 1602 6033
rect 1636 5999 1671 6033
rect 1705 5999 1740 6033
rect 1774 5999 1809 6033
rect 1843 5999 1878 6033
rect 1912 5999 1947 6033
rect 1981 5999 2016 6033
rect 2050 5999 2085 6033
rect 2119 5999 2154 6033
rect 2188 5999 2223 6033
rect 2257 5999 2292 6033
rect 2326 5999 2361 6033
rect 2395 5999 2430 6033
rect 2464 5999 2499 6033
rect 2533 5999 2568 6033
rect 2602 5999 2637 6033
rect 2671 5999 2706 6033
rect 2740 5999 2775 6033
rect 2809 5999 2844 6033
rect 2878 5999 2913 6033
rect 2947 5999 2982 6033
rect 3016 5999 3051 6033
rect 3085 5999 3120 6033
rect 3154 5999 3189 6033
rect 3223 5999 3257 6033
rect 3291 5999 3325 6033
rect 3359 5999 3393 6033
rect 3427 5999 3461 6033
rect 3495 5999 3529 6033
rect 3563 5999 3597 6033
rect 3631 5999 3665 6033
rect 3699 5999 3733 6033
rect 3767 5999 3801 6033
rect 3835 5999 3869 6033
rect 3903 5999 3937 6033
rect 3971 5999 4005 6033
rect 4039 5999 4073 6033
rect 4107 5999 4141 6033
rect 4175 5999 4209 6033
rect 4243 5999 4277 6033
rect 4311 5999 4345 6033
rect 4379 5999 4413 6033
rect 4447 5999 4481 6033
rect 4515 5999 4549 6033
rect 4583 5999 4617 6033
rect 4651 5999 4685 6033
rect 4719 5999 4753 6033
rect 4787 5999 4821 6033
rect 4855 5999 4889 6033
rect 4923 5999 4957 6033
rect 4991 5999 5025 6033
rect 5059 5999 5093 6033
rect 5127 5999 5161 6033
rect 5195 5999 5229 6033
rect 5263 5999 5297 6033
rect 5331 5999 5365 6033
rect 5399 5999 5433 6033
rect 5467 5999 5501 6033
rect 5535 5999 5569 6033
rect 5603 5999 5637 6033
rect 5671 5999 5705 6033
rect 5739 5999 5773 6033
rect 5807 5999 5841 6033
rect 5875 5999 5909 6033
rect 5943 5999 5977 6033
rect 6011 5999 6045 6033
rect 6079 5999 6113 6033
rect 6147 5999 6181 6033
rect 6215 5999 6249 6033
rect 6283 5999 6317 6033
rect 6351 5999 6385 6033
rect 6419 5999 6453 6033
rect 6487 5999 6521 6033
rect 6555 5999 6589 6033
rect 6623 5999 6657 6033
rect 6691 5999 6725 6033
rect 6759 5999 6793 6033
rect 6827 5999 6861 6033
rect 6895 5999 6929 6033
rect 6963 5999 6997 6033
rect 7031 5999 7065 6033
rect 7099 5999 7133 6033
rect 7167 5999 7201 6033
rect 7235 5999 7269 6033
rect 7303 5999 7337 6033
rect 7371 5999 7405 6033
rect 7439 5999 7473 6033
rect 7507 5999 7541 6033
rect 7575 5999 7609 6033
rect 7643 5999 7677 6033
rect 7711 5999 7745 6033
rect 7779 5999 7813 6033
rect 7847 5999 7881 6033
rect 7915 5999 7949 6033
rect 7983 5999 8017 6033
rect 8051 5999 8085 6033
rect 8119 5999 8153 6033
rect 8187 5999 8221 6033
rect 8255 5999 8289 6033
rect 8323 5999 8357 6033
rect 8391 5999 8425 6033
rect 8459 5999 8493 6033
rect 8527 5999 8561 6033
rect 8595 5999 8629 6033
rect 8663 5999 8697 6033
rect 8731 5999 8765 6033
rect 8799 5999 8833 6033
rect 8867 5999 8901 6033
rect 8935 5999 8969 6033
rect 9003 5999 9037 6033
rect 9071 5999 9105 6033
rect 9139 5999 9173 6033
rect 9207 5999 9241 6033
rect 9275 5999 9309 6033
rect 9343 5999 9377 6033
rect 9411 5999 9445 6033
rect 9479 5999 9513 6033
rect 9547 5999 9581 6033
rect 9615 5999 9649 6033
rect 9683 5999 9717 6033
rect 9751 5999 9785 6033
rect 9819 5999 9853 6033
rect 9887 5999 9921 6033
rect 9955 5999 9989 6033
rect 10023 5999 10057 6033
rect 10091 5999 10125 6033
rect 10159 5999 10193 6033
rect 10227 5999 10261 6033
rect 10295 5999 10329 6033
rect 10363 5999 10397 6033
rect 10431 5999 10465 6033
rect 10499 5999 10533 6033
rect 10567 5999 10601 6033
rect 10635 5999 10669 6033
rect 10703 5999 10737 6033
rect 10771 5999 10805 6033
rect 10839 5999 10873 6033
rect 10907 5999 10941 6033
rect 10975 5999 11009 6033
rect 11043 5999 11077 6033
rect 11111 5999 11145 6033
rect 11179 5999 11213 6033
rect 11247 5999 11281 6033
rect 11315 5999 11349 6033
rect 11383 5999 11417 6033
rect 11451 5999 11485 6033
rect 11519 5999 11553 6033
rect 11587 5999 11621 6033
rect 11655 5999 11689 6033
rect 11723 5999 11757 6033
rect 11791 5999 11825 6033
rect 11859 5999 11893 6033
rect 11927 5999 11961 6033
rect 11995 5999 12029 6033
rect 12063 5999 12097 6033
rect 12131 5999 12165 6033
rect 12199 5999 12233 6033
rect 12267 5999 12301 6033
rect 12335 5999 12369 6033
rect 12403 5999 12437 6033
rect 12471 5999 12505 6033
rect 12539 5999 12573 6033
rect 12607 5999 12641 6033
rect 12675 5999 12709 6033
rect 12743 5999 12777 6033
rect 12811 5999 12845 6033
rect 12879 5999 12913 6033
rect 12947 5999 12981 6033
rect 13015 5999 13049 6033
rect 13083 5999 13117 6033
rect 13151 5999 13185 6033
rect 13219 5999 13253 6033
rect 13287 5999 13321 6033
rect 13355 5999 13389 6033
rect 13423 5999 13457 6033
rect 13491 5999 13525 6033
rect 13559 5999 13593 6033
rect 13627 5999 13661 6033
rect 13695 5999 13729 6033
rect 13763 5999 13797 6033
rect 13831 5999 13865 6033
rect 13899 5999 13933 6033
rect 13967 5999 14001 6033
rect 14035 5999 14069 6033
rect 14103 5999 14137 6033
rect 14171 5999 14205 6033
rect 14239 5999 14273 6033
rect 14307 5999 14341 6033
rect 14375 5999 14409 6033
rect 14443 5999 14477 6033
rect 14511 5999 14545 6033
rect 14579 5999 14613 6033
rect 14647 6017 16032 6033
rect 14647 5999 14774 6017
rect 336 5983 14774 5999
rect 14808 5983 14844 6017
rect 14878 5983 14914 6017
rect 14948 5983 14984 6017
rect 15018 5983 15054 6017
rect 15088 5983 15124 6017
rect 15158 5983 15194 6017
rect 15228 5983 15264 6017
rect 15298 5983 15334 6017
rect 15368 5983 15404 6017
rect 15438 5983 15474 6017
rect 15508 5983 15544 6017
rect 15578 5983 15614 6017
rect 15648 5983 15684 6017
rect 15718 5983 15754 6017
rect 15788 5983 15824 6017
rect 15858 5983 15894 6017
rect 15928 5983 15964 6017
rect 15998 5983 16032 6017
rect 336 5975 16032 5983
rect 11482 5951 11564 5975
rect 11482 5917 11506 5951
rect 11540 5917 11564 5951
rect 14740 5948 16032 5975
rect 11482 5882 11564 5917
rect 11482 5848 11506 5882
rect 11540 5848 11564 5882
rect 11482 5813 11564 5848
rect 14740 5914 14774 5948
rect 14808 5914 14844 5948
rect 14878 5914 14914 5948
rect 14948 5914 14984 5948
rect 15018 5914 15054 5948
rect 15088 5914 15124 5948
rect 15158 5914 15194 5948
rect 15228 5914 15264 5948
rect 15298 5914 15334 5948
rect 15368 5914 15404 5948
rect 15438 5914 15474 5948
rect 15508 5914 15544 5948
rect 15578 5914 15614 5948
rect 15648 5914 15684 5948
rect 15718 5914 15754 5948
rect 15788 5914 15824 5948
rect 15858 5914 15894 5948
rect 15928 5914 15964 5948
rect 15998 5914 16032 5948
rect 14740 5879 16032 5914
rect 14740 5845 14774 5879
rect 14808 5845 14844 5879
rect 14878 5845 14914 5879
rect 14948 5845 14984 5879
rect 15018 5845 15054 5879
rect 15088 5845 15124 5879
rect 15158 5845 15194 5879
rect 15228 5845 15264 5879
rect 15298 5845 15334 5879
rect 15368 5845 15404 5879
rect 15438 5845 15474 5879
rect 15508 5845 15544 5879
rect 15578 5845 15614 5879
rect 15648 5845 15684 5879
rect 15718 5845 15754 5879
rect 15788 5845 15824 5879
rect 15858 5845 15894 5879
rect 15928 5845 15964 5879
rect 15998 5845 16032 5879
rect 11482 5779 11506 5813
rect 11540 5779 11564 5813
rect 11482 5744 11564 5779
rect 14740 5810 16032 5845
rect 14740 5776 14774 5810
rect 14808 5776 14844 5810
rect 14878 5776 14914 5810
rect 14948 5776 14984 5810
rect 15018 5776 15054 5810
rect 15088 5776 15124 5810
rect 15158 5776 15194 5810
rect 15228 5776 15264 5810
rect 15298 5776 15334 5810
rect 15368 5776 15404 5810
rect 15438 5776 15474 5810
rect 15508 5776 15544 5810
rect 15578 5776 15614 5810
rect 15648 5776 15684 5810
rect 15718 5776 15754 5810
rect 15788 5776 15824 5810
rect 15858 5776 15894 5810
rect 15928 5776 15964 5810
rect 15998 5776 16032 5810
rect 11482 5710 11506 5744
rect 11540 5710 11564 5744
rect 11482 5675 11564 5710
rect 11482 5641 11506 5675
rect 11540 5641 11564 5675
rect 14740 5741 16032 5776
rect 14740 5707 14774 5741
rect 14808 5707 14844 5741
rect 14878 5707 14914 5741
rect 14948 5707 14984 5741
rect 15018 5707 15054 5741
rect 15088 5707 15124 5741
rect 15158 5707 15194 5741
rect 15228 5707 15264 5741
rect 15298 5707 15334 5741
rect 15368 5707 15404 5741
rect 15438 5707 15474 5741
rect 15508 5707 15544 5741
rect 15578 5707 15614 5741
rect 15648 5707 15684 5741
rect 15718 5707 15754 5741
rect 15788 5707 15824 5741
rect 15858 5707 15894 5741
rect 15928 5707 15964 5741
rect 15998 5707 16032 5741
rect 14740 5672 16032 5707
rect 11482 5606 11564 5641
rect 14740 5638 14774 5672
rect 14808 5638 14844 5672
rect 14878 5638 14914 5672
rect 14948 5638 14984 5672
rect 15018 5638 15054 5672
rect 15088 5638 15124 5672
rect 15158 5638 15194 5672
rect 15228 5638 15264 5672
rect 15298 5638 15334 5672
rect 15368 5638 15404 5672
rect 15438 5638 15474 5672
rect 15508 5638 15544 5672
rect 15578 5638 15614 5672
rect 15648 5638 15684 5672
rect 15718 5638 15754 5672
rect 15788 5638 15824 5672
rect 15858 5638 15894 5672
rect 15928 5638 15964 5672
rect 15998 5638 16032 5672
rect 11482 5572 11506 5606
rect 11540 5572 11564 5606
rect 11482 5537 11564 5572
rect 11482 5503 11506 5537
rect 11540 5503 11564 5537
rect 14740 5603 16032 5638
rect 14740 5569 14774 5603
rect 14808 5569 14844 5603
rect 14878 5569 14914 5603
rect 14948 5569 14984 5603
rect 15018 5569 15054 5603
rect 15088 5569 15124 5603
rect 15158 5569 15194 5603
rect 15228 5569 15264 5603
rect 15298 5569 15334 5603
rect 15368 5569 15404 5603
rect 15438 5569 15474 5603
rect 15508 5569 15544 5603
rect 15578 5569 15614 5603
rect 15648 5569 15684 5603
rect 15718 5569 15754 5603
rect 15788 5569 15824 5603
rect 15858 5569 15894 5603
rect 15928 5569 15964 5603
rect 15998 5569 16032 5603
rect 14740 5534 16032 5569
rect 11482 5468 11564 5503
rect 11482 5434 11506 5468
rect 11540 5434 11564 5468
rect 14740 5500 14774 5534
rect 14808 5500 14844 5534
rect 14878 5500 14914 5534
rect 14948 5500 14984 5534
rect 15018 5500 15054 5534
rect 15088 5500 15124 5534
rect 15158 5500 15194 5534
rect 15228 5500 15264 5534
rect 15298 5500 15334 5534
rect 15368 5500 15404 5534
rect 15438 5500 15474 5534
rect 15508 5500 15544 5534
rect 15578 5500 15614 5534
rect 15648 5500 15684 5534
rect 15718 5500 15754 5534
rect 15788 5500 15824 5534
rect 15858 5500 15894 5534
rect 15928 5500 15964 5534
rect 15998 5500 16032 5534
rect 14740 5465 16032 5500
rect 11482 5399 11564 5434
rect 11482 5365 11506 5399
rect 11540 5365 11564 5399
rect 11482 5330 11564 5365
rect 14740 5431 14774 5465
rect 14808 5431 14844 5465
rect 14878 5431 14914 5465
rect 14948 5431 14984 5465
rect 15018 5431 15054 5465
rect 15088 5431 15124 5465
rect 15158 5431 15194 5465
rect 15228 5431 15264 5465
rect 15298 5431 15334 5465
rect 15368 5431 15404 5465
rect 15438 5431 15474 5465
rect 15508 5431 15544 5465
rect 15578 5431 15614 5465
rect 15648 5431 15684 5465
rect 15718 5431 15754 5465
rect 15788 5431 15824 5465
rect 15858 5431 15894 5465
rect 15928 5431 15964 5465
rect 15998 5431 16032 5465
rect 14740 5396 16032 5431
rect 14740 5362 14774 5396
rect 14808 5362 14844 5396
rect 14878 5362 14914 5396
rect 14948 5362 14984 5396
rect 15018 5362 15054 5396
rect 15088 5362 15124 5396
rect 15158 5362 15194 5396
rect 15228 5362 15264 5396
rect 15298 5362 15334 5396
rect 15368 5362 15404 5396
rect 15438 5362 15474 5396
rect 15508 5362 15544 5396
rect 15578 5362 15614 5396
rect 15648 5362 15684 5396
rect 15718 5362 15754 5396
rect 15788 5362 15824 5396
rect 15858 5362 15894 5396
rect 15928 5362 15964 5396
rect 15998 5362 16032 5396
rect 11482 5296 11506 5330
rect 11540 5296 11564 5330
rect 14740 5327 16032 5362
rect 11482 5261 11564 5296
rect 11482 5227 11506 5261
rect 11540 5227 11564 5261
rect 11482 5192 11564 5227
rect 14740 5293 14774 5327
rect 14808 5293 14844 5327
rect 14878 5293 14914 5327
rect 14948 5293 14984 5327
rect 15018 5293 15054 5327
rect 15088 5293 15124 5327
rect 15158 5293 15194 5327
rect 15228 5293 15264 5327
rect 15298 5293 15334 5327
rect 15368 5293 15404 5327
rect 15438 5293 15474 5327
rect 15508 5293 15544 5327
rect 15578 5293 15614 5327
rect 15648 5293 15684 5327
rect 15718 5293 15754 5327
rect 15788 5293 15824 5327
rect 15858 5293 15894 5327
rect 15928 5293 15964 5327
rect 15998 5293 16032 5327
rect 14740 5258 16032 5293
rect 14740 5224 14774 5258
rect 14808 5224 14844 5258
rect 14878 5224 14914 5258
rect 14948 5224 14984 5258
rect 15018 5224 15054 5258
rect 15088 5224 15124 5258
rect 15158 5224 15194 5258
rect 15228 5224 15264 5258
rect 15298 5224 15334 5258
rect 15368 5224 15404 5258
rect 15438 5224 15474 5258
rect 15508 5224 15544 5258
rect 15578 5224 15614 5258
rect 15648 5224 15684 5258
rect 15718 5224 15754 5258
rect 15788 5224 15824 5258
rect 15858 5224 15894 5258
rect 15928 5224 15964 5258
rect 15998 5224 16032 5258
rect 11482 5158 11506 5192
rect 11540 5158 11564 5192
rect 11482 5123 11564 5158
rect 14740 5190 16032 5224
rect 14740 5156 14774 5190
rect 14808 5156 14844 5190
rect 14878 5156 14914 5190
rect 14948 5156 14984 5190
rect 15018 5156 15054 5190
rect 15088 5156 15124 5190
rect 15158 5156 15194 5190
rect 15228 5156 15264 5190
rect 15298 5156 15334 5190
rect 15368 5156 15404 5190
rect 15438 5156 15474 5190
rect 15508 5156 15544 5190
rect 15578 5156 15614 5190
rect 15648 5156 15684 5190
rect 15718 5156 15754 5190
rect 15788 5156 15824 5190
rect 15858 5156 15894 5190
rect 15928 5156 15964 5190
rect 15998 5156 16032 5190
rect 11482 5089 11506 5123
rect 11540 5089 11564 5123
rect 11482 5054 11564 5089
rect 11482 5020 11506 5054
rect 11540 5020 11564 5054
rect 14740 5122 16032 5156
rect 14740 5088 14774 5122
rect 14808 5088 14844 5122
rect 14878 5088 14914 5122
rect 14948 5088 14984 5122
rect 15018 5088 15054 5122
rect 15088 5088 15124 5122
rect 15158 5088 15194 5122
rect 15228 5088 15264 5122
rect 15298 5088 15334 5122
rect 15368 5088 15404 5122
rect 15438 5088 15474 5122
rect 15508 5088 15544 5122
rect 15578 5088 15614 5122
rect 15648 5088 15684 5122
rect 15718 5088 15754 5122
rect 15788 5088 15824 5122
rect 15858 5088 15894 5122
rect 15928 5088 15964 5122
rect 15998 5088 16032 5122
rect 14740 5054 16032 5088
rect 11482 4985 11564 5020
rect 14740 5020 14774 5054
rect 14808 5020 14844 5054
rect 14878 5020 14914 5054
rect 14948 5020 14984 5054
rect 15018 5020 15054 5054
rect 15088 5020 15124 5054
rect 15158 5020 15194 5054
rect 15228 5020 15264 5054
rect 15298 5020 15334 5054
rect 15368 5020 15404 5054
rect 15438 5020 15474 5054
rect 15508 5020 15544 5054
rect 15578 5020 15614 5054
rect 15648 5020 15684 5054
rect 15718 5020 15754 5054
rect 15788 5020 15824 5054
rect 15858 5020 15894 5054
rect 15928 5020 15964 5054
rect 15998 5020 16032 5054
rect 11482 4951 11506 4985
rect 11540 4951 11564 4985
rect 11482 4916 11564 4951
rect 11482 4882 11506 4916
rect 11540 4882 11564 4916
rect 14740 4986 16032 5020
rect 14740 4952 14774 4986
rect 14808 4952 14844 4986
rect 14878 4952 14914 4986
rect 14948 4952 14984 4986
rect 15018 4952 15054 4986
rect 15088 4952 15124 4986
rect 15158 4952 15194 4986
rect 15228 4952 15264 4986
rect 15298 4952 15334 4986
rect 15368 4952 15404 4986
rect 15438 4952 15474 4986
rect 15508 4952 15544 4986
rect 15578 4952 15614 4986
rect 15648 4952 15684 4986
rect 15718 4952 15754 4986
rect 15788 4952 15824 4986
rect 15858 4952 15894 4986
rect 15928 4952 15964 4986
rect 15998 4952 16032 4986
rect 14740 4918 16032 4952
rect 11482 4847 11564 4882
rect 11482 4813 11506 4847
rect 11540 4813 11564 4847
rect 14740 4884 14774 4918
rect 14808 4884 14844 4918
rect 14878 4884 14914 4918
rect 14948 4884 14984 4918
rect 15018 4884 15054 4918
rect 15088 4884 15124 4918
rect 15158 4884 15194 4918
rect 15228 4884 15264 4918
rect 15298 4884 15334 4918
rect 15368 4884 15404 4918
rect 15438 4884 15474 4918
rect 15508 4884 15544 4918
rect 15578 4884 15614 4918
rect 15648 4884 15684 4918
rect 15718 4884 15754 4918
rect 15788 4884 15824 4918
rect 15858 4884 15894 4918
rect 15928 4884 15964 4918
rect 15998 4884 16032 4918
rect 14740 4850 16032 4884
rect 11482 4778 11564 4813
rect 11482 4744 11506 4778
rect 11540 4744 11564 4778
rect 11482 4709 11564 4744
rect 14740 4816 14774 4850
rect 14808 4816 14844 4850
rect 14878 4816 14914 4850
rect 14948 4816 14984 4850
rect 15018 4816 15054 4850
rect 15088 4816 15124 4850
rect 15158 4816 15194 4850
rect 15228 4816 15264 4850
rect 15298 4816 15334 4850
rect 15368 4816 15404 4850
rect 15438 4816 15474 4850
rect 15508 4816 15544 4850
rect 15578 4816 15614 4850
rect 15648 4816 15684 4850
rect 15718 4816 15754 4850
rect 15788 4816 15824 4850
rect 15858 4816 15894 4850
rect 15928 4816 15964 4850
rect 15998 4816 16032 4850
rect 14740 4782 16032 4816
rect 14740 4748 14774 4782
rect 14808 4748 14844 4782
rect 14878 4748 14914 4782
rect 14948 4748 14984 4782
rect 15018 4748 15054 4782
rect 15088 4748 15124 4782
rect 15158 4748 15194 4782
rect 15228 4748 15264 4782
rect 15298 4748 15334 4782
rect 15368 4748 15404 4782
rect 15438 4748 15474 4782
rect 15508 4748 15544 4782
rect 15578 4748 15614 4782
rect 15648 4748 15684 4782
rect 15718 4748 15754 4782
rect 15788 4748 15824 4782
rect 15858 4748 15894 4782
rect 15928 4748 15964 4782
rect 15998 4748 16032 4782
rect 11482 4675 11506 4709
rect 11540 4675 11564 4709
rect 14740 4714 16032 4748
rect 11482 4640 11564 4675
rect 11482 4606 11506 4640
rect 11540 4606 11564 4640
rect 11482 4571 11564 4606
rect 14740 4680 14774 4714
rect 14808 4680 14844 4714
rect 14878 4680 14914 4714
rect 14948 4680 14984 4714
rect 15018 4680 15054 4714
rect 15088 4680 15124 4714
rect 15158 4680 15194 4714
rect 15228 4680 15264 4714
rect 15298 4680 15334 4714
rect 15368 4680 15404 4714
rect 15438 4680 15474 4714
rect 15508 4680 15544 4714
rect 15578 4680 15614 4714
rect 15648 4680 15684 4714
rect 15718 4680 15754 4714
rect 15788 4680 15824 4714
rect 15858 4680 15894 4714
rect 15928 4680 15964 4714
rect 15998 4680 16032 4714
rect 14740 4646 16032 4680
rect 14740 4612 14774 4646
rect 14808 4612 14844 4646
rect 14878 4612 14914 4646
rect 14948 4612 14984 4646
rect 15018 4612 15054 4646
rect 15088 4612 15124 4646
rect 15158 4612 15194 4646
rect 15228 4612 15264 4646
rect 15298 4612 15334 4646
rect 15368 4612 15404 4646
rect 15438 4612 15474 4646
rect 15508 4612 15544 4646
rect 15578 4612 15614 4646
rect 15648 4612 15684 4646
rect 15718 4612 15754 4646
rect 15788 4612 15824 4646
rect 15858 4612 15894 4646
rect 15928 4612 15964 4646
rect 15998 4612 16032 4646
rect 11482 4537 11506 4571
rect 11540 4537 11564 4571
rect 11482 4502 11564 4537
rect 14740 4578 16032 4612
rect 14740 4544 14774 4578
rect 14808 4544 14844 4578
rect 14878 4544 14914 4578
rect 14948 4544 14984 4578
rect 15018 4544 15054 4578
rect 15088 4544 15124 4578
rect 15158 4544 15194 4578
rect 15228 4544 15264 4578
rect 15298 4544 15334 4578
rect 15368 4544 15404 4578
rect 15438 4544 15474 4578
rect 15508 4544 15544 4578
rect 15578 4544 15614 4578
rect 15648 4544 15684 4578
rect 15718 4544 15754 4578
rect 15788 4544 15824 4578
rect 15858 4544 15894 4578
rect 15928 4544 15964 4578
rect 15998 4544 16032 4578
rect 11482 4468 11506 4502
rect 11540 4468 11564 4502
rect 11482 4433 11564 4468
rect 14740 4510 16032 4544
rect 14740 4476 14774 4510
rect 14808 4476 14844 4510
rect 14878 4476 14914 4510
rect 14948 4476 14984 4510
rect 15018 4476 15054 4510
rect 15088 4476 15124 4510
rect 15158 4476 15194 4510
rect 15228 4476 15264 4510
rect 15298 4476 15334 4510
rect 15368 4476 15404 4510
rect 15438 4476 15474 4510
rect 15508 4476 15544 4510
rect 15578 4476 15614 4510
rect 15648 4476 15684 4510
rect 15718 4476 15754 4510
rect 15788 4476 15824 4510
rect 15858 4476 15894 4510
rect 15928 4476 15964 4510
rect 15998 4476 16032 4510
rect 14740 4442 16032 4476
rect 11482 4399 11506 4433
rect 11540 4399 11564 4433
rect 11482 4364 11564 4399
rect 14740 4408 14774 4442
rect 14808 4408 14844 4442
rect 14878 4408 14914 4442
rect 14948 4408 14984 4442
rect 15018 4408 15054 4442
rect 15088 4408 15124 4442
rect 15158 4408 15194 4442
rect 15228 4408 15264 4442
rect 15298 4408 15334 4442
rect 15368 4408 15404 4442
rect 15438 4408 15474 4442
rect 15508 4408 15544 4442
rect 15578 4408 15614 4442
rect 15648 4408 15684 4442
rect 15718 4408 15754 4442
rect 15788 4408 15824 4442
rect 15858 4408 15894 4442
rect 15928 4408 15964 4442
rect 15998 4408 16032 4442
rect 11482 4330 11506 4364
rect 11540 4330 11564 4364
rect 11482 4295 11564 4330
rect 11482 4261 11506 4295
rect 11540 4261 11564 4295
rect 14740 4374 16032 4408
rect 14740 4340 14774 4374
rect 14808 4340 14844 4374
rect 14878 4340 14914 4374
rect 14948 4340 14984 4374
rect 15018 4340 15054 4374
rect 15088 4340 15124 4374
rect 15158 4340 15194 4374
rect 15228 4340 15264 4374
rect 15298 4340 15334 4374
rect 15368 4340 15404 4374
rect 15438 4340 15474 4374
rect 15508 4340 15544 4374
rect 15578 4340 15614 4374
rect 15648 4340 15684 4374
rect 15718 4340 15754 4374
rect 15788 4340 15824 4374
rect 15858 4340 15894 4374
rect 15928 4340 15964 4374
rect 15998 4340 16032 4374
rect 14740 4306 16032 4340
rect 11482 4226 11564 4261
rect 14740 4272 14774 4306
rect 14808 4272 14844 4306
rect 14878 4272 14914 4306
rect 14948 4272 14984 4306
rect 15018 4272 15054 4306
rect 15088 4272 15124 4306
rect 15158 4272 15194 4306
rect 15228 4272 15264 4306
rect 15298 4272 15334 4306
rect 15368 4272 15404 4306
rect 15438 4272 15474 4306
rect 15508 4272 15544 4306
rect 15578 4272 15614 4306
rect 15648 4272 15684 4306
rect 15718 4272 15754 4306
rect 15788 4272 15824 4306
rect 15858 4272 15894 4306
rect 15928 4272 15964 4306
rect 15998 4272 16032 4306
rect 14740 4238 16032 4272
rect 11482 4192 11506 4226
rect 11540 4192 11564 4226
rect 11482 4157 11564 4192
rect 11482 4123 11506 4157
rect 11540 4123 11564 4157
rect 14740 4204 14774 4238
rect 14808 4204 14844 4238
rect 14878 4204 14914 4238
rect 14948 4204 14984 4238
rect 15018 4204 15054 4238
rect 15088 4204 15124 4238
rect 15158 4204 15194 4238
rect 15228 4204 15264 4238
rect 15298 4204 15334 4238
rect 15368 4204 15404 4238
rect 15438 4204 15474 4238
rect 15508 4204 15544 4238
rect 15578 4204 15614 4238
rect 15648 4204 15684 4238
rect 15718 4204 15754 4238
rect 15788 4204 15824 4238
rect 15858 4204 15894 4238
rect 15928 4204 15964 4238
rect 15998 4204 16032 4238
rect 14740 4170 16032 4204
rect 14740 4136 14774 4170
rect 14808 4136 14844 4170
rect 14878 4136 14914 4170
rect 14948 4136 14984 4170
rect 15018 4136 15054 4170
rect 15088 4136 15124 4170
rect 15158 4136 15194 4170
rect 15228 4136 15264 4170
rect 15298 4136 15334 4170
rect 15368 4136 15404 4170
rect 15438 4136 15474 4170
rect 15508 4136 15544 4170
rect 15578 4136 15614 4170
rect 15648 4136 15684 4170
rect 15718 4136 15754 4170
rect 15788 4136 15824 4170
rect 15858 4136 15894 4170
rect 15928 4136 15964 4170
rect 15998 4136 16032 4170
rect 11482 4088 11564 4123
rect 11482 4054 11506 4088
rect 11540 4054 11564 4088
rect 11482 4051 11564 4054
rect 14740 4102 16032 4136
rect 14740 4068 14774 4102
rect 14808 4068 14844 4102
rect 14878 4068 14914 4102
rect 14948 4068 14984 4102
rect 15018 4068 15054 4102
rect 15088 4068 15124 4102
rect 15158 4068 15194 4102
rect 15228 4068 15264 4102
rect 15298 4068 15334 4102
rect 15368 4068 15404 4102
rect 15438 4068 15474 4102
rect 15508 4068 15544 4102
rect 15578 4068 15614 4102
rect 15648 4068 15684 4102
rect 15718 4068 15754 4102
rect 15788 4068 15824 4102
rect 15858 4068 15894 4102
rect 15928 4068 15964 4102
rect 15998 4068 16032 4102
rect 14740 4051 16032 4068
rect 11482 4019 11588 4051
rect 11482 3985 11506 4019
rect 11540 4017 11588 4019
rect 11622 4017 11657 4051
rect 11691 4017 11726 4051
rect 11760 4017 11795 4051
rect 11829 4017 11864 4051
rect 11898 4017 11933 4051
rect 11967 4017 12002 4051
rect 12036 4017 12071 4051
rect 12105 4017 12140 4051
rect 12174 4017 12209 4051
rect 12243 4017 12278 4051
rect 12312 4017 12347 4051
rect 12381 4017 12416 4051
rect 12450 4017 12485 4051
rect 12519 4017 12554 4051
rect 12588 4017 12623 4051
rect 12657 4017 12692 4051
rect 12726 4017 12761 4051
rect 12795 4017 12830 4051
rect 12864 4017 12899 4051
rect 12933 4017 12968 4051
rect 13002 4017 13037 4051
rect 13071 4017 13106 4051
rect 13140 4017 13175 4051
rect 13209 4017 13244 4051
rect 13278 4017 13313 4051
rect 13347 4017 13382 4051
rect 13416 4017 13451 4051
rect 13485 4017 13520 4051
rect 13554 4017 13589 4051
rect 13623 4017 13658 4051
rect 13692 4017 13727 4051
rect 13761 4017 13796 4051
rect 13830 4017 13865 4051
rect 13899 4017 13934 4051
rect 13968 4017 14002 4051
rect 14036 4017 14070 4051
rect 14104 4017 14138 4051
rect 14172 4017 14206 4051
rect 14240 4017 14274 4051
rect 14308 4017 14342 4051
rect 14376 4017 14410 4051
rect 14444 4017 14478 4051
rect 14512 4017 14546 4051
rect 14580 4017 14614 4051
rect 14648 4017 14682 4051
rect 14716 4034 16032 4051
rect 14716 4017 14774 4034
rect 11540 3985 11564 4017
rect 11482 3950 11564 3985
rect 11482 3916 11506 3950
rect 11540 3916 11564 3950
rect 14740 4000 14774 4017
rect 14808 4000 14844 4034
rect 14878 4000 14914 4034
rect 14948 4000 14984 4034
rect 15018 4000 15054 4034
rect 15088 4000 15124 4034
rect 15158 4000 15194 4034
rect 15228 4000 15264 4034
rect 15298 4000 15334 4034
rect 15368 4000 15404 4034
rect 15438 4000 15474 4034
rect 15508 4000 15544 4034
rect 15578 4000 15614 4034
rect 15648 4000 15684 4034
rect 15718 4000 15754 4034
rect 15788 4000 15824 4034
rect 15858 4000 15894 4034
rect 15928 4000 15964 4034
rect 15998 4000 16032 4034
rect 14740 3966 16032 4000
rect 11482 3881 11564 3916
rect 11482 3847 11506 3881
rect 11540 3847 11564 3881
rect 11482 3812 11564 3847
rect 14740 3932 14774 3966
rect 14808 3932 14844 3966
rect 14878 3932 14914 3966
rect 14948 3932 14984 3966
rect 15018 3932 15054 3966
rect 15088 3932 15124 3966
rect 15158 3932 15194 3966
rect 15228 3932 15264 3966
rect 15298 3932 15334 3966
rect 15368 3932 15404 3966
rect 15438 3932 15474 3966
rect 15508 3932 15544 3966
rect 15578 3932 15614 3966
rect 15648 3932 15684 3966
rect 15718 3932 15754 3966
rect 15788 3932 15824 3966
rect 15858 3932 15894 3966
rect 15928 3932 15964 3966
rect 15998 3932 16032 3966
rect 14740 3898 16032 3932
rect 14740 3864 14774 3898
rect 14808 3864 14844 3898
rect 14878 3864 14914 3898
rect 14948 3864 14984 3898
rect 15018 3864 15054 3898
rect 15088 3864 15124 3898
rect 15158 3864 15194 3898
rect 15228 3864 15264 3898
rect 15298 3864 15334 3898
rect 15368 3864 15404 3898
rect 15438 3864 15474 3898
rect 15508 3864 15544 3898
rect 15578 3864 15614 3898
rect 15648 3864 15684 3898
rect 15718 3864 15754 3898
rect 15788 3864 15824 3898
rect 15858 3864 15894 3898
rect 15928 3864 15964 3898
rect 15998 3864 16032 3898
rect 11482 3778 11506 3812
rect 11540 3778 11564 3812
rect 14740 3830 16032 3864
rect 14740 3796 14774 3830
rect 14808 3796 14844 3830
rect 14878 3796 14914 3830
rect 14948 3796 14984 3830
rect 15018 3796 15054 3830
rect 15088 3796 15124 3830
rect 15158 3796 15194 3830
rect 15228 3796 15264 3830
rect 15298 3796 15334 3830
rect 15368 3796 15404 3830
rect 15438 3796 15474 3830
rect 15508 3796 15544 3830
rect 15578 3796 15614 3830
rect 15648 3796 15684 3830
rect 15718 3796 15754 3830
rect 15788 3796 15824 3830
rect 15858 3796 15894 3830
rect 15928 3796 15964 3830
rect 15998 3796 16032 3830
rect 11482 3743 11564 3778
rect 11482 3709 11506 3743
rect 11540 3709 11564 3743
rect 11482 3674 11564 3709
rect 14740 3762 16032 3796
rect 14740 3728 14774 3762
rect 14808 3728 14844 3762
rect 14878 3728 14914 3762
rect 14948 3728 14984 3762
rect 15018 3728 15054 3762
rect 15088 3728 15124 3762
rect 15158 3728 15194 3762
rect 15228 3728 15264 3762
rect 15298 3728 15334 3762
rect 15368 3728 15404 3762
rect 15438 3728 15474 3762
rect 15508 3728 15544 3762
rect 15578 3728 15614 3762
rect 15648 3728 15684 3762
rect 15718 3728 15754 3762
rect 15788 3728 15824 3762
rect 15858 3728 15894 3762
rect 15928 3728 15964 3762
rect 15998 3728 16032 3762
rect 14740 3694 16032 3728
rect 11482 3640 11506 3674
rect 11540 3640 11564 3674
rect 11482 3605 11564 3640
rect 14740 3660 14774 3694
rect 14808 3660 14844 3694
rect 14878 3660 14914 3694
rect 14948 3660 14984 3694
rect 15018 3660 15054 3694
rect 15088 3660 15124 3694
rect 15158 3660 15194 3694
rect 15228 3660 15264 3694
rect 15298 3660 15334 3694
rect 15368 3660 15404 3694
rect 15438 3660 15474 3694
rect 15508 3660 15544 3694
rect 15578 3660 15614 3694
rect 15648 3660 15684 3694
rect 15718 3660 15754 3694
rect 15788 3660 15824 3694
rect 15858 3660 15894 3694
rect 15928 3660 15964 3694
rect 15998 3660 16032 3694
rect 11482 3571 11506 3605
rect 11540 3571 11564 3605
rect 11482 3536 11564 3571
rect 11482 3502 11506 3536
rect 11540 3502 11564 3536
rect 14740 3626 16032 3660
rect 14740 3592 14774 3626
rect 14808 3592 14844 3626
rect 14878 3592 14914 3626
rect 14948 3592 14984 3626
rect 15018 3592 15054 3626
rect 15088 3592 15124 3626
rect 15158 3592 15194 3626
rect 15228 3592 15264 3626
rect 15298 3592 15334 3626
rect 15368 3592 15404 3626
rect 15438 3592 15474 3626
rect 15508 3592 15544 3626
rect 15578 3592 15614 3626
rect 15648 3592 15684 3626
rect 15718 3592 15754 3626
rect 15788 3592 15824 3626
rect 15858 3592 15894 3626
rect 15928 3592 15964 3626
rect 15998 3592 16032 3626
rect 14740 3558 16032 3592
rect 11482 3467 11564 3502
rect 14740 3524 14774 3558
rect 14808 3524 14844 3558
rect 14878 3524 14914 3558
rect 14948 3524 14984 3558
rect 15018 3524 15054 3558
rect 15088 3524 15124 3558
rect 15158 3524 15194 3558
rect 15228 3524 15264 3558
rect 15298 3524 15334 3558
rect 15368 3524 15404 3558
rect 15438 3524 15474 3558
rect 15508 3524 15544 3558
rect 15578 3524 15614 3558
rect 15648 3524 15684 3558
rect 15718 3524 15754 3558
rect 15788 3524 15824 3558
rect 15858 3524 15894 3558
rect 15928 3524 15964 3558
rect 15998 3524 16032 3558
rect 14740 3490 16032 3524
rect 11482 3433 11506 3467
rect 11540 3433 11564 3467
rect 11482 3398 11564 3433
rect 11482 3364 11506 3398
rect 11540 3364 11564 3398
rect 14740 3456 14774 3490
rect 14808 3456 14844 3490
rect 14878 3456 14914 3490
rect 14948 3456 14984 3490
rect 15018 3456 15054 3490
rect 15088 3456 15124 3490
rect 15158 3456 15194 3490
rect 15228 3456 15264 3490
rect 15298 3456 15334 3490
rect 15368 3456 15404 3490
rect 15438 3456 15474 3490
rect 15508 3456 15544 3490
rect 15578 3456 15614 3490
rect 15648 3456 15684 3490
rect 15718 3456 15754 3490
rect 15788 3456 15824 3490
rect 15858 3456 15894 3490
rect 15928 3456 15964 3490
rect 15998 3456 16032 3490
rect 14740 3422 16032 3456
rect 14740 3388 14774 3422
rect 14808 3388 14844 3422
rect 14878 3388 14914 3422
rect 14948 3388 14984 3422
rect 15018 3388 15054 3422
rect 15088 3388 15124 3422
rect 15158 3388 15194 3422
rect 15228 3388 15264 3422
rect 15298 3388 15334 3422
rect 15368 3388 15404 3422
rect 15438 3388 15474 3422
rect 15508 3388 15544 3422
rect 15578 3388 15614 3422
rect 15648 3388 15684 3422
rect 15718 3388 15754 3422
rect 15788 3388 15824 3422
rect 15858 3388 15894 3422
rect 15928 3388 15964 3422
rect 15998 3388 16032 3422
rect 11482 3329 11564 3364
rect 11482 3295 11506 3329
rect 11540 3295 11564 3329
rect 14740 3354 16032 3388
rect 11482 3260 11564 3295
rect 11482 3226 11506 3260
rect 11540 3226 11564 3260
rect 11482 3191 11564 3226
rect 14740 3320 14774 3354
rect 14808 3320 14844 3354
rect 14878 3320 14914 3354
rect 14948 3320 14984 3354
rect 15018 3320 15054 3354
rect 15088 3320 15124 3354
rect 15158 3320 15194 3354
rect 15228 3320 15264 3354
rect 15298 3320 15334 3354
rect 15368 3320 15404 3354
rect 15438 3320 15474 3354
rect 15508 3320 15544 3354
rect 15578 3320 15614 3354
rect 15648 3320 15684 3354
rect 15718 3320 15754 3354
rect 15788 3320 15824 3354
rect 15858 3320 15894 3354
rect 15928 3320 15964 3354
rect 15998 3320 16032 3354
rect 14740 3286 16032 3320
rect 14740 3252 14774 3286
rect 14808 3252 14844 3286
rect 14878 3252 14914 3286
rect 14948 3252 14984 3286
rect 15018 3252 15054 3286
rect 15088 3252 15124 3286
rect 15158 3252 15194 3286
rect 15228 3252 15264 3286
rect 15298 3252 15334 3286
rect 15368 3252 15404 3286
rect 15438 3252 15474 3286
rect 15508 3252 15544 3286
rect 15578 3252 15614 3286
rect 15648 3252 15684 3286
rect 15718 3252 15754 3286
rect 15788 3252 15824 3286
rect 15858 3252 15894 3286
rect 15928 3252 15964 3286
rect 15998 3252 16032 3286
rect 11482 3157 11506 3191
rect 11540 3157 11564 3191
rect 14740 3218 16032 3252
rect 14740 3184 14774 3218
rect 14808 3184 14844 3218
rect 14878 3184 14914 3218
rect 14948 3184 14984 3218
rect 15018 3184 15054 3218
rect 15088 3184 15124 3218
rect 15158 3184 15194 3218
rect 15228 3184 15264 3218
rect 15298 3184 15334 3218
rect 15368 3184 15404 3218
rect 15438 3184 15474 3218
rect 15508 3184 15544 3218
rect 15578 3184 15614 3218
rect 15648 3184 15684 3218
rect 15718 3184 15754 3218
rect 15788 3184 15824 3218
rect 15858 3184 15894 3218
rect 15928 3184 15964 3218
rect 15998 3184 16032 3218
rect 11482 3122 11564 3157
rect 11482 3088 11506 3122
rect 11540 3088 11564 3122
rect 11482 3053 11564 3088
rect 14740 3150 16032 3184
rect 14740 3116 14774 3150
rect 14808 3116 14844 3150
rect 14878 3116 14914 3150
rect 14948 3116 14984 3150
rect 15018 3116 15054 3150
rect 15088 3116 15124 3150
rect 15158 3116 15194 3150
rect 15228 3116 15264 3150
rect 15298 3116 15334 3150
rect 15368 3116 15404 3150
rect 15438 3116 15474 3150
rect 15508 3116 15544 3150
rect 15578 3116 15614 3150
rect 15648 3116 15684 3150
rect 15718 3116 15754 3150
rect 15788 3116 15824 3150
rect 15858 3116 15894 3150
rect 15928 3116 15964 3150
rect 15998 3116 16032 3150
rect 14740 3082 16032 3116
rect 11482 3019 11506 3053
rect 11540 3019 11564 3053
rect 11482 2984 11564 3019
rect 14740 3048 14774 3082
rect 14808 3048 14844 3082
rect 14878 3048 14914 3082
rect 14948 3048 14984 3082
rect 15018 3048 15054 3082
rect 15088 3048 15124 3082
rect 15158 3048 15194 3082
rect 15228 3048 15264 3082
rect 15298 3048 15334 3082
rect 15368 3048 15404 3082
rect 15438 3048 15474 3082
rect 15508 3048 15544 3082
rect 15578 3048 15614 3082
rect 15648 3048 15684 3082
rect 15718 3048 15754 3082
rect 15788 3048 15824 3082
rect 15858 3048 15894 3082
rect 15928 3048 15964 3082
rect 15998 3048 16032 3082
rect 11482 2950 11506 2984
rect 11540 2950 11564 2984
rect 11482 2915 11564 2950
rect 14740 3014 16032 3048
rect 14740 2980 14774 3014
rect 14808 2980 14844 3014
rect 14878 2980 14914 3014
rect 14948 2980 14984 3014
rect 15018 2980 15054 3014
rect 15088 2980 15124 3014
rect 15158 2980 15194 3014
rect 15228 2980 15264 3014
rect 15298 2980 15334 3014
rect 15368 2980 15404 3014
rect 15438 2980 15474 3014
rect 15508 2980 15544 3014
rect 15578 2980 15614 3014
rect 15648 2980 15684 3014
rect 15718 2980 15754 3014
rect 15788 2980 15824 3014
rect 15858 2980 15894 3014
rect 15928 2980 15964 3014
rect 15998 2980 16032 3014
rect 14740 2946 16032 2980
rect 11482 2881 11506 2915
rect 11540 2881 11564 2915
rect 11482 2846 11564 2881
rect 14740 2912 14774 2946
rect 14808 2912 14844 2946
rect 14878 2912 14914 2946
rect 14948 2912 14984 2946
rect 15018 2912 15054 2946
rect 15088 2912 15124 2946
rect 15158 2912 15194 2946
rect 15228 2912 15264 2946
rect 15298 2912 15334 2946
rect 15368 2912 15404 2946
rect 15438 2912 15474 2946
rect 15508 2912 15544 2946
rect 15578 2912 15614 2946
rect 15648 2912 15684 2946
rect 15718 2912 15754 2946
rect 15788 2912 15824 2946
rect 15858 2912 15894 2946
rect 15928 2912 15964 2946
rect 15998 2912 16032 2946
rect 14740 2878 16032 2912
rect 11482 2812 11506 2846
rect 11540 2812 11564 2846
rect 11482 2777 11564 2812
rect 11482 2743 11506 2777
rect 11540 2743 11564 2777
rect 14740 2844 14774 2878
rect 14808 2844 14844 2878
rect 14878 2844 14914 2878
rect 14948 2844 14984 2878
rect 15018 2844 15054 2878
rect 15088 2844 15124 2878
rect 15158 2844 15194 2878
rect 15228 2844 15264 2878
rect 15298 2844 15334 2878
rect 15368 2844 15404 2878
rect 15438 2844 15474 2878
rect 15508 2844 15544 2878
rect 15578 2844 15614 2878
rect 15648 2844 15684 2878
rect 15718 2844 15754 2878
rect 15788 2844 15824 2878
rect 15858 2844 15894 2878
rect 15928 2844 15964 2878
rect 15998 2844 16032 2878
rect 14740 2810 16032 2844
rect 14740 2776 14774 2810
rect 14808 2776 14844 2810
rect 14878 2776 14914 2810
rect 14948 2776 14984 2810
rect 15018 2776 15054 2810
rect 15088 2776 15124 2810
rect 15158 2776 15194 2810
rect 15228 2776 15264 2810
rect 15298 2776 15334 2810
rect 15368 2776 15404 2810
rect 15438 2776 15474 2810
rect 15508 2776 15544 2810
rect 15578 2776 15614 2810
rect 15648 2776 15684 2810
rect 15718 2776 15754 2810
rect 15788 2776 15824 2810
rect 15858 2776 15894 2810
rect 15928 2776 15964 2810
rect 15998 2776 16032 2810
rect 11482 2708 11564 2743
rect 14740 2742 16032 2776
rect 11482 2674 11506 2708
rect 11540 2674 11564 2708
rect 11482 2639 11564 2674
rect 11482 2605 11506 2639
rect 11540 2605 11564 2639
rect 14740 2708 14774 2742
rect 14808 2708 14844 2742
rect 14878 2708 14914 2742
rect 14948 2708 14984 2742
rect 15018 2708 15054 2742
rect 15088 2708 15124 2742
rect 15158 2708 15194 2742
rect 15228 2708 15264 2742
rect 15298 2708 15334 2742
rect 15368 2708 15404 2742
rect 15438 2708 15474 2742
rect 15508 2708 15544 2742
rect 15578 2708 15614 2742
rect 15648 2708 15684 2742
rect 15718 2708 15754 2742
rect 15788 2708 15824 2742
rect 15858 2708 15894 2742
rect 15928 2708 15964 2742
rect 15998 2708 16032 2742
rect 14740 2674 16032 2708
rect 14740 2640 14774 2674
rect 14808 2640 14844 2674
rect 14878 2640 14914 2674
rect 14948 2640 14984 2674
rect 15018 2640 15054 2674
rect 15088 2640 15124 2674
rect 15158 2640 15194 2674
rect 15228 2640 15264 2674
rect 15298 2640 15334 2674
rect 15368 2640 15404 2674
rect 15438 2640 15474 2674
rect 15508 2640 15544 2674
rect 15578 2640 15614 2674
rect 15648 2640 15684 2674
rect 15718 2640 15754 2674
rect 15788 2640 15824 2674
rect 15858 2640 15894 2674
rect 15928 2640 15964 2674
rect 15998 2640 16032 2674
rect 11482 2570 11564 2605
rect 11482 2536 11506 2570
rect 11540 2536 11564 2570
rect 14740 2606 16032 2640
rect 14740 2572 14774 2606
rect 14808 2572 14844 2606
rect 14878 2572 14914 2606
rect 14948 2572 14984 2606
rect 15018 2572 15054 2606
rect 15088 2572 15124 2606
rect 15158 2572 15194 2606
rect 15228 2572 15264 2606
rect 15298 2572 15334 2606
rect 15368 2572 15404 2606
rect 15438 2572 15474 2606
rect 15508 2572 15544 2606
rect 15578 2572 15614 2606
rect 15648 2572 15684 2606
rect 15718 2572 15754 2606
rect 15788 2572 15824 2606
rect 15858 2572 15894 2606
rect 15928 2572 15964 2606
rect 15998 2572 16032 2606
rect 11482 2501 11564 2536
rect 11482 2467 11506 2501
rect 11540 2467 11564 2501
rect 11482 2431 11564 2467
rect 14740 2538 16032 2572
rect 14740 2504 14774 2538
rect 14808 2504 14844 2538
rect 14878 2504 14914 2538
rect 14948 2504 14984 2538
rect 15018 2504 15054 2538
rect 15088 2504 15124 2538
rect 15158 2504 15194 2538
rect 15228 2504 15264 2538
rect 15298 2504 15334 2538
rect 15368 2504 15404 2538
rect 15438 2504 15474 2538
rect 15508 2504 15544 2538
rect 15578 2504 15614 2538
rect 15648 2504 15684 2538
rect 15718 2504 15754 2538
rect 15788 2504 15824 2538
rect 15858 2504 15894 2538
rect 15928 2504 15964 2538
rect 15998 2504 16032 2538
rect 14740 2470 16032 2504
rect 11482 2397 11506 2431
rect 11540 2397 11564 2431
rect 14740 2436 14774 2470
rect 14808 2436 14844 2470
rect 14878 2436 14914 2470
rect 14948 2436 14984 2470
rect 15018 2436 15054 2470
rect 15088 2436 15124 2470
rect 15158 2436 15194 2470
rect 15228 2436 15264 2470
rect 15298 2436 15334 2470
rect 15368 2436 15404 2470
rect 15438 2436 15474 2470
rect 15508 2436 15544 2470
rect 15578 2436 15614 2470
rect 15648 2436 15684 2470
rect 15718 2436 15754 2470
rect 15788 2436 15824 2470
rect 15858 2436 15894 2470
rect 15928 2436 15964 2470
rect 15998 2436 16032 2470
rect 14740 2402 16032 2436
rect 11482 2361 11564 2397
rect 11482 2327 11506 2361
rect 11540 2327 11564 2361
rect 11482 2291 11564 2327
rect 14740 2368 14774 2402
rect 14808 2368 14844 2402
rect 14878 2368 14914 2402
rect 14948 2368 14984 2402
rect 15018 2368 15054 2402
rect 15088 2368 15124 2402
rect 15158 2368 15194 2402
rect 15228 2368 15264 2402
rect 15298 2368 15334 2402
rect 15368 2368 15404 2402
rect 15438 2368 15474 2402
rect 15508 2368 15544 2402
rect 15578 2368 15614 2402
rect 15648 2368 15684 2402
rect 15718 2368 15754 2402
rect 15788 2368 15824 2402
rect 15858 2368 15894 2402
rect 15928 2368 15964 2402
rect 15998 2368 16032 2402
rect 14740 2334 16032 2368
rect 11482 2257 11506 2291
rect 11540 2257 11564 2291
rect 11482 2221 11564 2257
rect 14740 2300 14774 2334
rect 14808 2300 14844 2334
rect 14878 2300 14914 2334
rect 14948 2300 14984 2334
rect 15018 2300 15054 2334
rect 15088 2300 15124 2334
rect 15158 2300 15194 2334
rect 15228 2300 15264 2334
rect 15298 2300 15334 2334
rect 15368 2300 15404 2334
rect 15438 2300 15474 2334
rect 15508 2300 15544 2334
rect 15578 2300 15614 2334
rect 15648 2300 15684 2334
rect 15718 2300 15754 2334
rect 15788 2300 15824 2334
rect 15858 2300 15894 2334
rect 15928 2300 15964 2334
rect 15998 2300 16032 2334
rect 14740 2266 16032 2300
rect 11482 2187 11506 2221
rect 11540 2187 11564 2221
rect 11482 2151 11564 2187
rect 11482 2117 11506 2151
rect 11540 2117 11564 2151
rect 14740 2232 14774 2266
rect 14808 2232 14844 2266
rect 14878 2232 14914 2266
rect 14948 2232 14984 2266
rect 15018 2232 15054 2266
rect 15088 2232 15124 2266
rect 15158 2232 15194 2266
rect 15228 2232 15264 2266
rect 15298 2232 15334 2266
rect 15368 2232 15404 2266
rect 15438 2232 15474 2266
rect 15508 2232 15544 2266
rect 15578 2232 15614 2266
rect 15648 2232 15684 2266
rect 15718 2232 15754 2266
rect 15788 2232 15824 2266
rect 15858 2232 15894 2266
rect 15928 2232 15964 2266
rect 15998 2232 16032 2266
rect 14740 2198 16032 2232
rect 14740 2164 14774 2198
rect 14808 2164 14844 2198
rect 14878 2164 14914 2198
rect 14948 2164 14984 2198
rect 15018 2164 15054 2198
rect 15088 2164 15124 2198
rect 15158 2164 15194 2198
rect 15228 2164 15264 2198
rect 15298 2164 15334 2198
rect 15368 2164 15404 2198
rect 15438 2164 15474 2198
rect 15508 2164 15544 2198
rect 15578 2164 15614 2198
rect 15648 2164 15684 2198
rect 15718 2164 15754 2198
rect 15788 2164 15824 2198
rect 15858 2164 15894 2198
rect 15928 2164 15964 2198
rect 15998 2164 16032 2198
rect 11482 2093 11564 2117
rect 14740 2130 16032 2164
rect 14740 2096 14774 2130
rect 14808 2096 14844 2130
rect 14878 2096 14914 2130
rect 14948 2096 14984 2130
rect 15018 2096 15054 2130
rect 15088 2096 15124 2130
rect 15158 2096 15194 2130
rect 15228 2096 15264 2130
rect 15298 2096 15334 2130
rect 15368 2096 15404 2130
rect 15438 2096 15474 2130
rect 15508 2096 15544 2130
rect 15578 2096 15614 2130
rect 15648 2096 15684 2130
rect 15718 2096 15754 2130
rect 15788 2096 15824 2130
rect 15858 2096 15894 2130
rect 15928 2096 15964 2130
rect 15998 2096 16032 2130
rect 14740 2093 16032 2096
rect 336 2069 16032 2093
rect 370 2035 405 2069
rect 439 2035 474 2069
rect 508 2035 543 2069
rect 577 2035 612 2069
rect 646 2035 681 2069
rect 715 2035 750 2069
rect 784 2035 819 2069
rect 853 2035 888 2069
rect 922 2035 957 2069
rect 991 2035 1026 2069
rect 1060 2035 1095 2069
rect 1129 2035 1164 2069
rect 1198 2035 1233 2069
rect 1267 2035 1302 2069
rect 1336 2035 1371 2069
rect 1405 2035 1440 2069
rect 1474 2035 1509 2069
rect 1543 2035 1578 2069
rect 1612 2035 1647 2069
rect 1681 2035 1716 2069
rect 1750 2035 1785 2069
rect 1819 2035 1854 2069
rect 1888 2035 1923 2069
rect 1957 2035 1992 2069
rect 2026 2035 2061 2069
rect 2095 2035 2130 2069
rect 2164 2035 2199 2069
rect 2233 2035 2268 2069
rect 2302 2035 2337 2069
rect 2371 2035 2406 2069
rect 2440 2035 2475 2069
rect 2509 2035 2544 2069
rect 2578 2035 2613 2069
rect 2647 2035 2682 2069
rect 2716 2035 2751 2069
rect 2785 2035 2820 2069
rect 2854 2035 2889 2069
rect 2923 2035 2958 2069
rect 2992 2035 3027 2069
rect 3061 2035 3096 2069
rect 3130 2035 3165 2069
rect 3199 2035 3234 2069
rect 3268 2035 3303 2069
rect 3337 2035 3372 2069
rect 3406 2035 3441 2069
rect 3475 2035 3510 2069
rect 3544 2035 3579 2069
rect 3613 2035 3648 2069
rect 3682 2035 3717 2069
rect 3751 2035 3786 2069
rect 3820 2035 3855 2069
rect 3889 2035 3924 2069
rect 3958 2035 3993 2069
rect 4027 2035 4062 2069
rect 4096 2035 4131 2069
rect 4165 2035 4200 2069
rect 4234 2035 4269 2069
rect 4303 2035 4338 2069
rect 4372 2035 4407 2069
rect 4441 2035 4475 2069
rect 4509 2035 4543 2069
rect 4577 2035 4611 2069
rect 4645 2035 4679 2069
rect 4713 2035 4747 2069
rect 4781 2035 4815 2069
rect 4849 2035 4883 2069
rect 4917 2035 4951 2069
rect 4985 2035 5019 2069
rect 5053 2035 5087 2069
rect 5121 2035 5155 2069
rect 5189 2035 5223 2069
rect 5257 2035 5291 2069
rect 5325 2035 5359 2069
rect 5393 2035 5427 2069
rect 5461 2035 5495 2069
rect 5529 2035 5563 2069
rect 5597 2035 5631 2069
rect 5665 2035 5699 2069
rect 5733 2035 5767 2069
rect 5801 2035 5835 2069
rect 5869 2035 5903 2069
rect 5937 2035 5971 2069
rect 6005 2035 6039 2069
rect 6073 2035 6107 2069
rect 6141 2035 6175 2069
rect 6209 2035 6243 2069
rect 6277 2035 6311 2069
rect 6345 2035 6379 2069
rect 6413 2035 6447 2069
rect 6481 2035 6515 2069
rect 6549 2035 6583 2069
rect 6617 2035 6651 2069
rect 6685 2035 6719 2069
rect 6753 2035 6787 2069
rect 6821 2035 6855 2069
rect 6889 2035 6923 2069
rect 6957 2035 6991 2069
rect 7025 2035 7059 2069
rect 7093 2035 7127 2069
rect 7161 2035 7195 2069
rect 7229 2035 7263 2069
rect 7297 2035 7331 2069
rect 7365 2035 7399 2069
rect 7433 2035 7467 2069
rect 7501 2035 7535 2069
rect 7569 2035 7603 2069
rect 7637 2035 7671 2069
rect 7705 2035 7739 2069
rect 7773 2035 7807 2069
rect 7841 2035 7875 2069
rect 7909 2035 7943 2069
rect 7977 2035 8011 2069
rect 8045 2035 8079 2069
rect 8113 2035 8147 2069
rect 8181 2035 8215 2069
rect 8249 2035 8283 2069
rect 8317 2035 8351 2069
rect 8385 2035 8419 2069
rect 8453 2035 8487 2069
rect 8521 2035 8555 2069
rect 8589 2035 8623 2069
rect 8657 2035 8691 2069
rect 8725 2035 8759 2069
rect 8793 2035 8827 2069
rect 8861 2035 8895 2069
rect 8929 2035 8963 2069
rect 8997 2035 9031 2069
rect 9065 2035 9099 2069
rect 9133 2035 9167 2069
rect 9201 2035 9235 2069
rect 9269 2035 9303 2069
rect 9337 2035 9371 2069
rect 9405 2035 9439 2069
rect 9473 2035 9507 2069
rect 9541 2035 9575 2069
rect 9609 2035 9643 2069
rect 9677 2035 9711 2069
rect 9745 2035 9779 2069
rect 9813 2035 9847 2069
rect 9881 2035 9915 2069
rect 9949 2035 9983 2069
rect 10017 2035 10051 2069
rect 10085 2035 10119 2069
rect 10153 2035 10187 2069
rect 10221 2035 10255 2069
rect 10289 2035 10323 2069
rect 10357 2035 10391 2069
rect 10425 2035 10459 2069
rect 10493 2035 10527 2069
rect 10561 2035 10595 2069
rect 10629 2035 10663 2069
rect 10697 2035 10731 2069
rect 10765 2035 10799 2069
rect 10833 2035 10867 2069
rect 10901 2035 10935 2069
rect 10969 2035 11003 2069
rect 11037 2035 11071 2069
rect 11105 2035 11139 2069
rect 11173 2035 11207 2069
rect 11241 2035 11275 2069
rect 11309 2035 11343 2069
rect 11377 2035 11411 2069
rect 11445 2035 11479 2069
rect 11513 2035 11547 2069
rect 11581 2035 11615 2069
rect 11649 2035 11683 2069
rect 11717 2035 11751 2069
rect 11785 2035 11819 2069
rect 11853 2035 11887 2069
rect 11921 2035 11955 2069
rect 11989 2035 12023 2069
rect 12057 2035 12091 2069
rect 12125 2035 12159 2069
rect 12193 2035 12227 2069
rect 12261 2035 12295 2069
rect 12329 2035 12363 2069
rect 12397 2035 12431 2069
rect 12465 2035 12499 2069
rect 12533 2035 12567 2069
rect 12601 2035 12635 2069
rect 12669 2035 12703 2069
rect 12737 2035 12771 2069
rect 12805 2035 12839 2069
rect 12873 2035 12907 2069
rect 12941 2035 12975 2069
rect 13009 2035 13043 2069
rect 13077 2035 13111 2069
rect 13145 2035 13179 2069
rect 13213 2035 13247 2069
rect 13281 2035 13315 2069
rect 13349 2035 13383 2069
rect 13417 2035 13451 2069
rect 13485 2035 13519 2069
rect 13553 2035 13587 2069
rect 13621 2035 13655 2069
rect 13689 2035 13723 2069
rect 13757 2035 13791 2069
rect 13825 2035 13859 2069
rect 13893 2035 13927 2069
rect 13961 2035 13995 2069
rect 14029 2035 14063 2069
rect 14097 2035 14131 2069
rect 14165 2035 14199 2069
rect 14233 2035 14267 2069
rect 14301 2035 14335 2069
rect 14369 2035 14403 2069
rect 14437 2035 14471 2069
rect 14505 2035 14539 2069
rect 14573 2035 14607 2069
rect 14641 2035 14675 2069
rect 14709 2062 16032 2069
rect 14709 2035 14774 2062
rect 336 2028 14774 2035
rect 14808 2028 14844 2062
rect 14878 2028 14914 2062
rect 14948 2028 14984 2062
rect 15018 2028 15054 2062
rect 15088 2028 15124 2062
rect 15158 2028 15194 2062
rect 15228 2028 15264 2062
rect 15298 2028 15334 2062
rect 15368 2028 15404 2062
rect 15438 2028 15474 2062
rect 15508 2028 15544 2062
rect 15578 2028 15614 2062
rect 15648 2028 15684 2062
rect 15718 2028 15754 2062
rect 15788 2028 15824 2062
rect 15858 2028 15894 2062
rect 15928 2028 15964 2062
rect 15998 2028 16032 2062
rect 336 2011 16032 2028
rect 336 1959 418 2011
rect 336 1925 360 1959
rect 394 1925 418 1959
rect 13152 2001 16032 2011
rect 13152 1967 13194 2001
rect 13228 1967 13264 2001
rect 13298 1967 13334 2001
rect 13368 1967 13404 2001
rect 13438 1967 13474 2001
rect 13508 1967 13544 2001
rect 13578 1967 13614 2001
rect 13648 1967 13684 2001
rect 13718 1967 13754 2001
rect 13788 1967 13824 2001
rect 13858 1967 13894 2001
rect 13928 1967 13964 2001
rect 13998 1967 14034 2001
rect 14068 1967 14104 2001
rect 14138 1967 14174 2001
rect 14208 1967 14244 2001
rect 14278 1967 14314 2001
rect 14348 1967 14384 2001
rect 14418 1967 14454 2001
rect 14488 1967 14524 2001
rect 14558 1967 14594 2001
rect 14628 1967 14664 2001
rect 14698 1994 16032 2001
rect 14698 1967 14774 1994
rect 13152 1960 14774 1967
rect 14808 1960 14844 1994
rect 14878 1960 14914 1994
rect 14948 1960 14984 1994
rect 15018 1960 15054 1994
rect 15088 1960 15124 1994
rect 15158 1960 15194 1994
rect 15228 1960 15264 1994
rect 15298 1960 15334 1994
rect 15368 1960 15404 1994
rect 15438 1960 15474 1994
rect 15508 1960 15544 1994
rect 15578 1960 15614 1994
rect 15648 1960 15684 1994
rect 15718 1960 15754 1994
rect 15788 1960 15824 1994
rect 15858 1960 15894 1994
rect 15928 1960 15964 1994
rect 15998 1960 16032 1994
rect 336 1889 418 1925
rect 336 1855 360 1889
rect 394 1855 418 1889
rect 13152 1931 16032 1960
rect 13152 1897 13194 1931
rect 13228 1897 13264 1931
rect 13298 1897 13334 1931
rect 13368 1897 13404 1931
rect 13438 1897 13474 1931
rect 13508 1897 13544 1931
rect 13578 1897 13614 1931
rect 13648 1897 13684 1931
rect 13718 1897 13754 1931
rect 13788 1897 13824 1931
rect 13858 1897 13894 1931
rect 13928 1897 13964 1931
rect 13998 1897 14034 1931
rect 14068 1897 14104 1931
rect 14138 1897 14174 1931
rect 14208 1897 14244 1931
rect 14278 1897 14314 1931
rect 14348 1897 14384 1931
rect 14418 1897 14454 1931
rect 14488 1897 14524 1931
rect 14558 1897 14594 1931
rect 14628 1897 14664 1931
rect 14698 1926 16032 1931
rect 14698 1897 14774 1926
rect 13152 1892 14774 1897
rect 14808 1892 14844 1926
rect 14878 1892 14914 1926
rect 14948 1892 14984 1926
rect 15018 1892 15054 1926
rect 15088 1892 15124 1926
rect 15158 1892 15194 1926
rect 15228 1892 15264 1926
rect 15298 1892 15334 1926
rect 15368 1892 15404 1926
rect 15438 1892 15474 1926
rect 15508 1892 15544 1926
rect 15578 1892 15614 1926
rect 15648 1892 15684 1926
rect 15718 1892 15754 1926
rect 15788 1892 15824 1926
rect 15858 1892 15894 1926
rect 15928 1892 15964 1926
rect 15998 1892 16032 1926
rect 13152 1861 16032 1892
rect 336 1819 418 1855
rect 336 1785 360 1819
rect 394 1785 418 1819
rect 13152 1827 13194 1861
rect 13228 1827 13264 1861
rect 13298 1827 13334 1861
rect 13368 1827 13404 1861
rect 13438 1827 13474 1861
rect 13508 1827 13544 1861
rect 13578 1827 13614 1861
rect 13648 1827 13684 1861
rect 13718 1827 13754 1861
rect 13788 1827 13824 1861
rect 13858 1827 13894 1861
rect 13928 1827 13964 1861
rect 13998 1827 14034 1861
rect 14068 1827 14104 1861
rect 14138 1827 14174 1861
rect 14208 1827 14244 1861
rect 14278 1827 14314 1861
rect 14348 1827 14384 1861
rect 14418 1827 14454 1861
rect 14488 1827 14524 1861
rect 14558 1827 14594 1861
rect 14628 1827 14664 1861
rect 14698 1858 16032 1861
rect 14698 1827 14774 1858
rect 13152 1824 14774 1827
rect 14808 1824 14844 1858
rect 14878 1824 14914 1858
rect 14948 1824 14984 1858
rect 15018 1824 15054 1858
rect 15088 1824 15124 1858
rect 15158 1824 15194 1858
rect 15228 1824 15264 1858
rect 15298 1824 15334 1858
rect 15368 1824 15404 1858
rect 15438 1824 15474 1858
rect 15508 1824 15544 1858
rect 15578 1824 15614 1858
rect 15648 1824 15684 1858
rect 15718 1824 15754 1858
rect 15788 1824 15824 1858
rect 15858 1824 15894 1858
rect 15928 1824 15964 1858
rect 15998 1824 16032 1858
rect 336 1749 418 1785
rect 336 1715 360 1749
rect 394 1715 418 1749
rect 336 1679 418 1715
rect 13152 1791 16032 1824
rect 13152 1757 13194 1791
rect 13228 1757 13264 1791
rect 13298 1757 13334 1791
rect 13368 1757 13404 1791
rect 13438 1757 13474 1791
rect 13508 1757 13544 1791
rect 13578 1757 13614 1791
rect 13648 1757 13684 1791
rect 13718 1757 13754 1791
rect 13788 1757 13824 1791
rect 13858 1757 13894 1791
rect 13928 1757 13964 1791
rect 13998 1757 14034 1791
rect 14068 1757 14104 1791
rect 14138 1757 14174 1791
rect 14208 1757 14244 1791
rect 14278 1757 14314 1791
rect 14348 1757 14384 1791
rect 14418 1757 14454 1791
rect 14488 1757 14524 1791
rect 14558 1757 14594 1791
rect 14628 1757 14664 1791
rect 14698 1790 16032 1791
rect 14698 1757 14774 1790
rect 13152 1756 14774 1757
rect 14808 1756 14844 1790
rect 14878 1756 14914 1790
rect 14948 1756 14984 1790
rect 15018 1756 15054 1790
rect 15088 1756 15124 1790
rect 15158 1756 15194 1790
rect 15228 1756 15264 1790
rect 15298 1756 15334 1790
rect 15368 1756 15404 1790
rect 15438 1756 15474 1790
rect 15508 1756 15544 1790
rect 15578 1756 15614 1790
rect 15648 1756 15684 1790
rect 15718 1756 15754 1790
rect 15788 1756 15824 1790
rect 15858 1756 15894 1790
rect 15928 1756 15964 1790
rect 15998 1756 16032 1790
rect 13152 1722 16032 1756
rect 13152 1721 14774 1722
rect 336 1645 360 1679
rect 394 1645 418 1679
rect 13152 1687 13194 1721
rect 13228 1687 13264 1721
rect 13298 1687 13334 1721
rect 13368 1687 13404 1721
rect 13438 1687 13474 1721
rect 13508 1687 13544 1721
rect 13578 1687 13614 1721
rect 13648 1687 13684 1721
rect 13718 1687 13754 1721
rect 13788 1687 13824 1721
rect 13858 1687 13894 1721
rect 13928 1687 13964 1721
rect 13998 1687 14034 1721
rect 14068 1687 14104 1721
rect 14138 1687 14174 1721
rect 14208 1687 14244 1721
rect 14278 1687 14314 1721
rect 14348 1687 14384 1721
rect 14418 1687 14454 1721
rect 14488 1687 14524 1721
rect 14558 1687 14594 1721
rect 14628 1687 14664 1721
rect 14698 1688 14774 1721
rect 14808 1688 14844 1722
rect 14878 1688 14914 1722
rect 14948 1688 14984 1722
rect 15018 1688 15054 1722
rect 15088 1688 15124 1722
rect 15158 1688 15194 1722
rect 15228 1688 15264 1722
rect 15298 1688 15334 1722
rect 15368 1688 15404 1722
rect 15438 1688 15474 1722
rect 15508 1688 15544 1722
rect 15578 1688 15614 1722
rect 15648 1688 15684 1722
rect 15718 1688 15754 1722
rect 15788 1688 15824 1722
rect 15858 1688 15894 1722
rect 15928 1688 15964 1722
rect 15998 1688 16032 1722
rect 14698 1687 16032 1688
rect 13152 1654 16032 1687
rect 13152 1651 14774 1654
rect 336 1609 418 1645
rect 336 1575 360 1609
rect 394 1575 418 1609
rect 336 1539 418 1575
rect 13152 1617 13194 1651
rect 13228 1617 13264 1651
rect 13298 1617 13334 1651
rect 13368 1617 13404 1651
rect 13438 1617 13474 1651
rect 13508 1617 13544 1651
rect 13578 1617 13614 1651
rect 13648 1617 13684 1651
rect 13718 1617 13754 1651
rect 13788 1617 13824 1651
rect 13858 1617 13894 1651
rect 13928 1617 13964 1651
rect 13998 1617 14034 1651
rect 14068 1617 14104 1651
rect 14138 1617 14174 1651
rect 14208 1617 14244 1651
rect 14278 1617 14314 1651
rect 14348 1617 14384 1651
rect 14418 1617 14454 1651
rect 14488 1617 14524 1651
rect 14558 1617 14594 1651
rect 14628 1617 14664 1651
rect 14698 1620 14774 1651
rect 14808 1620 14844 1654
rect 14878 1620 14914 1654
rect 14948 1620 14984 1654
rect 15018 1620 15054 1654
rect 15088 1620 15124 1654
rect 15158 1620 15194 1654
rect 15228 1620 15264 1654
rect 15298 1620 15334 1654
rect 15368 1620 15404 1654
rect 15438 1620 15474 1654
rect 15508 1620 15544 1654
rect 15578 1620 15614 1654
rect 15648 1620 15684 1654
rect 15718 1620 15754 1654
rect 15788 1620 15824 1654
rect 15858 1620 15894 1654
rect 15928 1620 15964 1654
rect 15998 1620 16032 1654
rect 14698 1617 16032 1620
rect 13152 1586 16032 1617
rect 13152 1581 14774 1586
rect 336 1505 360 1539
rect 394 1505 418 1539
rect 336 1469 418 1505
rect 13152 1547 13194 1581
rect 13228 1547 13264 1581
rect 13298 1547 13334 1581
rect 13368 1547 13404 1581
rect 13438 1547 13474 1581
rect 13508 1547 13544 1581
rect 13578 1547 13614 1581
rect 13648 1547 13684 1581
rect 13718 1547 13754 1581
rect 13788 1547 13824 1581
rect 13858 1547 13894 1581
rect 13928 1547 13964 1581
rect 13998 1547 14034 1581
rect 14068 1547 14104 1581
rect 14138 1547 14174 1581
rect 14208 1547 14244 1581
rect 14278 1547 14314 1581
rect 14348 1547 14384 1581
rect 14418 1547 14454 1581
rect 14488 1547 14524 1581
rect 14558 1547 14594 1581
rect 14628 1547 14664 1581
rect 14698 1552 14774 1581
rect 14808 1552 14844 1586
rect 14878 1552 14914 1586
rect 14948 1552 14984 1586
rect 15018 1552 15054 1586
rect 15088 1552 15124 1586
rect 15158 1552 15194 1586
rect 15228 1552 15264 1586
rect 15298 1552 15334 1586
rect 15368 1552 15404 1586
rect 15438 1552 15474 1586
rect 15508 1552 15544 1586
rect 15578 1552 15614 1586
rect 15648 1552 15684 1586
rect 15718 1552 15754 1586
rect 15788 1552 15824 1586
rect 15858 1552 15894 1586
rect 15928 1552 15964 1586
rect 15998 1552 16032 1586
rect 14698 1547 16032 1552
rect 13152 1518 16032 1547
rect 13152 1511 14774 1518
rect 336 1435 360 1469
rect 394 1435 418 1469
rect 336 1399 418 1435
rect 336 1365 360 1399
rect 394 1365 418 1399
rect 13152 1477 13194 1511
rect 13228 1477 13264 1511
rect 13298 1477 13334 1511
rect 13368 1477 13404 1511
rect 13438 1477 13474 1511
rect 13508 1477 13544 1511
rect 13578 1477 13614 1511
rect 13648 1477 13684 1511
rect 13718 1477 13754 1511
rect 13788 1477 13824 1511
rect 13858 1477 13894 1511
rect 13928 1477 13964 1511
rect 13998 1477 14034 1511
rect 14068 1477 14104 1511
rect 14138 1477 14174 1511
rect 14208 1477 14244 1511
rect 14278 1477 14314 1511
rect 14348 1477 14384 1511
rect 14418 1477 14454 1511
rect 14488 1477 14524 1511
rect 14558 1477 14594 1511
rect 14628 1477 14664 1511
rect 14698 1484 14774 1511
rect 14808 1484 14844 1518
rect 14878 1484 14914 1518
rect 14948 1484 14984 1518
rect 15018 1484 15054 1518
rect 15088 1484 15124 1518
rect 15158 1484 15194 1518
rect 15228 1484 15264 1518
rect 15298 1484 15334 1518
rect 15368 1484 15404 1518
rect 15438 1484 15474 1518
rect 15508 1484 15544 1518
rect 15578 1484 15614 1518
rect 15648 1484 15684 1518
rect 15718 1484 15754 1518
rect 15788 1484 15824 1518
rect 15858 1484 15894 1518
rect 15928 1484 15964 1518
rect 15998 1484 16032 1518
rect 14698 1477 16032 1484
rect 13152 1450 16032 1477
rect 13152 1441 14774 1450
rect 13152 1407 13194 1441
rect 13228 1407 13264 1441
rect 13298 1407 13334 1441
rect 13368 1407 13404 1441
rect 13438 1407 13474 1441
rect 13508 1407 13544 1441
rect 13578 1407 13614 1441
rect 13648 1407 13684 1441
rect 13718 1407 13754 1441
rect 13788 1407 13824 1441
rect 13858 1407 13894 1441
rect 13928 1407 13964 1441
rect 13998 1407 14034 1441
rect 14068 1407 14104 1441
rect 14138 1407 14174 1441
rect 14208 1407 14244 1441
rect 14278 1407 14314 1441
rect 14348 1407 14384 1441
rect 14418 1407 14454 1441
rect 14488 1407 14524 1441
rect 14558 1407 14594 1441
rect 14628 1407 14664 1441
rect 14698 1416 14774 1441
rect 14808 1416 14844 1450
rect 14878 1416 14914 1450
rect 14948 1416 14984 1450
rect 15018 1416 15054 1450
rect 15088 1416 15124 1450
rect 15158 1416 15194 1450
rect 15228 1416 15264 1450
rect 15298 1416 15334 1450
rect 15368 1416 15404 1450
rect 15438 1416 15474 1450
rect 15508 1416 15544 1450
rect 15578 1416 15614 1450
rect 15648 1416 15684 1450
rect 15718 1416 15754 1450
rect 15788 1416 15824 1450
rect 15858 1416 15894 1450
rect 15928 1416 15964 1450
rect 15998 1416 16032 1450
rect 14698 1407 16032 1416
rect 336 1329 418 1365
rect 13152 1382 16032 1407
rect 13152 1371 14774 1382
rect 336 1295 360 1329
rect 394 1295 418 1329
rect 336 1259 418 1295
rect 336 1225 360 1259
rect 394 1225 418 1259
rect 13152 1337 13194 1371
rect 13228 1337 13264 1371
rect 13298 1337 13334 1371
rect 13368 1337 13404 1371
rect 13438 1337 13474 1371
rect 13508 1337 13544 1371
rect 13578 1337 13614 1371
rect 13648 1337 13684 1371
rect 13718 1337 13754 1371
rect 13788 1337 13824 1371
rect 13858 1337 13894 1371
rect 13928 1337 13964 1371
rect 13998 1337 14034 1371
rect 14068 1337 14104 1371
rect 14138 1337 14174 1371
rect 14208 1337 14244 1371
rect 14278 1337 14314 1371
rect 14348 1337 14384 1371
rect 14418 1337 14454 1371
rect 14488 1337 14524 1371
rect 14558 1337 14594 1371
rect 14628 1337 14664 1371
rect 14698 1348 14774 1371
rect 14808 1348 14844 1382
rect 14878 1348 14914 1382
rect 14948 1348 14984 1382
rect 15018 1348 15054 1382
rect 15088 1348 15124 1382
rect 15158 1348 15194 1382
rect 15228 1348 15264 1382
rect 15298 1348 15334 1382
rect 15368 1348 15404 1382
rect 15438 1348 15474 1382
rect 15508 1348 15544 1382
rect 15578 1348 15614 1382
rect 15648 1348 15684 1382
rect 15718 1348 15754 1382
rect 15788 1348 15824 1382
rect 15858 1348 15894 1382
rect 15928 1348 15964 1382
rect 15998 1348 16032 1382
rect 14698 1337 16032 1348
rect 13152 1314 16032 1337
rect 13152 1301 14774 1314
rect 13152 1267 13194 1301
rect 13228 1267 13264 1301
rect 13298 1267 13334 1301
rect 13368 1267 13404 1301
rect 13438 1267 13474 1301
rect 13508 1267 13544 1301
rect 13578 1267 13614 1301
rect 13648 1267 13684 1301
rect 13718 1267 13754 1301
rect 13788 1267 13824 1301
rect 13858 1267 13894 1301
rect 13928 1267 13964 1301
rect 13998 1267 14034 1301
rect 14068 1267 14104 1301
rect 14138 1267 14174 1301
rect 14208 1267 14244 1301
rect 14278 1267 14314 1301
rect 14348 1267 14384 1301
rect 14418 1267 14454 1301
rect 14488 1267 14524 1301
rect 14558 1267 14594 1301
rect 14628 1267 14664 1301
rect 14698 1280 14774 1301
rect 14808 1280 14844 1314
rect 14878 1280 14914 1314
rect 14948 1280 14984 1314
rect 15018 1280 15054 1314
rect 15088 1280 15124 1314
rect 15158 1280 15194 1314
rect 15228 1280 15264 1314
rect 15298 1280 15334 1314
rect 15368 1280 15404 1314
rect 15438 1280 15474 1314
rect 15508 1280 15544 1314
rect 15578 1280 15614 1314
rect 15648 1280 15684 1314
rect 15718 1280 15754 1314
rect 15788 1280 15824 1314
rect 15858 1280 15894 1314
rect 15928 1280 15964 1314
rect 15998 1280 16032 1314
rect 14698 1267 16032 1280
rect 13152 1246 16032 1267
rect 336 1189 418 1225
rect 336 1155 360 1189
rect 394 1155 418 1189
rect 13152 1231 14774 1246
rect 13152 1197 13194 1231
rect 13228 1197 13264 1231
rect 13298 1197 13334 1231
rect 13368 1197 13404 1231
rect 13438 1197 13474 1231
rect 13508 1197 13544 1231
rect 13578 1197 13614 1231
rect 13648 1197 13684 1231
rect 13718 1197 13754 1231
rect 13788 1197 13824 1231
rect 13858 1197 13894 1231
rect 13928 1197 13964 1231
rect 13998 1197 14034 1231
rect 14068 1197 14104 1231
rect 14138 1197 14174 1231
rect 14208 1197 14244 1231
rect 14278 1197 14314 1231
rect 14348 1197 14384 1231
rect 14418 1197 14454 1231
rect 14488 1197 14524 1231
rect 14558 1197 14594 1231
rect 14628 1197 14664 1231
rect 14698 1212 14774 1231
rect 14808 1212 14844 1246
rect 14878 1212 14914 1246
rect 14948 1212 14984 1246
rect 15018 1212 15054 1246
rect 15088 1212 15124 1246
rect 15158 1212 15194 1246
rect 15228 1212 15264 1246
rect 15298 1212 15334 1246
rect 15368 1212 15404 1246
rect 15438 1212 15474 1246
rect 15508 1212 15544 1246
rect 15578 1212 15614 1246
rect 15648 1212 15684 1246
rect 15718 1212 15754 1246
rect 15788 1212 15824 1246
rect 15858 1212 15894 1246
rect 15928 1212 15964 1246
rect 15998 1212 16032 1246
rect 14698 1197 16032 1212
rect 336 1119 418 1155
rect 336 1085 360 1119
rect 394 1085 418 1119
rect 13152 1178 16032 1197
rect 13152 1161 14774 1178
rect 13152 1127 13194 1161
rect 13228 1127 13264 1161
rect 13298 1127 13334 1161
rect 13368 1127 13404 1161
rect 13438 1127 13474 1161
rect 13508 1127 13544 1161
rect 13578 1127 13614 1161
rect 13648 1127 13684 1161
rect 13718 1127 13754 1161
rect 13788 1127 13824 1161
rect 13858 1127 13894 1161
rect 13928 1127 13964 1161
rect 13998 1127 14034 1161
rect 14068 1127 14104 1161
rect 14138 1127 14174 1161
rect 14208 1127 14244 1161
rect 14278 1127 14314 1161
rect 14348 1127 14384 1161
rect 14418 1127 14454 1161
rect 14488 1127 14524 1161
rect 14558 1127 14594 1161
rect 14628 1127 14664 1161
rect 14698 1144 14774 1161
rect 14808 1144 14844 1178
rect 14878 1144 14914 1178
rect 14948 1144 14984 1178
rect 15018 1144 15054 1178
rect 15088 1144 15124 1178
rect 15158 1144 15194 1178
rect 15228 1144 15264 1178
rect 15298 1144 15334 1178
rect 15368 1144 15404 1178
rect 15438 1144 15474 1178
rect 15508 1144 15544 1178
rect 15578 1144 15614 1178
rect 15648 1144 15684 1178
rect 15718 1144 15754 1178
rect 15788 1144 15824 1178
rect 15858 1144 15894 1178
rect 15928 1144 15964 1178
rect 15998 1144 16032 1178
rect 14698 1127 16032 1144
rect 13152 1110 16032 1127
rect 13152 1091 14774 1110
rect 336 1050 418 1085
rect 336 1016 360 1050
rect 394 1016 418 1050
rect 13152 1057 13194 1091
rect 13228 1057 13264 1091
rect 13298 1057 13334 1091
rect 13368 1057 13404 1091
rect 13438 1057 13474 1091
rect 13508 1057 13544 1091
rect 13578 1057 13614 1091
rect 13648 1057 13684 1091
rect 13718 1057 13754 1091
rect 13788 1057 13824 1091
rect 13858 1057 13894 1091
rect 13928 1057 13964 1091
rect 13998 1057 14034 1091
rect 14068 1057 14104 1091
rect 14138 1057 14174 1091
rect 14208 1057 14244 1091
rect 14278 1057 14314 1091
rect 14348 1057 14384 1091
rect 14418 1057 14454 1091
rect 14488 1057 14524 1091
rect 14558 1057 14594 1091
rect 14628 1057 14664 1091
rect 14698 1076 14774 1091
rect 14808 1076 14844 1110
rect 14878 1076 14914 1110
rect 14948 1076 14984 1110
rect 15018 1076 15054 1110
rect 15088 1076 15124 1110
rect 15158 1076 15194 1110
rect 15228 1076 15264 1110
rect 15298 1076 15334 1110
rect 15368 1076 15404 1110
rect 15438 1076 15474 1110
rect 15508 1076 15544 1110
rect 15578 1076 15614 1110
rect 15648 1076 15684 1110
rect 15718 1076 15754 1110
rect 15788 1076 15824 1110
rect 15858 1076 15894 1110
rect 15928 1076 15964 1110
rect 15998 1076 16032 1110
rect 14698 1057 16032 1076
rect 13152 1042 16032 1057
rect 336 981 418 1016
rect 336 947 360 981
rect 394 947 418 981
rect 336 912 418 947
rect 13152 1021 14774 1042
rect 13152 987 13194 1021
rect 13228 987 13264 1021
rect 13298 987 13334 1021
rect 13368 987 13404 1021
rect 13438 987 13474 1021
rect 13508 987 13544 1021
rect 13578 987 13614 1021
rect 13648 987 13684 1021
rect 13718 987 13754 1021
rect 13788 987 13824 1021
rect 13858 987 13894 1021
rect 13928 987 13964 1021
rect 13998 987 14034 1021
rect 14068 987 14104 1021
rect 14138 987 14174 1021
rect 14208 987 14244 1021
rect 14278 987 14314 1021
rect 14348 987 14384 1021
rect 14418 987 14454 1021
rect 14488 987 14524 1021
rect 14558 987 14594 1021
rect 14628 987 14664 1021
rect 14698 1008 14774 1021
rect 14808 1008 14844 1042
rect 14878 1008 14914 1042
rect 14948 1008 14984 1042
rect 15018 1008 15054 1042
rect 15088 1008 15124 1042
rect 15158 1008 15194 1042
rect 15228 1008 15264 1042
rect 15298 1008 15334 1042
rect 15368 1008 15404 1042
rect 15438 1008 15474 1042
rect 15508 1008 15544 1042
rect 15578 1008 15614 1042
rect 15648 1008 15684 1042
rect 15718 1008 15754 1042
rect 15788 1008 15824 1042
rect 15858 1008 15894 1042
rect 15928 1008 15964 1042
rect 15998 1008 16032 1042
rect 14698 987 16032 1008
rect 13152 974 16032 987
rect 13152 951 14774 974
rect 336 878 360 912
rect 394 878 418 912
rect 13152 917 13194 951
rect 13228 917 13264 951
rect 13298 917 13334 951
rect 13368 917 13404 951
rect 13438 917 13474 951
rect 13508 917 13544 951
rect 13578 917 13614 951
rect 13648 917 13684 951
rect 13718 917 13754 951
rect 13788 917 13824 951
rect 13858 917 13894 951
rect 13928 917 13964 951
rect 13998 917 14034 951
rect 14068 917 14104 951
rect 14138 917 14174 951
rect 14208 917 14244 951
rect 14278 917 14314 951
rect 14348 917 14384 951
rect 14418 917 14454 951
rect 14488 917 14524 951
rect 14558 917 14594 951
rect 14628 917 14664 951
rect 14698 940 14774 951
rect 14808 940 14844 974
rect 14878 940 14914 974
rect 14948 940 14984 974
rect 15018 940 15054 974
rect 15088 940 15124 974
rect 15158 940 15194 974
rect 15228 940 15264 974
rect 15298 940 15334 974
rect 15368 940 15404 974
rect 15438 940 15474 974
rect 15508 940 15544 974
rect 15578 940 15614 974
rect 15648 940 15684 974
rect 15718 940 15754 974
rect 15788 940 15824 974
rect 15858 940 15894 974
rect 15928 940 15964 974
rect 15998 940 16032 974
rect 14698 917 16032 940
rect 13152 906 16032 917
rect 13152 881 14774 906
rect 336 843 418 878
rect 336 809 360 843
rect 394 809 418 843
rect 336 774 418 809
rect 13152 847 13194 881
rect 13228 847 13264 881
rect 13298 847 13334 881
rect 13368 847 13404 881
rect 13438 847 13474 881
rect 13508 847 13544 881
rect 13578 847 13614 881
rect 13648 847 13684 881
rect 13718 847 13754 881
rect 13788 847 13824 881
rect 13858 847 13894 881
rect 13928 847 13964 881
rect 13998 847 14034 881
rect 14068 847 14104 881
rect 14138 847 14174 881
rect 14208 847 14244 881
rect 14278 847 14314 881
rect 14348 847 14384 881
rect 14418 847 14454 881
rect 14488 847 14524 881
rect 14558 847 14594 881
rect 14628 847 14664 881
rect 14698 872 14774 881
rect 14808 872 14844 906
rect 14878 872 14914 906
rect 14948 872 14984 906
rect 15018 872 15054 906
rect 15088 872 15124 906
rect 15158 872 15194 906
rect 15228 872 15264 906
rect 15298 872 15334 906
rect 15368 872 15404 906
rect 15438 872 15474 906
rect 15508 872 15544 906
rect 15578 872 15614 906
rect 15648 872 15684 906
rect 15718 872 15754 906
rect 15788 872 15824 906
rect 15858 872 15894 906
rect 15928 872 15964 906
rect 15998 872 16032 906
rect 14698 847 16032 872
rect 13152 838 16032 847
rect 13152 811 14774 838
rect 336 740 360 774
rect 394 740 418 774
rect 336 705 418 740
rect 13152 777 13194 811
rect 13228 777 13264 811
rect 13298 777 13334 811
rect 13368 777 13404 811
rect 13438 777 13474 811
rect 13508 777 13544 811
rect 13578 777 13614 811
rect 13648 777 13684 811
rect 13718 777 13754 811
rect 13788 777 13824 811
rect 13858 777 13894 811
rect 13928 777 13964 811
rect 13998 777 14034 811
rect 14068 777 14104 811
rect 14138 777 14174 811
rect 14208 777 14244 811
rect 14278 777 14314 811
rect 14348 777 14384 811
rect 14418 777 14454 811
rect 14488 777 14524 811
rect 14558 777 14594 811
rect 14628 777 14664 811
rect 14698 804 14774 811
rect 14808 804 14844 838
rect 14878 804 14914 838
rect 14948 804 14984 838
rect 15018 804 15054 838
rect 15088 804 15124 838
rect 15158 804 15194 838
rect 15228 804 15264 838
rect 15298 804 15334 838
rect 15368 804 15404 838
rect 15438 804 15474 838
rect 15508 804 15544 838
rect 15578 804 15614 838
rect 15648 804 15684 838
rect 15718 804 15754 838
rect 15788 804 15824 838
rect 15858 804 15894 838
rect 15928 804 15964 838
rect 15998 804 16032 838
rect 14698 777 16032 804
rect 13152 770 16032 777
rect 13152 741 14774 770
rect 336 671 360 705
rect 394 671 418 705
rect 336 636 418 671
rect 336 602 360 636
rect 394 602 418 636
rect 13152 707 13194 741
rect 13228 707 13264 741
rect 13298 707 13334 741
rect 13368 707 13404 741
rect 13438 707 13474 741
rect 13508 707 13544 741
rect 13578 707 13614 741
rect 13648 707 13684 741
rect 13718 707 13754 741
rect 13788 707 13824 741
rect 13858 707 13894 741
rect 13928 707 13964 741
rect 13998 707 14034 741
rect 14068 707 14104 741
rect 14138 707 14174 741
rect 14208 707 14244 741
rect 14278 707 14314 741
rect 14348 707 14384 741
rect 14418 707 14454 741
rect 14488 707 14524 741
rect 14558 707 14594 741
rect 14628 707 14664 741
rect 14698 736 14774 741
rect 14808 736 14844 770
rect 14878 736 14914 770
rect 14948 736 14984 770
rect 15018 736 15054 770
rect 15088 736 15124 770
rect 15158 736 15194 770
rect 15228 736 15264 770
rect 15298 736 15334 770
rect 15368 736 15404 770
rect 15438 736 15474 770
rect 15508 736 15544 770
rect 15578 736 15614 770
rect 15648 736 15684 770
rect 15718 736 15754 770
rect 15788 736 15824 770
rect 15858 736 15894 770
rect 15928 736 15964 770
rect 15998 736 16032 770
rect 14698 707 16032 736
rect 13152 702 16032 707
rect 13152 671 14774 702
rect 13152 637 13194 671
rect 13228 637 13264 671
rect 13298 637 13334 671
rect 13368 637 13404 671
rect 13438 637 13474 671
rect 13508 637 13544 671
rect 13578 637 13614 671
rect 13648 637 13684 671
rect 13718 637 13754 671
rect 13788 637 13824 671
rect 13858 637 13894 671
rect 13928 637 13964 671
rect 13998 637 14034 671
rect 14068 637 14104 671
rect 14138 637 14174 671
rect 14208 637 14244 671
rect 14278 637 14314 671
rect 14348 637 14384 671
rect 14418 637 14454 671
rect 14488 637 14524 671
rect 14558 637 14594 671
rect 14628 637 14664 671
rect 14698 668 14774 671
rect 14808 668 14844 702
rect 14878 668 14914 702
rect 14948 668 14984 702
rect 15018 668 15054 702
rect 15088 668 15124 702
rect 15158 668 15194 702
rect 15228 668 15264 702
rect 15298 668 15334 702
rect 15368 668 15404 702
rect 15438 668 15474 702
rect 15508 668 15544 702
rect 15578 668 15614 702
rect 15648 668 15684 702
rect 15718 668 15754 702
rect 15788 668 15824 702
rect 15858 668 15894 702
rect 15928 668 15964 702
rect 15998 668 16032 702
rect 14698 637 16032 668
rect 13152 634 16032 637
rect 336 567 418 602
rect 13152 601 14774 634
rect 336 533 360 567
rect 394 533 418 567
rect 336 498 418 533
rect 336 464 360 498
rect 394 464 418 498
rect 13152 567 13194 601
rect 13228 567 13264 601
rect 13298 567 13334 601
rect 13368 567 13404 601
rect 13438 567 13474 601
rect 13508 567 13544 601
rect 13578 567 13614 601
rect 13648 567 13684 601
rect 13718 567 13754 601
rect 13788 567 13824 601
rect 13858 567 13894 601
rect 13928 567 13964 601
rect 13998 567 14034 601
rect 14068 567 14104 601
rect 14138 567 14174 601
rect 14208 567 14244 601
rect 14278 567 14314 601
rect 14348 567 14384 601
rect 14418 567 14454 601
rect 14488 567 14524 601
rect 14558 567 14594 601
rect 14628 567 14664 601
rect 14698 600 14774 601
rect 14808 600 14844 634
rect 14878 600 14914 634
rect 14948 600 14984 634
rect 15018 600 15054 634
rect 15088 600 15124 634
rect 15158 600 15194 634
rect 15228 600 15264 634
rect 15298 600 15334 634
rect 15368 600 15404 634
rect 15438 600 15474 634
rect 15508 600 15544 634
rect 15578 600 15614 634
rect 15648 600 15684 634
rect 15718 600 15754 634
rect 15788 600 15824 634
rect 15858 600 15894 634
rect 15928 600 15964 634
rect 15998 600 16032 634
rect 14698 567 16032 600
rect 13152 566 16032 567
rect 13152 532 14774 566
rect 14808 532 14844 566
rect 14878 532 14914 566
rect 14948 532 14984 566
rect 15018 532 15054 566
rect 15088 532 15124 566
rect 15158 532 15194 566
rect 15228 532 15264 566
rect 15298 532 15334 566
rect 15368 532 15404 566
rect 15438 532 15474 566
rect 15508 532 15544 566
rect 15578 532 15614 566
rect 15648 532 15684 566
rect 15718 532 15754 566
rect 15788 532 15824 566
rect 15858 532 15894 566
rect 15928 532 15964 566
rect 15998 532 16032 566
rect 13152 531 16032 532
rect 13152 497 13194 531
rect 13228 497 13264 531
rect 13298 497 13334 531
rect 13368 497 13404 531
rect 13438 497 13474 531
rect 13508 497 13544 531
rect 13578 497 13614 531
rect 13648 497 13684 531
rect 13718 497 13754 531
rect 13788 497 13824 531
rect 13858 497 13894 531
rect 13928 497 13964 531
rect 13998 497 14034 531
rect 14068 497 14104 531
rect 14138 497 14174 531
rect 14208 497 14244 531
rect 14278 497 14314 531
rect 14348 497 14384 531
rect 14418 497 14454 531
rect 14488 497 14524 531
rect 14558 497 14594 531
rect 14628 497 14664 531
rect 14698 498 16032 531
rect 14698 497 14774 498
rect 336 429 418 464
rect 336 395 360 429
rect 394 395 418 429
rect 13152 464 14774 497
rect 14808 464 14844 498
rect 14878 464 14914 498
rect 14948 464 14984 498
rect 15018 464 15054 498
rect 15088 464 15124 498
rect 15158 464 15194 498
rect 15228 464 15264 498
rect 15298 464 15334 498
rect 15368 464 15404 498
rect 15438 464 15474 498
rect 15508 464 15544 498
rect 15578 464 15614 498
rect 15648 464 15684 498
rect 15718 464 15754 498
rect 15788 464 15824 498
rect 15858 464 15894 498
rect 15928 464 15964 498
rect 15998 464 16032 498
rect 13152 461 16032 464
rect 13152 427 13194 461
rect 13228 427 13264 461
rect 13298 427 13334 461
rect 13368 427 13404 461
rect 13438 427 13474 461
rect 13508 427 13544 461
rect 13578 427 13614 461
rect 13648 427 13684 461
rect 13718 427 13754 461
rect 13788 427 13824 461
rect 13858 427 13894 461
rect 13928 427 13964 461
rect 13998 427 14034 461
rect 14068 427 14104 461
rect 14138 427 14174 461
rect 14208 427 14244 461
rect 14278 427 14314 461
rect 14348 427 14384 461
rect 14418 427 14454 461
rect 14488 427 14524 461
rect 14558 427 14594 461
rect 14628 427 14664 461
rect 14698 430 16032 461
rect 14698 427 14774 430
rect 336 360 418 395
rect 336 326 360 360
rect 394 326 418 360
rect 336 291 418 326
rect 13152 396 14774 427
rect 14808 396 14844 430
rect 14878 396 14914 430
rect 14948 396 14984 430
rect 15018 396 15054 430
rect 15088 396 15124 430
rect 15158 396 15194 430
rect 15228 396 15264 430
rect 15298 396 15334 430
rect 15368 396 15404 430
rect 15438 396 15474 430
rect 15508 396 15544 430
rect 15578 396 15614 430
rect 15648 396 15684 430
rect 15718 396 15754 430
rect 15788 396 15824 430
rect 15858 396 15894 430
rect 15928 396 15964 430
rect 15998 396 16032 430
rect 13152 391 16032 396
rect 13152 357 13194 391
rect 13228 357 13264 391
rect 13298 357 13334 391
rect 13368 357 13404 391
rect 13438 357 13474 391
rect 13508 357 13544 391
rect 13578 357 13614 391
rect 13648 357 13684 391
rect 13718 357 13754 391
rect 13788 357 13824 391
rect 13858 357 13894 391
rect 13928 357 13964 391
rect 13998 357 14034 391
rect 14068 357 14104 391
rect 14138 357 14174 391
rect 14208 357 14244 391
rect 14278 357 14314 391
rect 14348 357 14384 391
rect 14418 357 14454 391
rect 14488 357 14524 391
rect 14558 357 14594 391
rect 14628 357 14664 391
rect 14698 362 16032 391
rect 14698 357 14774 362
rect 13152 328 14774 357
rect 14808 328 14844 362
rect 14878 328 14914 362
rect 14948 328 14984 362
rect 15018 328 15054 362
rect 15088 328 15124 362
rect 15158 328 15194 362
rect 15228 328 15264 362
rect 15298 328 15334 362
rect 15368 328 15404 362
rect 15438 328 15474 362
rect 15508 328 15544 362
rect 15578 328 15614 362
rect 15648 328 15684 362
rect 15718 328 15754 362
rect 15788 328 15824 362
rect 15858 328 15894 362
rect 15928 328 15964 362
rect 15998 328 16032 362
rect 13152 321 16032 328
rect 336 257 360 291
rect 394 257 418 291
rect 13152 287 13194 321
rect 13228 287 13264 321
rect 13298 287 13334 321
rect 13368 287 13404 321
rect 13438 287 13474 321
rect 13508 287 13544 321
rect 13578 287 13614 321
rect 13648 287 13684 321
rect 13718 287 13754 321
rect 13788 287 13824 321
rect 13858 287 13894 321
rect 13928 287 13964 321
rect 13998 287 14034 321
rect 14068 287 14104 321
rect 14138 287 14174 321
rect 14208 287 14244 321
rect 14278 287 14314 321
rect 14348 287 14384 321
rect 14418 287 14454 321
rect 14488 287 14524 321
rect 14558 287 14594 321
rect 14628 287 14664 321
rect 14698 294 16032 321
rect 14698 287 14774 294
rect 336 222 418 257
rect 336 188 360 222
rect 394 188 418 222
rect 336 153 418 188
rect 13152 260 14774 287
rect 14808 260 14844 294
rect 14878 260 14914 294
rect 14948 260 14984 294
rect 15018 260 15054 294
rect 15088 260 15124 294
rect 15158 260 15194 294
rect 15228 260 15264 294
rect 15298 260 15334 294
rect 15368 260 15404 294
rect 15438 260 15474 294
rect 15508 260 15544 294
rect 15578 260 15614 294
rect 15648 260 15684 294
rect 15718 260 15754 294
rect 15788 260 15824 294
rect 15858 260 15894 294
rect 15928 260 15964 294
rect 15998 260 16032 294
rect 13152 251 16032 260
rect 13152 217 13194 251
rect 13228 217 13264 251
rect 13298 217 13334 251
rect 13368 217 13404 251
rect 13438 217 13474 251
rect 13508 217 13544 251
rect 13578 217 13614 251
rect 13648 217 13684 251
rect 13718 217 13754 251
rect 13788 217 13824 251
rect 13858 217 13894 251
rect 13928 217 13964 251
rect 13998 217 14034 251
rect 14068 217 14104 251
rect 14138 217 14174 251
rect 14208 217 14244 251
rect 14278 217 14314 251
rect 14348 217 14384 251
rect 14418 217 14454 251
rect 14488 217 14524 251
rect 14558 217 14594 251
rect 14628 217 14664 251
rect 14698 226 16032 251
rect 14698 217 14774 226
rect 13152 192 14774 217
rect 14808 192 14844 226
rect 14878 192 14914 226
rect 14948 192 14984 226
rect 15018 192 15054 226
rect 15088 192 15124 226
rect 15158 192 15194 226
rect 15228 192 15264 226
rect 15298 192 15334 226
rect 15368 192 15404 226
rect 15438 192 15474 226
rect 15508 192 15544 226
rect 15578 192 15614 226
rect 15648 192 15684 226
rect 15718 192 15754 226
rect 15788 192 15824 226
rect 15858 192 15894 226
rect 15928 192 15964 226
rect 15998 192 16032 226
rect 13152 181 16032 192
rect 336 119 360 153
rect 394 119 418 153
rect 336 108 418 119
rect 13152 147 13194 181
rect 13228 147 13264 181
rect 13298 147 13334 181
rect 13368 147 13404 181
rect 13438 147 13474 181
rect 13508 147 13544 181
rect 13578 147 13614 181
rect 13648 147 13684 181
rect 13718 147 13754 181
rect 13788 147 13824 181
rect 13858 147 13894 181
rect 13928 147 13964 181
rect 13998 147 14034 181
rect 14068 147 14104 181
rect 14138 147 14174 181
rect 14208 147 14244 181
rect 14278 147 14314 181
rect 14348 147 14384 181
rect 14418 147 14454 181
rect 14488 147 14524 181
rect 14558 147 14594 181
rect 14628 147 14664 181
rect 14698 158 16032 181
rect 14698 147 14774 158
rect 13152 124 14774 147
rect 14808 124 14844 158
rect 14878 124 14914 158
rect 14948 124 14984 158
rect 15018 124 15054 158
rect 15088 124 15124 158
rect 15158 124 15194 158
rect 15228 124 15264 158
rect 15298 124 15334 158
rect 15368 124 15404 158
rect 15438 124 15474 158
rect 15508 124 15544 158
rect 15578 124 15614 158
rect 15648 124 15684 158
rect 15718 124 15754 158
rect 15788 124 15824 158
rect 15858 124 15894 158
rect 15928 124 15964 158
rect 15998 124 16032 158
rect 13152 108 16032 124
rect 336 84 16032 108
rect 336 50 360 84
rect 394 50 429 84
rect 463 50 498 84
rect 532 50 567 84
rect 601 50 636 84
rect 670 50 705 84
rect 739 50 774 84
rect 808 50 843 84
rect 877 50 912 84
rect 946 50 981 84
rect 1015 50 1050 84
rect 1084 50 1119 84
rect 1153 50 1188 84
rect 1222 50 1257 84
rect 1291 50 1326 84
rect 1360 50 1395 84
rect 1429 50 1464 84
rect 1498 50 1533 84
rect 1567 50 1602 84
rect 1636 50 1671 84
rect 1705 50 1740 84
rect 1774 50 1809 84
rect 1843 50 1878 84
rect 1912 50 1947 84
rect 1981 50 2016 84
rect 2050 50 2085 84
rect 2119 50 2154 84
rect 2188 50 2223 84
rect 2257 50 2292 84
rect 2326 50 2361 84
rect 2395 50 2430 84
rect 2464 50 2499 84
rect 2533 50 2568 84
rect 2602 50 2637 84
rect 2671 50 2706 84
rect 2740 50 2775 84
rect 2809 50 2844 84
rect 2878 50 2913 84
rect 2947 50 2982 84
rect 3016 50 3051 84
rect 3085 50 3120 84
rect 3154 50 3189 84
rect 3223 50 3258 84
rect 3292 50 3327 84
rect 3361 50 3396 84
rect 3430 50 3465 84
rect 3499 50 3534 84
rect 3568 50 3603 84
rect 3637 50 3672 84
rect 3706 50 3741 84
rect 3775 50 3810 84
rect 3844 50 3879 84
rect 3913 50 3948 84
rect 3982 50 4017 84
rect 4051 50 4086 84
rect 4120 50 4155 84
rect 4189 50 4224 84
rect 4258 50 4293 84
rect 4327 50 4362 84
rect 4396 50 4431 84
rect 4465 50 4500 84
rect 4534 50 4569 84
rect 4603 50 4638 84
rect 4672 50 4707 84
rect 4741 50 4776 84
rect 4810 50 4845 84
rect 4879 50 4914 84
rect 4948 50 4982 84
rect 5016 50 5050 84
rect 5084 50 5118 84
rect 5152 50 5186 84
rect 5220 50 5254 84
rect 5288 50 5322 84
rect 5356 50 5390 84
rect 5424 50 5458 84
rect 5492 50 5526 84
rect 5560 50 5594 84
rect 5628 50 5662 84
rect 5696 50 5730 84
rect 5764 50 5798 84
rect 5832 50 5866 84
rect 5900 50 5934 84
rect 5968 50 6002 84
rect 6036 50 6070 84
rect 6104 50 6138 84
rect 6172 50 6206 84
rect 6240 50 6274 84
rect 6308 50 6342 84
rect 6376 50 6410 84
rect 6444 50 6478 84
rect 6512 50 6546 84
rect 6580 50 6614 84
rect 6648 50 6682 84
rect 6716 50 6750 84
rect 6784 50 6818 84
rect 6852 50 6886 84
rect 6920 50 6954 84
rect 6988 50 7022 84
rect 7056 50 7090 84
rect 7124 50 7158 84
rect 7192 50 7226 84
rect 7260 50 7294 84
rect 7328 50 7362 84
rect 7396 50 7430 84
rect 7464 50 7498 84
rect 7532 50 7566 84
rect 7600 50 7634 84
rect 7668 50 7702 84
rect 7736 50 7770 84
rect 7804 50 7838 84
rect 7872 50 7906 84
rect 7940 50 7974 84
rect 8008 50 8042 84
rect 8076 50 8110 84
rect 8144 50 8178 84
rect 8212 50 8246 84
rect 8280 50 8314 84
rect 8348 50 8382 84
rect 8416 50 8450 84
rect 8484 50 8518 84
rect 8552 50 8586 84
rect 8620 50 8654 84
rect 8688 50 8722 84
rect 8756 50 8790 84
rect 8824 50 8858 84
rect 8892 50 8926 84
rect 8960 50 8994 84
rect 9028 50 9062 84
rect 9096 50 9130 84
rect 9164 50 9198 84
rect 9232 50 9266 84
rect 9300 50 9334 84
rect 9368 50 9402 84
rect 9436 50 9470 84
rect 9504 50 9538 84
rect 9572 50 9606 84
rect 9640 50 9674 84
rect 9708 50 9742 84
rect 9776 50 9810 84
rect 9844 50 9878 84
rect 9912 50 9946 84
rect 9980 50 10014 84
rect 10048 50 10082 84
rect 10116 50 10150 84
rect 10184 50 10218 84
rect 10252 50 10286 84
rect 10320 50 10354 84
rect 10388 50 10422 84
rect 10456 50 10490 84
rect 10524 50 10558 84
rect 10592 50 10626 84
rect 10660 50 10694 84
rect 10728 50 10762 84
rect 10796 50 10830 84
rect 10864 50 10898 84
rect 10932 50 10966 84
rect 11000 50 11034 84
rect 11068 50 11102 84
rect 11136 50 11170 84
rect 11204 50 11238 84
rect 11272 50 11306 84
rect 11340 50 11374 84
rect 11408 50 11442 84
rect 11476 50 11510 84
rect 11544 50 11578 84
rect 11612 50 11646 84
rect 11680 50 11714 84
rect 11748 50 11782 84
rect 11816 50 11850 84
rect 11884 50 11918 84
rect 11952 50 11986 84
rect 12020 50 12054 84
rect 12088 50 12122 84
rect 12156 50 12190 84
rect 12224 50 12258 84
rect 12292 50 12326 84
rect 12360 50 12394 84
rect 12428 50 12462 84
rect 12496 50 12530 84
rect 12564 50 12598 84
rect 12632 50 12666 84
rect 12700 50 12734 84
rect 12768 50 12802 84
rect 12836 50 12870 84
rect 12904 50 12938 84
rect 12972 50 13006 84
rect 13040 50 13074 84
rect 13108 50 13142 84
rect 13176 50 13210 84
rect 13244 50 13278 84
rect 13312 50 13346 84
rect 13380 50 13414 84
rect 13448 50 13482 84
rect 13516 50 13550 84
rect 13584 50 13618 84
rect 13652 50 13686 84
rect 13720 50 13754 84
rect 13788 50 13822 84
rect 13856 50 13890 84
rect 13924 50 13958 84
rect 13992 50 14026 84
rect 14060 50 14094 84
rect 14128 50 14162 84
rect 14196 50 14230 84
rect 14264 50 14298 84
rect 14332 50 14366 84
rect 14400 50 14434 84
rect 14468 50 14502 84
rect 14536 50 14570 84
rect 14604 50 14638 84
rect 14672 50 14706 84
rect 14740 50 14774 84
rect 14808 50 14842 84
rect 14876 50 14910 84
rect 14944 50 14978 84
rect 15012 50 15046 84
rect 15080 50 15114 84
rect 15148 50 15182 84
rect 15216 50 15250 84
rect 15284 50 15318 84
rect 15352 50 15386 84
rect 15420 50 15454 84
rect 15488 50 15522 84
rect 15556 50 15590 84
rect 15624 50 15658 84
rect 15692 50 15726 84
rect 15760 50 15794 84
rect 15828 50 15862 84
rect 15896 50 15930 84
rect 15964 50 15998 84
rect 336 26 16032 50
<< mvpsubdiff >>
rect 336 3909 10970 3933
rect 336 3906 470 3909
rect 336 3872 360 3906
rect 394 3875 470 3906
rect 504 3875 538 3909
rect 572 3875 606 3909
rect 640 3875 674 3909
rect 708 3875 742 3909
rect 776 3875 810 3909
rect 844 3875 878 3909
rect 912 3875 946 3909
rect 980 3875 1014 3909
rect 1048 3875 1082 3909
rect 1116 3875 1150 3909
rect 1184 3875 1218 3909
rect 1252 3875 1286 3909
rect 1320 3875 1354 3909
rect 1388 3875 1422 3909
rect 1456 3875 1490 3909
rect 1524 3875 1558 3909
rect 1592 3875 1626 3909
rect 1660 3875 1694 3909
rect 1728 3875 1762 3909
rect 1796 3875 1830 3909
rect 1864 3875 1898 3909
rect 1932 3875 1966 3909
rect 2000 3875 2034 3909
rect 2068 3875 2102 3909
rect 2136 3875 2170 3909
rect 2204 3875 2238 3909
rect 2272 3875 2306 3909
rect 2340 3875 2374 3909
rect 2408 3875 2442 3909
rect 2476 3875 2510 3909
rect 2544 3875 2578 3909
rect 2612 3875 2646 3909
rect 2680 3875 2714 3909
rect 2748 3875 2782 3909
rect 2816 3875 2850 3909
rect 2884 3875 2918 3909
rect 2952 3875 2986 3909
rect 3020 3875 3054 3909
rect 3088 3875 3122 3909
rect 3156 3875 3190 3909
rect 3224 3875 3258 3909
rect 3292 3875 3326 3909
rect 3360 3875 3394 3909
rect 3428 3875 3462 3909
rect 3496 3875 3530 3909
rect 3564 3875 3598 3909
rect 3632 3875 3666 3909
rect 3700 3875 3734 3909
rect 3768 3875 3802 3909
rect 3836 3875 3870 3909
rect 3904 3875 3938 3909
rect 3972 3875 4006 3909
rect 4040 3875 4074 3909
rect 4108 3875 4142 3909
rect 4176 3875 4210 3909
rect 4244 3875 4278 3909
rect 4312 3875 4346 3909
rect 4380 3875 4414 3909
rect 4448 3875 4482 3909
rect 4516 3875 4550 3909
rect 4584 3875 4618 3909
rect 4652 3875 4686 3909
rect 4720 3875 4754 3909
rect 4788 3875 4822 3909
rect 4856 3875 4890 3909
rect 4924 3875 4958 3909
rect 4992 3875 5026 3909
rect 5060 3875 5094 3909
rect 5128 3875 5162 3909
rect 5196 3875 5230 3909
rect 5264 3875 5298 3909
rect 5332 3875 5366 3909
rect 5400 3875 5434 3909
rect 5468 3875 5502 3909
rect 5536 3875 5570 3909
rect 5604 3875 5638 3909
rect 5672 3875 5706 3909
rect 5740 3875 5774 3909
rect 5808 3875 5842 3909
rect 5876 3875 5910 3909
rect 5944 3875 5978 3909
rect 6012 3875 6046 3909
rect 6080 3875 6114 3909
rect 6148 3875 6182 3909
rect 6216 3875 6250 3909
rect 6284 3875 6318 3909
rect 6352 3875 6386 3909
rect 6420 3875 6454 3909
rect 6488 3875 6522 3909
rect 6556 3875 6590 3909
rect 6624 3875 6658 3909
rect 6692 3875 6726 3909
rect 6760 3875 6794 3909
rect 6828 3875 6862 3909
rect 6896 3875 6930 3909
rect 6964 3875 6998 3909
rect 7032 3875 7066 3909
rect 7100 3875 7134 3909
rect 7168 3875 7202 3909
rect 7236 3875 7270 3909
rect 7304 3875 7338 3909
rect 7372 3875 7406 3909
rect 7440 3875 7474 3909
rect 7508 3875 7542 3909
rect 7576 3875 7610 3909
rect 7644 3875 7678 3909
rect 7712 3875 7746 3909
rect 7780 3875 7814 3909
rect 7848 3875 7882 3909
rect 7916 3875 7950 3909
rect 7984 3875 8018 3909
rect 8052 3875 8086 3909
rect 8120 3875 8154 3909
rect 8188 3875 8222 3909
rect 8256 3875 8290 3909
rect 8324 3875 8359 3909
rect 8393 3875 8428 3909
rect 8462 3875 8497 3909
rect 8531 3875 8566 3909
rect 8600 3875 8635 3909
rect 8669 3875 8704 3909
rect 8738 3875 8773 3909
rect 8807 3875 8842 3909
rect 8876 3875 8911 3909
rect 8945 3875 8980 3909
rect 9014 3875 9049 3909
rect 9083 3875 9118 3909
rect 9152 3875 9187 3909
rect 9221 3875 9256 3909
rect 9290 3875 9325 3909
rect 9359 3875 9394 3909
rect 9428 3875 9463 3909
rect 9497 3875 9532 3909
rect 9566 3875 9601 3909
rect 9635 3875 9670 3909
rect 9704 3875 9739 3909
rect 9773 3875 9808 3909
rect 9842 3875 9877 3909
rect 9911 3875 9946 3909
rect 9980 3875 10015 3909
rect 10049 3875 10084 3909
rect 10118 3875 10153 3909
rect 10187 3875 10222 3909
rect 10256 3875 10291 3909
rect 10325 3875 10360 3909
rect 10394 3875 10429 3909
rect 10463 3875 10498 3909
rect 10532 3875 10567 3909
rect 10601 3875 10636 3909
rect 10670 3875 10705 3909
rect 10739 3875 10774 3909
rect 10808 3875 10843 3909
rect 10877 3875 10912 3909
rect 10946 3875 10970 3909
rect 394 3872 10970 3875
rect 336 3851 10970 3872
rect 336 3835 418 3851
rect 336 3801 360 3835
rect 394 3801 418 3835
rect 10888 3839 10970 3851
rect 336 3764 418 3801
rect 336 3730 360 3764
rect 394 3730 418 3764
rect 336 3693 418 3730
rect 10888 3805 10912 3839
rect 10946 3805 10970 3839
rect 10888 3769 10970 3805
rect 10888 3735 10912 3769
rect 10946 3735 10970 3769
rect 336 3659 360 3693
rect 394 3659 418 3693
rect 336 3623 418 3659
rect 336 3589 360 3623
rect 394 3589 418 3623
rect 336 3553 418 3589
rect 336 3519 360 3553
rect 394 3519 418 3553
rect 336 3483 418 3519
rect 336 3449 360 3483
rect 394 3449 418 3483
rect 336 3413 418 3449
rect 336 3379 360 3413
rect 394 3379 418 3413
rect 336 3343 418 3379
rect 336 3309 360 3343
rect 394 3309 418 3343
rect 336 3273 418 3309
rect 336 3239 360 3273
rect 394 3239 418 3273
rect 336 3203 418 3239
rect 336 3169 360 3203
rect 394 3169 418 3203
rect 336 3133 418 3169
rect 336 3099 360 3133
rect 394 3099 418 3133
rect 336 3063 418 3099
rect 336 3029 360 3063
rect 394 3029 418 3063
rect 336 2993 418 3029
rect 336 2959 360 2993
rect 394 2959 418 2993
rect 336 2923 418 2959
rect 336 2889 360 2923
rect 394 2889 418 2923
rect 336 2853 418 2889
rect 336 2819 360 2853
rect 394 2819 418 2853
rect 336 2783 418 2819
rect 336 2749 360 2783
rect 394 2749 418 2783
rect 336 2713 418 2749
rect 336 2679 360 2713
rect 394 2679 418 2713
rect 336 2643 418 2679
rect 336 2609 360 2643
rect 394 2609 418 2643
rect 336 2573 418 2609
rect 336 2539 360 2573
rect 394 2539 418 2573
rect 336 2503 418 2539
rect 336 2469 360 2503
rect 394 2469 418 2503
rect 336 2433 418 2469
rect 336 2399 360 2433
rect 394 2399 418 2433
rect 336 2363 418 2399
rect 336 2329 360 2363
rect 394 2329 418 2363
rect 336 2293 418 2329
rect 10888 3699 10970 3735
rect 10888 3665 10912 3699
rect 10946 3665 10970 3699
rect 10888 3629 10970 3665
rect 10888 3595 10912 3629
rect 10946 3595 10970 3629
rect 10888 3559 10970 3595
rect 10888 3525 10912 3559
rect 10946 3525 10970 3559
rect 10888 3489 10970 3525
rect 10888 3455 10912 3489
rect 10946 3455 10970 3489
rect 10888 3419 10970 3455
rect 10888 3385 10912 3419
rect 10946 3385 10970 3419
rect 10888 3349 10970 3385
rect 10888 3315 10912 3349
rect 10946 3315 10970 3349
rect 10888 3279 10970 3315
rect 10888 3245 10912 3279
rect 10946 3245 10970 3279
rect 10888 3209 10970 3245
rect 10888 3175 10912 3209
rect 10946 3175 10970 3209
rect 10888 3139 10970 3175
rect 10888 3105 10912 3139
rect 10946 3105 10970 3139
rect 10888 3069 10970 3105
rect 10888 3035 10912 3069
rect 10946 3035 10970 3069
rect 10888 2999 10970 3035
rect 10888 2965 10912 2999
rect 10946 2965 10970 2999
rect 10888 2929 10970 2965
rect 10888 2895 10912 2929
rect 10946 2895 10970 2929
rect 10888 2859 10970 2895
rect 10888 2825 10912 2859
rect 10946 2825 10970 2859
rect 10888 2789 10970 2825
rect 10888 2755 10912 2789
rect 10946 2755 10970 2789
rect 10888 2719 10970 2755
rect 10888 2685 10912 2719
rect 10946 2685 10970 2719
rect 10888 2649 10970 2685
rect 10888 2615 10912 2649
rect 10946 2615 10970 2649
rect 10888 2578 10970 2615
rect 10888 2544 10912 2578
rect 10946 2544 10970 2578
rect 10888 2507 10970 2544
rect 10888 2473 10912 2507
rect 10946 2473 10970 2507
rect 10888 2436 10970 2473
rect 10888 2402 10912 2436
rect 10946 2402 10970 2436
rect 10888 2365 10970 2402
rect 10888 2331 10912 2365
rect 10946 2331 10970 2365
rect 336 2259 360 2293
rect 394 2259 418 2293
rect 336 2247 418 2259
rect 10888 2294 10970 2331
rect 10888 2260 10912 2294
rect 10946 2260 10970 2294
rect 10888 2247 10970 2260
rect 336 2223 10970 2247
rect 336 2189 360 2223
rect 394 2189 429 2223
rect 463 2189 498 2223
rect 532 2189 567 2223
rect 601 2189 636 2223
rect 670 2189 705 2223
rect 739 2189 774 2223
rect 808 2189 843 2223
rect 877 2189 912 2223
rect 946 2189 981 2223
rect 1015 2189 1050 2223
rect 1084 2189 1119 2223
rect 1153 2189 1188 2223
rect 1222 2189 1256 2223
rect 1290 2189 1324 2223
rect 1358 2189 1392 2223
rect 1426 2189 1460 2223
rect 1494 2189 1528 2223
rect 1562 2189 1596 2223
rect 1630 2189 1664 2223
rect 1698 2189 1732 2223
rect 1766 2189 1800 2223
rect 1834 2189 1868 2223
rect 1902 2189 1936 2223
rect 1970 2189 2004 2223
rect 2038 2189 2072 2223
rect 2106 2189 2140 2223
rect 2174 2189 2208 2223
rect 2242 2189 2276 2223
rect 2310 2189 2344 2223
rect 2378 2189 2412 2223
rect 2446 2189 2480 2223
rect 2514 2189 2548 2223
rect 2582 2189 2616 2223
rect 2650 2189 2684 2223
rect 2718 2189 2752 2223
rect 2786 2189 2820 2223
rect 2854 2189 2888 2223
rect 2922 2189 2956 2223
rect 2990 2189 3024 2223
rect 3058 2189 3092 2223
rect 3126 2189 3160 2223
rect 3194 2189 3228 2223
rect 3262 2189 3296 2223
rect 3330 2189 3364 2223
rect 3398 2189 3432 2223
rect 3466 2189 3500 2223
rect 3534 2189 3568 2223
rect 3602 2189 3636 2223
rect 3670 2189 3704 2223
rect 3738 2189 3772 2223
rect 3806 2189 3840 2223
rect 3874 2189 3908 2223
rect 3942 2189 3976 2223
rect 4010 2189 4044 2223
rect 4078 2189 4112 2223
rect 4146 2189 4180 2223
rect 4214 2189 4248 2223
rect 4282 2189 4316 2223
rect 4350 2189 4384 2223
rect 4418 2189 4452 2223
rect 4486 2189 4520 2223
rect 4554 2189 4588 2223
rect 4622 2189 4656 2223
rect 4690 2189 4724 2223
rect 4758 2189 4792 2223
rect 4826 2189 4860 2223
rect 4894 2189 4928 2223
rect 4962 2189 4996 2223
rect 5030 2189 5064 2223
rect 5098 2189 5132 2223
rect 5166 2189 5200 2223
rect 5234 2189 5268 2223
rect 5302 2189 5336 2223
rect 5370 2189 5404 2223
rect 5438 2189 5472 2223
rect 5506 2189 5540 2223
rect 5574 2189 5608 2223
rect 5642 2189 5676 2223
rect 5710 2189 5744 2223
rect 5778 2189 5812 2223
rect 5846 2189 5880 2223
rect 5914 2189 5948 2223
rect 5982 2189 6016 2223
rect 6050 2189 6084 2223
rect 6118 2189 6152 2223
rect 6186 2189 6220 2223
rect 6254 2189 6288 2223
rect 6322 2189 6356 2223
rect 6390 2189 6424 2223
rect 6458 2189 6492 2223
rect 6526 2189 6560 2223
rect 6594 2189 6628 2223
rect 6662 2189 6696 2223
rect 6730 2189 6764 2223
rect 6798 2189 6832 2223
rect 6866 2189 6900 2223
rect 6934 2189 6968 2223
rect 7002 2189 7036 2223
rect 7070 2189 7104 2223
rect 7138 2189 7172 2223
rect 7206 2189 7240 2223
rect 7274 2189 7308 2223
rect 7342 2189 7376 2223
rect 7410 2189 7444 2223
rect 7478 2189 7512 2223
rect 7546 2189 7580 2223
rect 7614 2189 7648 2223
rect 7682 2189 7716 2223
rect 7750 2189 7784 2223
rect 7818 2189 7852 2223
rect 7886 2189 7920 2223
rect 7954 2189 7988 2223
rect 8022 2189 8056 2223
rect 8090 2189 8124 2223
rect 8158 2189 8192 2223
rect 8226 2189 8260 2223
rect 8294 2189 8328 2223
rect 8362 2189 8396 2223
rect 8430 2189 8464 2223
rect 8498 2189 8532 2223
rect 8566 2189 8600 2223
rect 8634 2189 8668 2223
rect 8702 2189 8736 2223
rect 8770 2189 8804 2223
rect 8838 2189 8872 2223
rect 8906 2189 8940 2223
rect 8974 2189 9008 2223
rect 9042 2189 9076 2223
rect 9110 2189 9144 2223
rect 9178 2189 9212 2223
rect 9246 2189 9280 2223
rect 9314 2189 9348 2223
rect 9382 2189 9416 2223
rect 9450 2189 9484 2223
rect 9518 2189 9552 2223
rect 9586 2189 9620 2223
rect 9654 2189 9688 2223
rect 9722 2189 9756 2223
rect 9790 2189 9824 2223
rect 9858 2189 9892 2223
rect 9926 2189 9960 2223
rect 9994 2189 10028 2223
rect 10062 2189 10096 2223
rect 10130 2189 10164 2223
rect 10198 2189 10232 2223
rect 10266 2189 10300 2223
rect 10334 2189 10368 2223
rect 10402 2189 10436 2223
rect 10470 2189 10504 2223
rect 10538 2189 10572 2223
rect 10606 2189 10640 2223
rect 10674 2189 10708 2223
rect 10742 2189 10776 2223
rect 10810 2189 10844 2223
rect 10878 2189 10912 2223
rect 10946 2189 10970 2223
rect 336 2165 10970 2189
<< mvnsubdiff >>
rect 336 5799 10930 5823
rect 336 5765 360 5799
rect 394 5765 428 5799
rect 462 5765 496 5799
rect 530 5765 564 5799
rect 598 5765 632 5799
rect 666 5765 700 5799
rect 734 5765 768 5799
rect 802 5765 836 5799
rect 870 5765 904 5799
rect 938 5765 972 5799
rect 1006 5765 1040 5799
rect 1074 5765 1108 5799
rect 1142 5765 1176 5799
rect 1210 5765 1244 5799
rect 1278 5765 1312 5799
rect 1346 5765 1380 5799
rect 1414 5765 1448 5799
rect 1482 5765 1516 5799
rect 1550 5765 1584 5799
rect 1618 5765 1652 5799
rect 1686 5765 1720 5799
rect 1754 5765 1788 5799
rect 1822 5765 1856 5799
rect 1890 5765 1924 5799
rect 1958 5765 1992 5799
rect 2026 5765 2060 5799
rect 2094 5765 2128 5799
rect 2162 5765 2196 5799
rect 2230 5765 2264 5799
rect 2298 5765 2332 5799
rect 2366 5765 2400 5799
rect 2434 5765 2468 5799
rect 2502 5765 2536 5799
rect 2570 5765 2604 5799
rect 2638 5765 2672 5799
rect 2706 5765 2740 5799
rect 2774 5765 2808 5799
rect 2842 5765 2876 5799
rect 2910 5765 2944 5799
rect 2978 5765 3012 5799
rect 3046 5765 3080 5799
rect 3114 5765 3148 5799
rect 3182 5765 3216 5799
rect 3250 5765 3284 5799
rect 3318 5765 3352 5799
rect 3386 5765 3420 5799
rect 3454 5765 3488 5799
rect 3522 5765 3556 5799
rect 3590 5765 3624 5799
rect 3658 5765 3692 5799
rect 3726 5765 3760 5799
rect 3794 5765 3828 5799
rect 3862 5765 3896 5799
rect 3930 5765 3964 5799
rect 3998 5765 4032 5799
rect 4066 5765 4100 5799
rect 4134 5765 4168 5799
rect 4202 5765 4236 5799
rect 4270 5765 4304 5799
rect 4338 5765 4372 5799
rect 4406 5765 4440 5799
rect 4474 5765 4508 5799
rect 4542 5765 4576 5799
rect 4610 5765 4644 5799
rect 4678 5765 4712 5799
rect 4746 5765 4780 5799
rect 4814 5765 4848 5799
rect 4882 5765 4916 5799
rect 4950 5765 4984 5799
rect 5018 5765 5052 5799
rect 5086 5765 5120 5799
rect 5154 5765 5188 5799
rect 5222 5765 5256 5799
rect 5290 5765 5324 5799
rect 5358 5765 5392 5799
rect 5426 5765 5460 5799
rect 5494 5765 5528 5799
rect 5562 5765 5596 5799
rect 5630 5765 5664 5799
rect 5698 5765 5732 5799
rect 5766 5765 5800 5799
rect 5834 5765 5868 5799
rect 5902 5765 5936 5799
rect 5970 5765 6004 5799
rect 6038 5765 6072 5799
rect 6106 5765 6140 5799
rect 6174 5765 6208 5799
rect 6242 5765 6276 5799
rect 6310 5765 6344 5799
rect 6378 5765 6412 5799
rect 6446 5765 6480 5799
rect 6514 5765 6548 5799
rect 6582 5765 6616 5799
rect 6650 5765 6684 5799
rect 6718 5765 6752 5799
rect 6786 5765 6820 5799
rect 6854 5765 6888 5799
rect 6922 5765 6956 5799
rect 6990 5765 7024 5799
rect 7058 5765 7092 5799
rect 7126 5765 7160 5799
rect 7194 5765 7228 5799
rect 7262 5765 7296 5799
rect 7330 5765 7364 5799
rect 7398 5765 7432 5799
rect 7466 5765 7500 5799
rect 7534 5765 7568 5799
rect 7602 5765 7636 5799
rect 7670 5765 7704 5799
rect 7738 5765 7772 5799
rect 7806 5765 7840 5799
rect 7874 5765 7908 5799
rect 7942 5765 7976 5799
rect 8010 5765 8044 5799
rect 8078 5765 8112 5799
rect 8146 5765 8181 5799
rect 8215 5765 8250 5799
rect 8284 5765 8319 5799
rect 8353 5765 8388 5799
rect 8422 5765 8457 5799
rect 8491 5765 8526 5799
rect 8560 5765 8595 5799
rect 8629 5765 8664 5799
rect 8698 5765 8733 5799
rect 8767 5765 8802 5799
rect 8836 5765 8871 5799
rect 8905 5765 8940 5799
rect 8974 5765 9009 5799
rect 9043 5765 9078 5799
rect 9112 5765 9147 5799
rect 9181 5765 9216 5799
rect 9250 5765 9285 5799
rect 9319 5765 9354 5799
rect 9388 5765 9423 5799
rect 9457 5765 9492 5799
rect 9526 5765 9561 5799
rect 9595 5765 9630 5799
rect 9664 5765 9699 5799
rect 9733 5765 9768 5799
rect 9802 5765 9837 5799
rect 9871 5765 9906 5799
rect 9940 5765 9975 5799
rect 10009 5765 10044 5799
rect 10078 5765 10113 5799
rect 10147 5765 10182 5799
rect 10216 5765 10251 5799
rect 10285 5765 10320 5799
rect 10354 5765 10389 5799
rect 10423 5765 10458 5799
rect 10492 5765 10527 5799
rect 10561 5765 10596 5799
rect 10630 5765 10665 5799
rect 10699 5765 10734 5799
rect 10768 5765 10803 5799
rect 10837 5765 10872 5799
rect 10906 5765 10930 5799
rect 336 5741 10930 5765
rect 336 5724 418 5741
rect 336 5690 360 5724
rect 394 5690 418 5724
rect 10848 5730 10930 5741
rect 336 5649 418 5690
rect 10848 5696 10872 5730
rect 10906 5696 10930 5730
rect 336 5615 360 5649
rect 394 5615 418 5649
rect 336 5575 418 5615
rect 336 5541 360 5575
rect 394 5541 418 5575
rect 336 5501 418 5541
rect 336 5467 360 5501
rect 394 5467 418 5501
rect 336 5427 418 5467
rect 336 5393 360 5427
rect 394 5393 418 5427
rect 336 5321 418 5393
rect 336 5287 360 5321
rect 394 5287 418 5321
rect 336 5251 418 5287
rect 336 5217 360 5251
rect 394 5217 418 5251
rect 336 5181 418 5217
rect 336 5147 360 5181
rect 394 5147 418 5181
rect 336 5111 418 5147
rect 336 5077 360 5111
rect 394 5077 418 5111
rect 336 5041 418 5077
rect 336 5007 360 5041
rect 394 5007 418 5041
rect 336 4971 418 5007
rect 336 4937 360 4971
rect 394 4937 418 4971
rect 336 4902 418 4937
rect 336 4868 360 4902
rect 394 4868 418 4902
rect 336 4833 418 4868
rect 336 4799 360 4833
rect 394 4799 418 4833
rect 336 4764 418 4799
rect 336 4730 360 4764
rect 394 4730 418 4764
rect 336 4695 418 4730
rect 336 4661 360 4695
rect 394 4661 418 4695
rect 336 4626 418 4661
rect 336 4592 360 4626
rect 394 4592 418 4626
rect 336 4557 418 4592
rect 336 4523 360 4557
rect 394 4523 418 4557
rect 336 4488 418 4523
rect 336 4454 360 4488
rect 394 4454 418 4488
rect 336 4419 418 4454
rect 336 4385 360 4419
rect 394 4385 418 4419
rect 336 4350 418 4385
rect 336 4316 360 4350
rect 394 4316 418 4350
rect 336 4281 418 4316
rect 10848 5661 10930 5696
rect 10848 5627 10872 5661
rect 10906 5627 10930 5661
rect 10848 5592 10930 5627
rect 10848 5558 10872 5592
rect 10906 5558 10930 5592
rect 10848 5523 10930 5558
rect 10848 5489 10872 5523
rect 10906 5489 10930 5523
rect 10848 5454 10930 5489
rect 10848 5420 10872 5454
rect 10906 5420 10930 5454
rect 10848 5385 10930 5420
rect 10848 5351 10872 5385
rect 10906 5351 10930 5385
rect 10848 5316 10930 5351
rect 10848 5282 10872 5316
rect 10906 5282 10930 5316
rect 10848 5247 10930 5282
rect 10848 5213 10872 5247
rect 10906 5213 10930 5247
rect 10848 5178 10930 5213
rect 10848 5144 10872 5178
rect 10906 5144 10930 5178
rect 10848 5109 10930 5144
rect 10848 5075 10872 5109
rect 10906 5075 10930 5109
rect 10848 5040 10930 5075
rect 10848 5006 10872 5040
rect 10906 5006 10930 5040
rect 10848 4971 10930 5006
rect 10848 4937 10872 4971
rect 10906 4937 10930 4971
rect 10848 4902 10930 4937
rect 10848 4868 10872 4902
rect 10906 4868 10930 4902
rect 10848 4833 10930 4868
rect 10848 4799 10872 4833
rect 10906 4799 10930 4833
rect 10848 4764 10930 4799
rect 10848 4730 10872 4764
rect 10906 4730 10930 4764
rect 10848 4695 10930 4730
rect 10848 4661 10872 4695
rect 10906 4661 10930 4695
rect 10848 4626 10930 4661
rect 10848 4592 10872 4626
rect 10906 4592 10930 4626
rect 10848 4557 10930 4592
rect 10848 4523 10872 4557
rect 10906 4523 10930 4557
rect 10848 4488 10930 4523
rect 10848 4454 10872 4488
rect 10906 4454 10930 4488
rect 10848 4419 10930 4454
rect 10848 4385 10872 4419
rect 10906 4385 10930 4419
rect 10848 4350 10930 4385
rect 10848 4316 10872 4350
rect 10906 4316 10930 4350
rect 336 4247 360 4281
rect 394 4247 418 4281
rect 336 4212 418 4247
rect 336 4178 360 4212
rect 394 4178 418 4212
rect 10848 4281 10930 4316
rect 10848 4247 10872 4281
rect 10906 4247 10930 4281
rect 10848 4212 10930 4247
rect 336 4167 418 4178
rect 10848 4178 10872 4212
rect 10906 4178 10930 4212
rect 10848 4167 10930 4178
rect 336 4143 10930 4167
rect 336 4109 360 4143
rect 394 4109 429 4143
rect 463 4109 498 4143
rect 532 4109 567 4143
rect 601 4109 636 4143
rect 670 4109 705 4143
rect 739 4109 774 4143
rect 808 4109 843 4143
rect 877 4109 912 4143
rect 946 4109 981 4143
rect 1015 4109 1050 4143
rect 1084 4109 1119 4143
rect 1153 4109 1188 4143
rect 1222 4109 1257 4143
rect 1291 4109 1326 4143
rect 1360 4109 1395 4143
rect 1429 4109 1464 4143
rect 1498 4109 1533 4143
rect 1567 4109 1602 4143
rect 1636 4109 1671 4143
rect 1705 4109 1740 4143
rect 1774 4109 1809 4143
rect 1843 4109 1878 4143
rect 1912 4109 1947 4143
rect 1981 4109 2016 4143
rect 2050 4109 2085 4143
rect 2119 4109 2154 4143
rect 2188 4109 2223 4143
rect 2257 4109 2292 4143
rect 2326 4109 2361 4143
rect 2395 4109 2430 4143
rect 2464 4109 2499 4143
rect 2533 4109 2568 4143
rect 2602 4109 2637 4143
rect 2671 4109 2706 4143
rect 2740 4109 2775 4143
rect 2809 4109 2844 4143
rect 2878 4109 2913 4143
rect 2947 4109 2982 4143
rect 3016 4109 3051 4143
rect 3085 4109 3120 4143
rect 3154 4109 3188 4143
rect 3222 4109 3256 4143
rect 3290 4109 3324 4143
rect 3358 4109 3392 4143
rect 3426 4109 3460 4143
rect 3494 4109 3528 4143
rect 3562 4109 3596 4143
rect 3630 4109 3664 4143
rect 3698 4109 3732 4143
rect 3766 4109 3800 4143
rect 3834 4109 3868 4143
rect 3902 4109 3936 4143
rect 3970 4109 4004 4143
rect 4038 4109 4072 4143
rect 4106 4109 4140 4143
rect 4174 4109 4208 4143
rect 4242 4109 4276 4143
rect 4310 4109 4344 4143
rect 4378 4109 4412 4143
rect 4446 4109 4480 4143
rect 4514 4109 4548 4143
rect 4582 4109 4616 4143
rect 4650 4109 4684 4143
rect 4718 4109 4752 4143
rect 4786 4109 4820 4143
rect 4854 4109 4888 4143
rect 4922 4109 4956 4143
rect 4990 4109 5024 4143
rect 5058 4109 5092 4143
rect 5126 4109 5160 4143
rect 5194 4109 5228 4143
rect 5262 4109 5296 4143
rect 5330 4109 5364 4143
rect 5398 4109 5432 4143
rect 5466 4109 5500 4143
rect 5534 4109 5568 4143
rect 5602 4109 5636 4143
rect 5670 4109 5704 4143
rect 5738 4109 5772 4143
rect 5806 4109 5840 4143
rect 5874 4109 5908 4143
rect 5942 4109 5976 4143
rect 6010 4109 6044 4143
rect 6078 4109 6112 4143
rect 6146 4109 6180 4143
rect 6214 4109 6248 4143
rect 6282 4109 6316 4143
rect 6350 4109 6384 4143
rect 6418 4109 6452 4143
rect 6486 4109 6520 4143
rect 6554 4109 6588 4143
rect 6622 4109 6656 4143
rect 6690 4109 6724 4143
rect 6758 4109 6792 4143
rect 6826 4109 6860 4143
rect 6894 4109 6928 4143
rect 6962 4109 6996 4143
rect 7030 4109 7064 4143
rect 7098 4109 7132 4143
rect 7166 4109 7200 4143
rect 7234 4109 7268 4143
rect 7302 4109 7336 4143
rect 7370 4109 7404 4143
rect 7438 4109 7472 4143
rect 7506 4109 7540 4143
rect 7574 4109 7608 4143
rect 7642 4109 7676 4143
rect 7710 4109 7744 4143
rect 7778 4109 7812 4143
rect 7846 4109 7880 4143
rect 7914 4109 7948 4143
rect 7982 4109 8016 4143
rect 8050 4109 8084 4143
rect 8118 4109 8152 4143
rect 8186 4109 8220 4143
rect 8254 4109 8288 4143
rect 8322 4109 8356 4143
rect 8390 4109 8424 4143
rect 8458 4109 8492 4143
rect 8526 4109 8560 4143
rect 8594 4109 8628 4143
rect 8662 4109 8696 4143
rect 8730 4109 8764 4143
rect 8798 4109 8832 4143
rect 8866 4109 8900 4143
rect 8934 4109 8968 4143
rect 9002 4109 9036 4143
rect 9070 4109 9104 4143
rect 9138 4109 9172 4143
rect 9206 4109 9240 4143
rect 9274 4109 9308 4143
rect 9342 4109 9376 4143
rect 9410 4109 9444 4143
rect 9478 4109 9512 4143
rect 9546 4109 9580 4143
rect 9614 4109 9648 4143
rect 9682 4109 9716 4143
rect 9750 4109 9784 4143
rect 9818 4109 9852 4143
rect 9886 4109 9920 4143
rect 9954 4109 9988 4143
rect 10022 4109 10056 4143
rect 10090 4109 10124 4143
rect 10158 4109 10192 4143
rect 10226 4109 10260 4143
rect 10294 4109 10328 4143
rect 10362 4109 10396 4143
rect 10430 4109 10464 4143
rect 10498 4109 10532 4143
rect 10566 4109 10600 4143
rect 10634 4109 10668 4143
rect 10702 4109 10736 4143
rect 10770 4109 10804 4143
rect 10838 4109 10872 4143
rect 10906 4109 10930 4143
rect 336 4085 10930 4109
<< psubdiffcont >>
rect 336 7984 370 8018
rect 405 7984 439 8018
rect 474 7984 508 8018
rect 543 7984 577 8018
rect 612 7984 646 8018
rect 681 7984 715 8018
rect 750 7984 784 8018
rect 819 7984 853 8018
rect 888 7984 922 8018
rect 957 7984 991 8018
rect 1026 7984 1060 8018
rect 1095 7984 1129 8018
rect 1164 7984 1198 8018
rect 1233 7984 1267 8018
rect 1302 7984 1336 8018
rect 1371 7984 1405 8018
rect 1440 7984 1474 8018
rect 1509 7984 1543 8018
rect 1578 7984 1612 8018
rect 1647 7984 1681 8018
rect 1716 7984 1750 8018
rect 1784 7984 1818 8018
rect 1852 7984 1886 8018
rect 1920 7984 1954 8018
rect 1988 7984 2022 8018
rect 2056 7984 2090 8018
rect 2124 7984 2158 8018
rect 2192 7984 2226 8018
rect 2260 7984 2294 8018
rect 2328 7984 2362 8018
rect 2396 7984 2430 8018
rect 2464 7984 2498 8018
rect 2532 7984 2566 8018
rect 2600 7984 2634 8018
rect 2668 7984 2702 8018
rect 2736 7984 2770 8018
rect 2804 7984 2838 8018
rect 2872 7984 2906 8018
rect 2940 7984 2974 8018
rect 3008 7984 3042 8018
rect 3076 7984 3110 8018
rect 3144 7984 3178 8018
rect 3212 7984 3246 8018
rect 3280 7984 3314 8018
rect 3348 7984 3382 8018
rect 3416 7984 3450 8018
rect 3484 7984 3518 8018
rect 3552 7984 3586 8018
rect 3620 7984 3654 8018
rect 3688 7984 3722 8018
rect 3756 7984 3790 8018
rect 3824 7984 3858 8018
rect 3892 7984 3926 8018
rect 3960 7984 3994 8018
rect 4028 7984 4062 8018
rect 4096 7984 4130 8018
rect 4164 7984 4198 8018
rect 4232 7984 4266 8018
rect 4300 7984 4334 8018
rect 4368 7984 4402 8018
rect 4436 7984 4470 8018
rect 4504 7984 4538 8018
rect 4572 7984 4606 8018
rect 4640 7984 4674 8018
rect 4708 7984 4742 8018
rect 4776 7984 4810 8018
rect 4844 7984 4878 8018
rect 4912 7984 4946 8018
rect 4980 7984 5014 8018
rect 5048 7984 5082 8018
rect 5116 7984 5150 8018
rect 5184 7984 5218 8018
rect 5252 7984 5286 8018
rect 5320 7984 5354 8018
rect 5388 7984 5422 8018
rect 5456 7984 5490 8018
rect 5524 7984 5558 8018
rect 5592 7984 5626 8018
rect 5660 7984 5694 8018
rect 5728 7984 5762 8018
rect 5796 7984 5830 8018
rect 5864 7984 5898 8018
rect 5932 7984 5966 8018
rect 6000 7984 6034 8018
rect 6068 7984 6102 8018
rect 6136 7984 6170 8018
rect 6204 7984 6238 8018
rect 6272 7984 6306 8018
rect 6340 7984 6374 8018
rect 6408 7984 6442 8018
rect 6476 7984 6510 8018
rect 6544 7984 6578 8018
rect 6612 7984 6646 8018
rect 6680 7984 6714 8018
rect 6748 7984 6782 8018
rect 6816 7984 6850 8018
rect 6884 7984 6918 8018
rect 6952 7984 6986 8018
rect 7020 7984 7054 8018
rect 7088 7984 7122 8018
rect 7156 7984 7190 8018
rect 7224 7984 7258 8018
rect 7292 7984 7326 8018
rect 7360 7984 7394 8018
rect 7428 7984 7462 8018
rect 7496 7984 7530 8018
rect 7564 7984 7598 8018
rect 7632 7984 7666 8018
rect 7700 7984 7734 8018
rect 7768 7984 7802 8018
rect 7836 7984 7870 8018
rect 7904 7984 7938 8018
rect 7972 7984 8006 8018
rect 8040 7984 8074 8018
rect 8108 7984 8142 8018
rect 8176 7984 8210 8018
rect 8244 7984 8278 8018
rect 8312 7984 8346 8018
rect 8380 7984 8414 8018
rect 8448 7984 8482 8018
rect 8516 7984 8550 8018
rect 8584 7984 8618 8018
rect 8652 7984 8686 8018
rect 8720 7984 8754 8018
rect 8788 7984 8822 8018
rect 8856 7984 8890 8018
rect 8924 7984 8958 8018
rect 8992 7984 9026 8018
rect 9060 7984 9094 8018
rect 9128 7984 9162 8018
rect 9196 7984 9230 8018
rect 9264 7984 9298 8018
rect 9332 7984 9366 8018
rect 9400 7984 9434 8018
rect 9468 7984 9502 8018
rect 9536 7984 9570 8018
rect 9604 7984 9638 8018
rect 9672 7984 9706 8018
rect 9740 7984 9774 8018
rect 9808 7984 9842 8018
rect 9876 7984 9910 8018
rect 9944 7984 9978 8018
rect 10012 7984 10046 8018
rect 10080 7984 10114 8018
rect 10148 7984 10182 8018
rect 10216 7984 10250 8018
rect 10284 7984 10318 8018
rect 10352 7984 10386 8018
rect 10420 7984 10454 8018
rect 10488 7984 10522 8018
rect 10556 7984 10590 8018
rect 10624 7984 10658 8018
rect 10692 7984 10726 8018
rect 10760 7984 10794 8018
rect 10828 7984 10862 8018
rect 10896 7984 10930 8018
rect 10964 7984 10998 8018
rect 11032 7984 11066 8018
rect 11100 7984 11134 8018
rect 11168 7984 11202 8018
rect 11236 7984 11270 8018
rect 11304 7984 11338 8018
rect 11372 7984 11406 8018
rect 11440 7984 11474 8018
rect 11508 7984 11542 8018
rect 11576 7984 11610 8018
rect 11644 7984 11678 8018
rect 11712 7984 11746 8018
rect 11780 7984 11814 8018
rect 11848 7984 11882 8018
rect 11916 7984 11950 8018
rect 11984 7984 12018 8018
rect 12052 7984 12086 8018
rect 12120 7984 12154 8018
rect 12188 7984 12222 8018
rect 12256 7984 12290 8018
rect 12324 7984 12358 8018
rect 12392 7984 12426 8018
rect 12460 7984 12494 8018
rect 12528 7984 12562 8018
rect 12596 7984 12630 8018
rect 12664 7984 12698 8018
rect 12732 7984 12766 8018
rect 12800 7984 12834 8018
rect 12868 7984 12902 8018
rect 12936 7984 12970 8018
rect 13004 7984 13038 8018
rect 13072 7984 13106 8018
rect 13140 7984 13174 8018
rect 13208 7984 13242 8018
rect 13276 7984 13310 8018
rect 13344 7984 13378 8018
rect 13412 7984 13446 8018
rect 13480 7984 13514 8018
rect 13548 7984 13582 8018
rect 13616 7984 13650 8018
rect 13684 7984 13718 8018
rect 13752 7984 13786 8018
rect 13820 7984 13854 8018
rect 13888 7984 13922 8018
rect 13956 7984 13990 8018
rect 14024 7984 14058 8018
rect 14092 7984 14126 8018
rect 14160 7984 14194 8018
rect 14228 7984 14262 8018
rect 14296 7984 14330 8018
rect 14364 7984 14398 8018
rect 14432 7984 14466 8018
rect 14500 7984 14534 8018
rect 14568 7984 14602 8018
rect 14636 7984 14670 8018
rect 14774 7984 14808 8018
rect 14844 7984 14878 8018
rect 14914 7984 14948 8018
rect 14984 7984 15018 8018
rect 15054 7984 15088 8018
rect 15124 7984 15158 8018
rect 15194 7984 15228 8018
rect 15264 7984 15298 8018
rect 15334 7984 15368 8018
rect 15404 7984 15438 8018
rect 15474 7984 15508 8018
rect 15544 7984 15578 8018
rect 15614 7984 15648 8018
rect 15684 7984 15718 8018
rect 15754 7984 15788 8018
rect 15824 7984 15858 8018
rect 15894 7984 15928 8018
rect 15964 7984 15998 8018
rect 360 7874 394 7908
rect 360 7804 394 7838
rect 13194 7894 13228 7928
rect 13264 7894 13298 7928
rect 13334 7894 13368 7928
rect 13404 7894 13438 7928
rect 13474 7894 13508 7928
rect 13544 7894 13578 7928
rect 13614 7894 13648 7928
rect 13684 7894 13718 7928
rect 13754 7894 13788 7928
rect 13824 7894 13858 7928
rect 13894 7894 13928 7928
rect 13964 7894 13998 7928
rect 14034 7894 14068 7928
rect 14104 7894 14138 7928
rect 14174 7894 14208 7928
rect 14244 7894 14278 7928
rect 14314 7894 14348 7928
rect 14384 7894 14418 7928
rect 14454 7894 14488 7928
rect 14524 7894 14558 7928
rect 14594 7894 14628 7928
rect 14664 7894 14698 7928
rect 14774 7915 14808 7949
rect 14844 7915 14878 7949
rect 14914 7915 14948 7949
rect 14984 7915 15018 7949
rect 15054 7915 15088 7949
rect 15124 7915 15158 7949
rect 15194 7915 15228 7949
rect 15264 7915 15298 7949
rect 15334 7915 15368 7949
rect 15404 7915 15438 7949
rect 15474 7915 15508 7949
rect 15544 7915 15578 7949
rect 15614 7915 15648 7949
rect 15684 7915 15718 7949
rect 15754 7915 15788 7949
rect 15824 7915 15858 7949
rect 15894 7915 15928 7949
rect 15964 7915 15998 7949
rect 13194 7824 13228 7858
rect 13264 7824 13298 7858
rect 13334 7824 13368 7858
rect 13404 7824 13438 7858
rect 13474 7824 13508 7858
rect 13544 7824 13578 7858
rect 13614 7824 13648 7858
rect 13684 7824 13718 7858
rect 13754 7824 13788 7858
rect 13824 7824 13858 7858
rect 13894 7824 13928 7858
rect 13964 7824 13998 7858
rect 14034 7824 14068 7858
rect 14104 7824 14138 7858
rect 14174 7824 14208 7858
rect 14244 7824 14278 7858
rect 14314 7824 14348 7858
rect 14384 7824 14418 7858
rect 14454 7824 14488 7858
rect 14524 7824 14558 7858
rect 14594 7824 14628 7858
rect 14664 7824 14698 7858
rect 14774 7846 14808 7880
rect 14844 7846 14878 7880
rect 14914 7846 14948 7880
rect 14984 7846 15018 7880
rect 15054 7846 15088 7880
rect 15124 7846 15158 7880
rect 15194 7846 15228 7880
rect 15264 7846 15298 7880
rect 15334 7846 15368 7880
rect 15404 7846 15438 7880
rect 15474 7846 15508 7880
rect 15544 7846 15578 7880
rect 15614 7846 15648 7880
rect 15684 7846 15718 7880
rect 15754 7846 15788 7880
rect 15824 7846 15858 7880
rect 15894 7846 15928 7880
rect 15964 7846 15998 7880
rect 360 7734 394 7768
rect 13194 7754 13228 7788
rect 13264 7754 13298 7788
rect 13334 7754 13368 7788
rect 13404 7754 13438 7788
rect 13474 7754 13508 7788
rect 13544 7754 13578 7788
rect 13614 7754 13648 7788
rect 13684 7754 13718 7788
rect 13754 7754 13788 7788
rect 13824 7754 13858 7788
rect 13894 7754 13928 7788
rect 13964 7754 13998 7788
rect 14034 7754 14068 7788
rect 14104 7754 14138 7788
rect 14174 7754 14208 7788
rect 14244 7754 14278 7788
rect 14314 7754 14348 7788
rect 14384 7754 14418 7788
rect 14454 7754 14488 7788
rect 14524 7754 14558 7788
rect 14594 7754 14628 7788
rect 14664 7754 14698 7788
rect 14774 7777 14808 7811
rect 14844 7777 14878 7811
rect 14914 7777 14948 7811
rect 14984 7777 15018 7811
rect 15054 7777 15088 7811
rect 15124 7777 15158 7811
rect 15194 7777 15228 7811
rect 15264 7777 15298 7811
rect 15334 7777 15368 7811
rect 15404 7777 15438 7811
rect 15474 7777 15508 7811
rect 15544 7777 15578 7811
rect 15614 7777 15648 7811
rect 15684 7777 15718 7811
rect 15754 7777 15788 7811
rect 15824 7777 15858 7811
rect 15894 7777 15928 7811
rect 15964 7777 15998 7811
rect 360 7664 394 7698
rect 13194 7684 13228 7718
rect 13264 7684 13298 7718
rect 13334 7684 13368 7718
rect 13404 7684 13438 7718
rect 13474 7684 13508 7718
rect 13544 7684 13578 7718
rect 13614 7684 13648 7718
rect 13684 7684 13718 7718
rect 13754 7684 13788 7718
rect 13824 7684 13858 7718
rect 13894 7684 13928 7718
rect 13964 7684 13998 7718
rect 14034 7684 14068 7718
rect 14104 7684 14138 7718
rect 14174 7684 14208 7718
rect 14244 7684 14278 7718
rect 14314 7684 14348 7718
rect 14384 7684 14418 7718
rect 14454 7684 14488 7718
rect 14524 7684 14558 7718
rect 14594 7684 14628 7718
rect 14664 7684 14698 7718
rect 14774 7708 14808 7742
rect 14844 7708 14878 7742
rect 14914 7708 14948 7742
rect 14984 7708 15018 7742
rect 15054 7708 15088 7742
rect 15124 7708 15158 7742
rect 15194 7708 15228 7742
rect 15264 7708 15298 7742
rect 15334 7708 15368 7742
rect 15404 7708 15438 7742
rect 15474 7708 15508 7742
rect 15544 7708 15578 7742
rect 15614 7708 15648 7742
rect 15684 7708 15718 7742
rect 15754 7708 15788 7742
rect 15824 7708 15858 7742
rect 15894 7708 15928 7742
rect 15964 7708 15998 7742
rect 360 7594 394 7628
rect 13194 7614 13228 7648
rect 13264 7614 13298 7648
rect 13334 7614 13368 7648
rect 13404 7614 13438 7648
rect 13474 7614 13508 7648
rect 13544 7614 13578 7648
rect 13614 7614 13648 7648
rect 13684 7614 13718 7648
rect 13754 7614 13788 7648
rect 13824 7614 13858 7648
rect 13894 7614 13928 7648
rect 13964 7614 13998 7648
rect 14034 7614 14068 7648
rect 14104 7614 14138 7648
rect 14174 7614 14208 7648
rect 14244 7614 14278 7648
rect 14314 7614 14348 7648
rect 14384 7614 14418 7648
rect 14454 7614 14488 7648
rect 14524 7614 14558 7648
rect 14594 7614 14628 7648
rect 14664 7614 14698 7648
rect 14774 7639 14808 7673
rect 14844 7639 14878 7673
rect 14914 7639 14948 7673
rect 14984 7639 15018 7673
rect 15054 7639 15088 7673
rect 15124 7639 15158 7673
rect 15194 7639 15228 7673
rect 15264 7639 15298 7673
rect 15334 7639 15368 7673
rect 15404 7639 15438 7673
rect 15474 7639 15508 7673
rect 15544 7639 15578 7673
rect 15614 7639 15648 7673
rect 15684 7639 15718 7673
rect 15754 7639 15788 7673
rect 15824 7639 15858 7673
rect 15894 7639 15928 7673
rect 15964 7639 15998 7673
rect 360 7524 394 7558
rect 13194 7544 13228 7578
rect 13264 7544 13298 7578
rect 13334 7544 13368 7578
rect 13404 7544 13438 7578
rect 13474 7544 13508 7578
rect 13544 7544 13578 7578
rect 13614 7544 13648 7578
rect 13684 7544 13718 7578
rect 13754 7544 13788 7578
rect 13824 7544 13858 7578
rect 13894 7544 13928 7578
rect 13964 7544 13998 7578
rect 14034 7544 14068 7578
rect 14104 7544 14138 7578
rect 14174 7544 14208 7578
rect 14244 7544 14278 7578
rect 14314 7544 14348 7578
rect 14384 7544 14418 7578
rect 14454 7544 14488 7578
rect 14524 7544 14558 7578
rect 14594 7544 14628 7578
rect 14664 7544 14698 7578
rect 14774 7570 14808 7604
rect 14844 7570 14878 7604
rect 14914 7570 14948 7604
rect 14984 7570 15018 7604
rect 15054 7570 15088 7604
rect 15124 7570 15158 7604
rect 15194 7570 15228 7604
rect 15264 7570 15298 7604
rect 15334 7570 15368 7604
rect 15404 7570 15438 7604
rect 15474 7570 15508 7604
rect 15544 7570 15578 7604
rect 15614 7570 15648 7604
rect 15684 7570 15718 7604
rect 15754 7570 15788 7604
rect 15824 7570 15858 7604
rect 15894 7570 15928 7604
rect 15964 7570 15998 7604
rect 360 7454 394 7488
rect 13194 7474 13228 7508
rect 13264 7474 13298 7508
rect 13334 7474 13368 7508
rect 13404 7474 13438 7508
rect 13474 7474 13508 7508
rect 13544 7474 13578 7508
rect 13614 7474 13648 7508
rect 13684 7474 13718 7508
rect 13754 7474 13788 7508
rect 13824 7474 13858 7508
rect 13894 7474 13928 7508
rect 13964 7474 13998 7508
rect 14034 7474 14068 7508
rect 14104 7474 14138 7508
rect 14174 7474 14208 7508
rect 14244 7474 14278 7508
rect 14314 7474 14348 7508
rect 14384 7474 14418 7508
rect 14454 7474 14488 7508
rect 14524 7474 14558 7508
rect 14594 7474 14628 7508
rect 14664 7474 14698 7508
rect 14774 7501 14808 7535
rect 14844 7501 14878 7535
rect 14914 7501 14948 7535
rect 14984 7501 15018 7535
rect 15054 7501 15088 7535
rect 15124 7501 15158 7535
rect 15194 7501 15228 7535
rect 15264 7501 15298 7535
rect 15334 7501 15368 7535
rect 15404 7501 15438 7535
rect 15474 7501 15508 7535
rect 15544 7501 15578 7535
rect 15614 7501 15648 7535
rect 15684 7501 15718 7535
rect 15754 7501 15788 7535
rect 15824 7501 15858 7535
rect 15894 7501 15928 7535
rect 15964 7501 15998 7535
rect 360 7384 394 7418
rect 360 7314 394 7348
rect 13194 7404 13228 7438
rect 13264 7404 13298 7438
rect 13334 7404 13368 7438
rect 13404 7404 13438 7438
rect 13474 7404 13508 7438
rect 13544 7404 13578 7438
rect 13614 7404 13648 7438
rect 13684 7404 13718 7438
rect 13754 7404 13788 7438
rect 13824 7404 13858 7438
rect 13894 7404 13928 7438
rect 13964 7404 13998 7438
rect 14034 7404 14068 7438
rect 14104 7404 14138 7438
rect 14174 7404 14208 7438
rect 14244 7404 14278 7438
rect 14314 7404 14348 7438
rect 14384 7404 14418 7438
rect 14454 7404 14488 7438
rect 14524 7404 14558 7438
rect 14594 7404 14628 7438
rect 14664 7404 14698 7438
rect 14774 7432 14808 7466
rect 14844 7432 14878 7466
rect 14914 7432 14948 7466
rect 14984 7432 15018 7466
rect 15054 7432 15088 7466
rect 15124 7432 15158 7466
rect 15194 7432 15228 7466
rect 15264 7432 15298 7466
rect 15334 7432 15368 7466
rect 15404 7432 15438 7466
rect 15474 7432 15508 7466
rect 15544 7432 15578 7466
rect 15614 7432 15648 7466
rect 15684 7432 15718 7466
rect 15754 7432 15788 7466
rect 15824 7432 15858 7466
rect 15894 7432 15928 7466
rect 15964 7432 15998 7466
rect 13194 7334 13228 7368
rect 13264 7334 13298 7368
rect 13334 7334 13368 7368
rect 13404 7334 13438 7368
rect 13474 7334 13508 7368
rect 13544 7334 13578 7368
rect 13614 7334 13648 7368
rect 13684 7334 13718 7368
rect 13754 7334 13788 7368
rect 13824 7334 13858 7368
rect 13894 7334 13928 7368
rect 13964 7334 13998 7368
rect 14034 7334 14068 7368
rect 14104 7334 14138 7368
rect 14174 7334 14208 7368
rect 14244 7334 14278 7368
rect 14314 7334 14348 7368
rect 14384 7334 14418 7368
rect 14454 7334 14488 7368
rect 14524 7334 14558 7368
rect 14594 7334 14628 7368
rect 14664 7334 14698 7368
rect 14774 7363 14808 7397
rect 14844 7363 14878 7397
rect 14914 7363 14948 7397
rect 14984 7363 15018 7397
rect 15054 7363 15088 7397
rect 15124 7363 15158 7397
rect 15194 7363 15228 7397
rect 15264 7363 15298 7397
rect 15334 7363 15368 7397
rect 15404 7363 15438 7397
rect 15474 7363 15508 7397
rect 15544 7363 15578 7397
rect 15614 7363 15648 7397
rect 15684 7363 15718 7397
rect 15754 7363 15788 7397
rect 15824 7363 15858 7397
rect 15894 7363 15928 7397
rect 15964 7363 15998 7397
rect 360 7244 394 7278
rect 360 7174 394 7208
rect 13194 7264 13228 7298
rect 13264 7264 13298 7298
rect 13334 7264 13368 7298
rect 13404 7264 13438 7298
rect 13474 7264 13508 7298
rect 13544 7264 13578 7298
rect 13614 7264 13648 7298
rect 13684 7264 13718 7298
rect 13754 7264 13788 7298
rect 13824 7264 13858 7298
rect 13894 7264 13928 7298
rect 13964 7264 13998 7298
rect 14034 7264 14068 7298
rect 14104 7264 14138 7298
rect 14174 7264 14208 7298
rect 14244 7264 14278 7298
rect 14314 7264 14348 7298
rect 14384 7264 14418 7298
rect 14454 7264 14488 7298
rect 14524 7264 14558 7298
rect 14594 7264 14628 7298
rect 14664 7264 14698 7298
rect 14774 7294 14808 7328
rect 14844 7294 14878 7328
rect 14914 7294 14948 7328
rect 14984 7294 15018 7328
rect 15054 7294 15088 7328
rect 15124 7294 15158 7328
rect 15194 7294 15228 7328
rect 15264 7294 15298 7328
rect 15334 7294 15368 7328
rect 15404 7294 15438 7328
rect 15474 7294 15508 7328
rect 15544 7294 15578 7328
rect 15614 7294 15648 7328
rect 15684 7294 15718 7328
rect 15754 7294 15788 7328
rect 15824 7294 15858 7328
rect 15894 7294 15928 7328
rect 15964 7294 15998 7328
rect 13194 7194 13228 7228
rect 13264 7194 13298 7228
rect 13334 7194 13368 7228
rect 13404 7194 13438 7228
rect 13474 7194 13508 7228
rect 13544 7194 13578 7228
rect 13614 7194 13648 7228
rect 13684 7194 13718 7228
rect 13754 7194 13788 7228
rect 13824 7194 13858 7228
rect 13894 7194 13928 7228
rect 13964 7194 13998 7228
rect 14034 7194 14068 7228
rect 14104 7194 14138 7228
rect 14174 7194 14208 7228
rect 14244 7194 14278 7228
rect 14314 7194 14348 7228
rect 14384 7194 14418 7228
rect 14454 7194 14488 7228
rect 14524 7194 14558 7228
rect 14594 7194 14628 7228
rect 14664 7194 14698 7228
rect 14774 7225 14808 7259
rect 14844 7225 14878 7259
rect 14914 7225 14948 7259
rect 14984 7225 15018 7259
rect 15054 7225 15088 7259
rect 15124 7225 15158 7259
rect 15194 7225 15228 7259
rect 15264 7225 15298 7259
rect 15334 7225 15368 7259
rect 15404 7225 15438 7259
rect 15474 7225 15508 7259
rect 15544 7225 15578 7259
rect 15614 7225 15648 7259
rect 15684 7225 15718 7259
rect 15754 7225 15788 7259
rect 15824 7225 15858 7259
rect 15894 7225 15928 7259
rect 15964 7225 15998 7259
rect 360 7104 394 7138
rect 360 7034 394 7068
rect 13194 7124 13228 7158
rect 13264 7124 13298 7158
rect 13334 7124 13368 7158
rect 13404 7124 13438 7158
rect 13474 7124 13508 7158
rect 13544 7124 13578 7158
rect 13614 7124 13648 7158
rect 13684 7124 13718 7158
rect 13754 7124 13788 7158
rect 13824 7124 13858 7158
rect 13894 7124 13928 7158
rect 13964 7124 13998 7158
rect 14034 7124 14068 7158
rect 14104 7124 14138 7158
rect 14174 7124 14208 7158
rect 14244 7124 14278 7158
rect 14314 7124 14348 7158
rect 14384 7124 14418 7158
rect 14454 7124 14488 7158
rect 14524 7124 14558 7158
rect 14594 7124 14628 7158
rect 14664 7124 14698 7158
rect 14774 7156 14808 7190
rect 14844 7156 14878 7190
rect 14914 7156 14948 7190
rect 14984 7156 15018 7190
rect 15054 7156 15088 7190
rect 15124 7156 15158 7190
rect 15194 7156 15228 7190
rect 15264 7156 15298 7190
rect 15334 7156 15368 7190
rect 15404 7156 15438 7190
rect 15474 7156 15508 7190
rect 15544 7156 15578 7190
rect 15614 7156 15648 7190
rect 15684 7156 15718 7190
rect 15754 7156 15788 7190
rect 15824 7156 15858 7190
rect 15894 7156 15928 7190
rect 15964 7156 15998 7190
rect 13194 7054 13228 7088
rect 13264 7054 13298 7088
rect 13334 7054 13368 7088
rect 13404 7054 13438 7088
rect 13474 7054 13508 7088
rect 13544 7054 13578 7088
rect 13614 7054 13648 7088
rect 13684 7054 13718 7088
rect 13754 7054 13788 7088
rect 13824 7054 13858 7088
rect 13894 7054 13928 7088
rect 13964 7054 13998 7088
rect 14034 7054 14068 7088
rect 14104 7054 14138 7088
rect 14174 7054 14208 7088
rect 14244 7054 14278 7088
rect 14314 7054 14348 7088
rect 14384 7054 14418 7088
rect 14454 7054 14488 7088
rect 14524 7054 14558 7088
rect 14594 7054 14628 7088
rect 14664 7054 14698 7088
rect 14774 7087 14808 7121
rect 14844 7087 14878 7121
rect 14914 7087 14948 7121
rect 14984 7087 15018 7121
rect 15054 7087 15088 7121
rect 15124 7087 15158 7121
rect 15194 7087 15228 7121
rect 15264 7087 15298 7121
rect 15334 7087 15368 7121
rect 15404 7087 15438 7121
rect 15474 7087 15508 7121
rect 15544 7087 15578 7121
rect 15614 7087 15648 7121
rect 15684 7087 15718 7121
rect 15754 7087 15788 7121
rect 15824 7087 15858 7121
rect 15894 7087 15928 7121
rect 15964 7087 15998 7121
rect 360 6965 394 6999
rect 14774 7018 14808 7052
rect 14844 7018 14878 7052
rect 14914 7018 14948 7052
rect 14984 7018 15018 7052
rect 15054 7018 15088 7052
rect 15124 7018 15158 7052
rect 15194 7018 15228 7052
rect 15264 7018 15298 7052
rect 15334 7018 15368 7052
rect 15404 7018 15438 7052
rect 15474 7018 15508 7052
rect 15544 7018 15578 7052
rect 15614 7018 15648 7052
rect 15684 7018 15718 7052
rect 15754 7018 15788 7052
rect 15824 7018 15858 7052
rect 15894 7018 15928 7052
rect 15964 7018 15998 7052
rect 13194 6984 13228 7018
rect 13264 6984 13298 7018
rect 13334 6984 13368 7018
rect 13404 6984 13438 7018
rect 13474 6984 13508 7018
rect 13544 6984 13578 7018
rect 13614 6984 13648 7018
rect 13684 6984 13718 7018
rect 13754 6984 13788 7018
rect 13824 6984 13858 7018
rect 13894 6984 13928 7018
rect 13964 6984 13998 7018
rect 14034 6984 14068 7018
rect 14104 6984 14138 7018
rect 14174 6984 14208 7018
rect 14244 6984 14278 7018
rect 14314 6984 14348 7018
rect 14384 6984 14418 7018
rect 14454 6984 14488 7018
rect 14524 6984 14558 7018
rect 14594 6984 14628 7018
rect 14664 6984 14698 7018
rect 360 6896 394 6930
rect 14774 6949 14808 6983
rect 14844 6949 14878 6983
rect 14914 6949 14948 6983
rect 14984 6949 15018 6983
rect 15054 6949 15088 6983
rect 15124 6949 15158 6983
rect 15194 6949 15228 6983
rect 15264 6949 15298 6983
rect 15334 6949 15368 6983
rect 15404 6949 15438 6983
rect 15474 6949 15508 6983
rect 15544 6949 15578 6983
rect 15614 6949 15648 6983
rect 15684 6949 15718 6983
rect 15754 6949 15788 6983
rect 15824 6949 15858 6983
rect 15894 6949 15928 6983
rect 15964 6949 15998 6983
rect 13194 6914 13228 6948
rect 13264 6914 13298 6948
rect 13334 6914 13368 6948
rect 13404 6914 13438 6948
rect 13474 6914 13508 6948
rect 13544 6914 13578 6948
rect 13614 6914 13648 6948
rect 13684 6914 13718 6948
rect 13754 6914 13788 6948
rect 13824 6914 13858 6948
rect 13894 6914 13928 6948
rect 13964 6914 13998 6948
rect 14034 6914 14068 6948
rect 14104 6914 14138 6948
rect 14174 6914 14208 6948
rect 14244 6914 14278 6948
rect 14314 6914 14348 6948
rect 14384 6914 14418 6948
rect 14454 6914 14488 6948
rect 14524 6914 14558 6948
rect 14594 6914 14628 6948
rect 14664 6914 14698 6948
rect 360 6827 394 6861
rect 14774 6880 14808 6914
rect 14844 6880 14878 6914
rect 14914 6880 14948 6914
rect 14984 6880 15018 6914
rect 15054 6880 15088 6914
rect 15124 6880 15158 6914
rect 15194 6880 15228 6914
rect 15264 6880 15298 6914
rect 15334 6880 15368 6914
rect 15404 6880 15438 6914
rect 15474 6880 15508 6914
rect 15544 6880 15578 6914
rect 15614 6880 15648 6914
rect 15684 6880 15718 6914
rect 15754 6880 15788 6914
rect 15824 6880 15858 6914
rect 15894 6880 15928 6914
rect 15964 6880 15998 6914
rect 13194 6844 13228 6878
rect 13264 6844 13298 6878
rect 13334 6844 13368 6878
rect 13404 6844 13438 6878
rect 13474 6844 13508 6878
rect 13544 6844 13578 6878
rect 13614 6844 13648 6878
rect 13684 6844 13718 6878
rect 13754 6844 13788 6878
rect 13824 6844 13858 6878
rect 13894 6844 13928 6878
rect 13964 6844 13998 6878
rect 14034 6844 14068 6878
rect 14104 6844 14138 6878
rect 14174 6844 14208 6878
rect 14244 6844 14278 6878
rect 14314 6844 14348 6878
rect 14384 6844 14418 6878
rect 14454 6844 14488 6878
rect 14524 6844 14558 6878
rect 14594 6844 14628 6878
rect 14664 6844 14698 6878
rect 360 6758 394 6792
rect 14774 6811 14808 6845
rect 14844 6811 14878 6845
rect 14914 6811 14948 6845
rect 14984 6811 15018 6845
rect 15054 6811 15088 6845
rect 15124 6811 15158 6845
rect 15194 6811 15228 6845
rect 15264 6811 15298 6845
rect 15334 6811 15368 6845
rect 15404 6811 15438 6845
rect 15474 6811 15508 6845
rect 15544 6811 15578 6845
rect 15614 6811 15648 6845
rect 15684 6811 15718 6845
rect 15754 6811 15788 6845
rect 15824 6811 15858 6845
rect 15894 6811 15928 6845
rect 15964 6811 15998 6845
rect 13194 6774 13228 6808
rect 13264 6774 13298 6808
rect 13334 6774 13368 6808
rect 13404 6774 13438 6808
rect 13474 6774 13508 6808
rect 13544 6774 13578 6808
rect 13614 6774 13648 6808
rect 13684 6774 13718 6808
rect 13754 6774 13788 6808
rect 13824 6774 13858 6808
rect 13894 6774 13928 6808
rect 13964 6774 13998 6808
rect 14034 6774 14068 6808
rect 14104 6774 14138 6808
rect 14174 6774 14208 6808
rect 14244 6774 14278 6808
rect 14314 6774 14348 6808
rect 14384 6774 14418 6808
rect 14454 6774 14488 6808
rect 14524 6774 14558 6808
rect 14594 6774 14628 6808
rect 14664 6774 14698 6808
rect 14774 6742 14808 6776
rect 14844 6742 14878 6776
rect 14914 6742 14948 6776
rect 14984 6742 15018 6776
rect 15054 6742 15088 6776
rect 15124 6742 15158 6776
rect 15194 6742 15228 6776
rect 15264 6742 15298 6776
rect 15334 6742 15368 6776
rect 15404 6742 15438 6776
rect 15474 6742 15508 6776
rect 15544 6742 15578 6776
rect 15614 6742 15648 6776
rect 15684 6742 15718 6776
rect 15754 6742 15788 6776
rect 15824 6742 15858 6776
rect 15894 6742 15928 6776
rect 15964 6742 15998 6776
rect 360 6689 394 6723
rect 13194 6704 13228 6738
rect 13264 6704 13298 6738
rect 13334 6704 13368 6738
rect 13404 6704 13438 6738
rect 13474 6704 13508 6738
rect 13544 6704 13578 6738
rect 13614 6704 13648 6738
rect 13684 6704 13718 6738
rect 13754 6704 13788 6738
rect 13824 6704 13858 6738
rect 13894 6704 13928 6738
rect 13964 6704 13998 6738
rect 14034 6704 14068 6738
rect 14104 6704 14138 6738
rect 14174 6704 14208 6738
rect 14244 6704 14278 6738
rect 14314 6704 14348 6738
rect 14384 6704 14418 6738
rect 14454 6704 14488 6738
rect 14524 6704 14558 6738
rect 14594 6704 14628 6738
rect 14664 6704 14698 6738
rect 360 6620 394 6654
rect 360 6551 394 6585
rect 14774 6673 14808 6707
rect 14844 6673 14878 6707
rect 14914 6673 14948 6707
rect 14984 6673 15018 6707
rect 15054 6673 15088 6707
rect 15124 6673 15158 6707
rect 15194 6673 15228 6707
rect 15264 6673 15298 6707
rect 15334 6673 15368 6707
rect 15404 6673 15438 6707
rect 15474 6673 15508 6707
rect 15544 6673 15578 6707
rect 15614 6673 15648 6707
rect 15684 6673 15718 6707
rect 15754 6673 15788 6707
rect 15824 6673 15858 6707
rect 15894 6673 15928 6707
rect 15964 6673 15998 6707
rect 13194 6634 13228 6668
rect 13264 6634 13298 6668
rect 13334 6634 13368 6668
rect 13404 6634 13438 6668
rect 13474 6634 13508 6668
rect 13544 6634 13578 6668
rect 13614 6634 13648 6668
rect 13684 6634 13718 6668
rect 13754 6634 13788 6668
rect 13824 6634 13858 6668
rect 13894 6634 13928 6668
rect 13964 6634 13998 6668
rect 14034 6634 14068 6668
rect 14104 6634 14138 6668
rect 14174 6634 14208 6668
rect 14244 6634 14278 6668
rect 14314 6634 14348 6668
rect 14384 6634 14418 6668
rect 14454 6634 14488 6668
rect 14524 6634 14558 6668
rect 14594 6634 14628 6668
rect 14664 6634 14698 6668
rect 14774 6604 14808 6638
rect 14844 6604 14878 6638
rect 14914 6604 14948 6638
rect 14984 6604 15018 6638
rect 15054 6604 15088 6638
rect 15124 6604 15158 6638
rect 15194 6604 15228 6638
rect 15264 6604 15298 6638
rect 15334 6604 15368 6638
rect 15404 6604 15438 6638
rect 15474 6604 15508 6638
rect 15544 6604 15578 6638
rect 15614 6604 15648 6638
rect 15684 6604 15718 6638
rect 15754 6604 15788 6638
rect 15824 6604 15858 6638
rect 15894 6604 15928 6638
rect 15964 6604 15998 6638
rect 13194 6564 13228 6598
rect 13264 6564 13298 6598
rect 13334 6564 13368 6598
rect 13404 6564 13438 6598
rect 13474 6564 13508 6598
rect 13544 6564 13578 6598
rect 13614 6564 13648 6598
rect 13684 6564 13718 6598
rect 13754 6564 13788 6598
rect 13824 6564 13858 6598
rect 13894 6564 13928 6598
rect 13964 6564 13998 6598
rect 14034 6564 14068 6598
rect 14104 6564 14138 6598
rect 14174 6564 14208 6598
rect 14244 6564 14278 6598
rect 14314 6564 14348 6598
rect 14384 6564 14418 6598
rect 14454 6564 14488 6598
rect 14524 6564 14558 6598
rect 14594 6564 14628 6598
rect 14664 6564 14698 6598
rect 14774 6535 14808 6569
rect 14844 6535 14878 6569
rect 14914 6535 14948 6569
rect 14984 6535 15018 6569
rect 15054 6535 15088 6569
rect 15124 6535 15158 6569
rect 15194 6535 15228 6569
rect 15264 6535 15298 6569
rect 15334 6535 15368 6569
rect 15404 6535 15438 6569
rect 15474 6535 15508 6569
rect 15544 6535 15578 6569
rect 15614 6535 15648 6569
rect 15684 6535 15718 6569
rect 15754 6535 15788 6569
rect 15824 6535 15858 6569
rect 15894 6535 15928 6569
rect 15964 6535 15998 6569
rect 360 6482 394 6516
rect 360 6413 394 6447
rect 13194 6494 13228 6528
rect 13264 6494 13298 6528
rect 13334 6494 13368 6528
rect 13404 6494 13438 6528
rect 13474 6494 13508 6528
rect 13544 6494 13578 6528
rect 13614 6494 13648 6528
rect 13684 6494 13718 6528
rect 13754 6494 13788 6528
rect 13824 6494 13858 6528
rect 13894 6494 13928 6528
rect 13964 6494 13998 6528
rect 14034 6494 14068 6528
rect 14104 6494 14138 6528
rect 14174 6494 14208 6528
rect 14244 6494 14278 6528
rect 14314 6494 14348 6528
rect 14384 6494 14418 6528
rect 14454 6494 14488 6528
rect 14524 6494 14558 6528
rect 14594 6494 14628 6528
rect 14664 6494 14698 6528
rect 14774 6466 14808 6500
rect 14844 6466 14878 6500
rect 14914 6466 14948 6500
rect 14984 6466 15018 6500
rect 15054 6466 15088 6500
rect 15124 6466 15158 6500
rect 15194 6466 15228 6500
rect 15264 6466 15298 6500
rect 15334 6466 15368 6500
rect 15404 6466 15438 6500
rect 15474 6466 15508 6500
rect 15544 6466 15578 6500
rect 15614 6466 15648 6500
rect 15684 6466 15718 6500
rect 15754 6466 15788 6500
rect 15824 6466 15858 6500
rect 15894 6466 15928 6500
rect 15964 6466 15998 6500
rect 13194 6424 13228 6458
rect 13264 6424 13298 6458
rect 13334 6424 13368 6458
rect 13404 6424 13438 6458
rect 13474 6424 13508 6458
rect 13544 6424 13578 6458
rect 13614 6424 13648 6458
rect 13684 6424 13718 6458
rect 13754 6424 13788 6458
rect 13824 6424 13858 6458
rect 13894 6424 13928 6458
rect 13964 6424 13998 6458
rect 14034 6424 14068 6458
rect 14104 6424 14138 6458
rect 14174 6424 14208 6458
rect 14244 6424 14278 6458
rect 14314 6424 14348 6458
rect 14384 6424 14418 6458
rect 14454 6424 14488 6458
rect 14524 6424 14558 6458
rect 14594 6424 14628 6458
rect 14664 6424 14698 6458
rect 360 6344 394 6378
rect 14774 6397 14808 6431
rect 14844 6397 14878 6431
rect 14914 6397 14948 6431
rect 14984 6397 15018 6431
rect 15054 6397 15088 6431
rect 15124 6397 15158 6431
rect 15194 6397 15228 6431
rect 15264 6397 15298 6431
rect 15334 6397 15368 6431
rect 15404 6397 15438 6431
rect 15474 6397 15508 6431
rect 15544 6397 15578 6431
rect 15614 6397 15648 6431
rect 15684 6397 15718 6431
rect 15754 6397 15788 6431
rect 15824 6397 15858 6431
rect 15894 6397 15928 6431
rect 15964 6397 15998 6431
rect 360 6275 394 6309
rect 13194 6354 13228 6388
rect 13264 6354 13298 6388
rect 13334 6354 13368 6388
rect 13404 6354 13438 6388
rect 13474 6354 13508 6388
rect 13544 6354 13578 6388
rect 13614 6354 13648 6388
rect 13684 6354 13718 6388
rect 13754 6354 13788 6388
rect 13824 6354 13858 6388
rect 13894 6354 13928 6388
rect 13964 6354 13998 6388
rect 14034 6354 14068 6388
rect 14104 6354 14138 6388
rect 14174 6354 14208 6388
rect 14244 6354 14278 6388
rect 14314 6354 14348 6388
rect 14384 6354 14418 6388
rect 14454 6354 14488 6388
rect 14524 6354 14558 6388
rect 14594 6354 14628 6388
rect 14664 6354 14698 6388
rect 14774 6328 14808 6362
rect 14844 6328 14878 6362
rect 14914 6328 14948 6362
rect 14984 6328 15018 6362
rect 15054 6328 15088 6362
rect 15124 6328 15158 6362
rect 15194 6328 15228 6362
rect 15264 6328 15298 6362
rect 15334 6328 15368 6362
rect 15404 6328 15438 6362
rect 15474 6328 15508 6362
rect 15544 6328 15578 6362
rect 15614 6328 15648 6362
rect 15684 6328 15718 6362
rect 15754 6328 15788 6362
rect 15824 6328 15858 6362
rect 15894 6328 15928 6362
rect 15964 6328 15998 6362
rect 13194 6284 13228 6318
rect 13264 6284 13298 6318
rect 13334 6284 13368 6318
rect 13404 6284 13438 6318
rect 13474 6284 13508 6318
rect 13544 6284 13578 6318
rect 13614 6284 13648 6318
rect 13684 6284 13718 6318
rect 13754 6284 13788 6318
rect 13824 6284 13858 6318
rect 13894 6284 13928 6318
rect 13964 6284 13998 6318
rect 14034 6284 14068 6318
rect 14104 6284 14138 6318
rect 14174 6284 14208 6318
rect 14244 6284 14278 6318
rect 14314 6284 14348 6318
rect 14384 6284 14418 6318
rect 14454 6284 14488 6318
rect 14524 6284 14558 6318
rect 14594 6284 14628 6318
rect 14664 6284 14698 6318
rect 360 6206 394 6240
rect 14774 6259 14808 6293
rect 14844 6259 14878 6293
rect 14914 6259 14948 6293
rect 14984 6259 15018 6293
rect 15054 6259 15088 6293
rect 15124 6259 15158 6293
rect 15194 6259 15228 6293
rect 15264 6259 15298 6293
rect 15334 6259 15368 6293
rect 15404 6259 15438 6293
rect 15474 6259 15508 6293
rect 15544 6259 15578 6293
rect 15614 6259 15648 6293
rect 15684 6259 15718 6293
rect 15754 6259 15788 6293
rect 15824 6259 15858 6293
rect 15894 6259 15928 6293
rect 15964 6259 15998 6293
rect 13194 6214 13228 6248
rect 13264 6214 13298 6248
rect 13334 6214 13368 6248
rect 13404 6214 13438 6248
rect 13474 6214 13508 6248
rect 13544 6214 13578 6248
rect 13614 6214 13648 6248
rect 13684 6214 13718 6248
rect 13754 6214 13788 6248
rect 13824 6214 13858 6248
rect 13894 6214 13928 6248
rect 13964 6214 13998 6248
rect 14034 6214 14068 6248
rect 14104 6214 14138 6248
rect 14174 6214 14208 6248
rect 14244 6214 14278 6248
rect 14314 6214 14348 6248
rect 14384 6214 14418 6248
rect 14454 6214 14488 6248
rect 14524 6214 14558 6248
rect 14594 6214 14628 6248
rect 14664 6214 14698 6248
rect 360 6137 394 6171
rect 14774 6190 14808 6224
rect 14844 6190 14878 6224
rect 14914 6190 14948 6224
rect 14984 6190 15018 6224
rect 15054 6190 15088 6224
rect 15124 6190 15158 6224
rect 15194 6190 15228 6224
rect 15264 6190 15298 6224
rect 15334 6190 15368 6224
rect 15404 6190 15438 6224
rect 15474 6190 15508 6224
rect 15544 6190 15578 6224
rect 15614 6190 15648 6224
rect 15684 6190 15718 6224
rect 15754 6190 15788 6224
rect 15824 6190 15858 6224
rect 15894 6190 15928 6224
rect 15964 6190 15998 6224
rect 13194 6144 13228 6178
rect 13264 6144 13298 6178
rect 13334 6144 13368 6178
rect 13404 6144 13438 6178
rect 13474 6144 13508 6178
rect 13544 6144 13578 6178
rect 13614 6144 13648 6178
rect 13684 6144 13718 6178
rect 13754 6144 13788 6178
rect 13824 6144 13858 6178
rect 13894 6144 13928 6178
rect 13964 6144 13998 6178
rect 14034 6144 14068 6178
rect 14104 6144 14138 6178
rect 14174 6144 14208 6178
rect 14244 6144 14278 6178
rect 14314 6144 14348 6178
rect 14384 6144 14418 6178
rect 14454 6144 14488 6178
rect 14524 6144 14558 6178
rect 14594 6144 14628 6178
rect 14664 6144 14698 6178
rect 14774 6121 14808 6155
rect 14844 6121 14878 6155
rect 14914 6121 14948 6155
rect 14984 6121 15018 6155
rect 15054 6121 15088 6155
rect 15124 6121 15158 6155
rect 15194 6121 15228 6155
rect 15264 6121 15298 6155
rect 15334 6121 15368 6155
rect 15404 6121 15438 6155
rect 15474 6121 15508 6155
rect 15544 6121 15578 6155
rect 15614 6121 15648 6155
rect 15684 6121 15718 6155
rect 15754 6121 15788 6155
rect 15824 6121 15858 6155
rect 15894 6121 15928 6155
rect 15964 6121 15998 6155
rect 360 6068 394 6102
rect 13194 6074 13228 6108
rect 13264 6074 13298 6108
rect 13334 6074 13368 6108
rect 13404 6074 13438 6108
rect 13474 6074 13508 6108
rect 13544 6074 13578 6108
rect 13614 6074 13648 6108
rect 13684 6074 13718 6108
rect 13754 6074 13788 6108
rect 13824 6074 13858 6108
rect 13894 6074 13928 6108
rect 13964 6074 13998 6108
rect 14034 6074 14068 6108
rect 14104 6074 14138 6108
rect 14174 6074 14208 6108
rect 14244 6074 14278 6108
rect 14314 6074 14348 6108
rect 14384 6074 14418 6108
rect 14454 6074 14488 6108
rect 14524 6074 14558 6108
rect 14594 6074 14628 6108
rect 14664 6074 14698 6108
rect 14774 6052 14808 6086
rect 14844 6052 14878 6086
rect 14914 6052 14948 6086
rect 14984 6052 15018 6086
rect 15054 6052 15088 6086
rect 15124 6052 15158 6086
rect 15194 6052 15228 6086
rect 15264 6052 15298 6086
rect 15334 6052 15368 6086
rect 15404 6052 15438 6086
rect 15474 6052 15508 6086
rect 15544 6052 15578 6086
rect 15614 6052 15648 6086
rect 15684 6052 15718 6086
rect 15754 6052 15788 6086
rect 15824 6052 15858 6086
rect 15894 6052 15928 6086
rect 15964 6052 15998 6086
rect 360 5999 394 6033
rect 429 5999 463 6033
rect 498 5999 532 6033
rect 567 5999 601 6033
rect 636 5999 670 6033
rect 705 5999 739 6033
rect 774 5999 808 6033
rect 843 5999 877 6033
rect 912 5999 946 6033
rect 981 5999 1015 6033
rect 1050 5999 1084 6033
rect 1119 5999 1153 6033
rect 1188 5999 1222 6033
rect 1257 5999 1291 6033
rect 1326 5999 1360 6033
rect 1395 5999 1429 6033
rect 1464 5999 1498 6033
rect 1533 5999 1567 6033
rect 1602 5999 1636 6033
rect 1671 5999 1705 6033
rect 1740 5999 1774 6033
rect 1809 5999 1843 6033
rect 1878 5999 1912 6033
rect 1947 5999 1981 6033
rect 2016 5999 2050 6033
rect 2085 5999 2119 6033
rect 2154 5999 2188 6033
rect 2223 5999 2257 6033
rect 2292 5999 2326 6033
rect 2361 5999 2395 6033
rect 2430 5999 2464 6033
rect 2499 5999 2533 6033
rect 2568 5999 2602 6033
rect 2637 5999 2671 6033
rect 2706 5999 2740 6033
rect 2775 5999 2809 6033
rect 2844 5999 2878 6033
rect 2913 5999 2947 6033
rect 2982 5999 3016 6033
rect 3051 5999 3085 6033
rect 3120 5999 3154 6033
rect 3189 5999 3223 6033
rect 3257 5999 3291 6033
rect 3325 5999 3359 6033
rect 3393 5999 3427 6033
rect 3461 5999 3495 6033
rect 3529 5999 3563 6033
rect 3597 5999 3631 6033
rect 3665 5999 3699 6033
rect 3733 5999 3767 6033
rect 3801 5999 3835 6033
rect 3869 5999 3903 6033
rect 3937 5999 3971 6033
rect 4005 5999 4039 6033
rect 4073 5999 4107 6033
rect 4141 5999 4175 6033
rect 4209 5999 4243 6033
rect 4277 5999 4311 6033
rect 4345 5999 4379 6033
rect 4413 5999 4447 6033
rect 4481 5999 4515 6033
rect 4549 5999 4583 6033
rect 4617 5999 4651 6033
rect 4685 5999 4719 6033
rect 4753 5999 4787 6033
rect 4821 5999 4855 6033
rect 4889 5999 4923 6033
rect 4957 5999 4991 6033
rect 5025 5999 5059 6033
rect 5093 5999 5127 6033
rect 5161 5999 5195 6033
rect 5229 5999 5263 6033
rect 5297 5999 5331 6033
rect 5365 5999 5399 6033
rect 5433 5999 5467 6033
rect 5501 5999 5535 6033
rect 5569 5999 5603 6033
rect 5637 5999 5671 6033
rect 5705 5999 5739 6033
rect 5773 5999 5807 6033
rect 5841 5999 5875 6033
rect 5909 5999 5943 6033
rect 5977 5999 6011 6033
rect 6045 5999 6079 6033
rect 6113 5999 6147 6033
rect 6181 5999 6215 6033
rect 6249 5999 6283 6033
rect 6317 5999 6351 6033
rect 6385 5999 6419 6033
rect 6453 5999 6487 6033
rect 6521 5999 6555 6033
rect 6589 5999 6623 6033
rect 6657 5999 6691 6033
rect 6725 5999 6759 6033
rect 6793 5999 6827 6033
rect 6861 5999 6895 6033
rect 6929 5999 6963 6033
rect 6997 5999 7031 6033
rect 7065 5999 7099 6033
rect 7133 5999 7167 6033
rect 7201 5999 7235 6033
rect 7269 5999 7303 6033
rect 7337 5999 7371 6033
rect 7405 5999 7439 6033
rect 7473 5999 7507 6033
rect 7541 5999 7575 6033
rect 7609 5999 7643 6033
rect 7677 5999 7711 6033
rect 7745 5999 7779 6033
rect 7813 5999 7847 6033
rect 7881 5999 7915 6033
rect 7949 5999 7983 6033
rect 8017 5999 8051 6033
rect 8085 5999 8119 6033
rect 8153 5999 8187 6033
rect 8221 5999 8255 6033
rect 8289 5999 8323 6033
rect 8357 5999 8391 6033
rect 8425 5999 8459 6033
rect 8493 5999 8527 6033
rect 8561 5999 8595 6033
rect 8629 5999 8663 6033
rect 8697 5999 8731 6033
rect 8765 5999 8799 6033
rect 8833 5999 8867 6033
rect 8901 5999 8935 6033
rect 8969 5999 9003 6033
rect 9037 5999 9071 6033
rect 9105 5999 9139 6033
rect 9173 5999 9207 6033
rect 9241 5999 9275 6033
rect 9309 5999 9343 6033
rect 9377 5999 9411 6033
rect 9445 5999 9479 6033
rect 9513 5999 9547 6033
rect 9581 5999 9615 6033
rect 9649 5999 9683 6033
rect 9717 5999 9751 6033
rect 9785 5999 9819 6033
rect 9853 5999 9887 6033
rect 9921 5999 9955 6033
rect 9989 5999 10023 6033
rect 10057 5999 10091 6033
rect 10125 5999 10159 6033
rect 10193 5999 10227 6033
rect 10261 5999 10295 6033
rect 10329 5999 10363 6033
rect 10397 5999 10431 6033
rect 10465 5999 10499 6033
rect 10533 5999 10567 6033
rect 10601 5999 10635 6033
rect 10669 5999 10703 6033
rect 10737 5999 10771 6033
rect 10805 5999 10839 6033
rect 10873 5999 10907 6033
rect 10941 5999 10975 6033
rect 11009 5999 11043 6033
rect 11077 5999 11111 6033
rect 11145 5999 11179 6033
rect 11213 5999 11247 6033
rect 11281 5999 11315 6033
rect 11349 5999 11383 6033
rect 11417 5999 11451 6033
rect 11485 5999 11519 6033
rect 11553 5999 11587 6033
rect 11621 5999 11655 6033
rect 11689 5999 11723 6033
rect 11757 5999 11791 6033
rect 11825 5999 11859 6033
rect 11893 5999 11927 6033
rect 11961 5999 11995 6033
rect 12029 5999 12063 6033
rect 12097 5999 12131 6033
rect 12165 5999 12199 6033
rect 12233 5999 12267 6033
rect 12301 5999 12335 6033
rect 12369 5999 12403 6033
rect 12437 5999 12471 6033
rect 12505 5999 12539 6033
rect 12573 5999 12607 6033
rect 12641 5999 12675 6033
rect 12709 5999 12743 6033
rect 12777 5999 12811 6033
rect 12845 5999 12879 6033
rect 12913 5999 12947 6033
rect 12981 5999 13015 6033
rect 13049 5999 13083 6033
rect 13117 5999 13151 6033
rect 13185 5999 13219 6033
rect 13253 5999 13287 6033
rect 13321 5999 13355 6033
rect 13389 5999 13423 6033
rect 13457 5999 13491 6033
rect 13525 5999 13559 6033
rect 13593 5999 13627 6033
rect 13661 5999 13695 6033
rect 13729 5999 13763 6033
rect 13797 5999 13831 6033
rect 13865 5999 13899 6033
rect 13933 5999 13967 6033
rect 14001 5999 14035 6033
rect 14069 5999 14103 6033
rect 14137 5999 14171 6033
rect 14205 5999 14239 6033
rect 14273 5999 14307 6033
rect 14341 5999 14375 6033
rect 14409 5999 14443 6033
rect 14477 5999 14511 6033
rect 14545 5999 14579 6033
rect 14613 5999 14647 6033
rect 14774 5983 14808 6017
rect 14844 5983 14878 6017
rect 14914 5983 14948 6017
rect 14984 5983 15018 6017
rect 15054 5983 15088 6017
rect 15124 5983 15158 6017
rect 15194 5983 15228 6017
rect 15264 5983 15298 6017
rect 15334 5983 15368 6017
rect 15404 5983 15438 6017
rect 15474 5983 15508 6017
rect 15544 5983 15578 6017
rect 15614 5983 15648 6017
rect 15684 5983 15718 6017
rect 15754 5983 15788 6017
rect 15824 5983 15858 6017
rect 15894 5983 15928 6017
rect 15964 5983 15998 6017
rect 11506 5917 11540 5951
rect 11506 5848 11540 5882
rect 14774 5914 14808 5948
rect 14844 5914 14878 5948
rect 14914 5914 14948 5948
rect 14984 5914 15018 5948
rect 15054 5914 15088 5948
rect 15124 5914 15158 5948
rect 15194 5914 15228 5948
rect 15264 5914 15298 5948
rect 15334 5914 15368 5948
rect 15404 5914 15438 5948
rect 15474 5914 15508 5948
rect 15544 5914 15578 5948
rect 15614 5914 15648 5948
rect 15684 5914 15718 5948
rect 15754 5914 15788 5948
rect 15824 5914 15858 5948
rect 15894 5914 15928 5948
rect 15964 5914 15998 5948
rect 14774 5845 14808 5879
rect 14844 5845 14878 5879
rect 14914 5845 14948 5879
rect 14984 5845 15018 5879
rect 15054 5845 15088 5879
rect 15124 5845 15158 5879
rect 15194 5845 15228 5879
rect 15264 5845 15298 5879
rect 15334 5845 15368 5879
rect 15404 5845 15438 5879
rect 15474 5845 15508 5879
rect 15544 5845 15578 5879
rect 15614 5845 15648 5879
rect 15684 5845 15718 5879
rect 15754 5845 15788 5879
rect 15824 5845 15858 5879
rect 15894 5845 15928 5879
rect 15964 5845 15998 5879
rect 11506 5779 11540 5813
rect 14774 5776 14808 5810
rect 14844 5776 14878 5810
rect 14914 5776 14948 5810
rect 14984 5776 15018 5810
rect 15054 5776 15088 5810
rect 15124 5776 15158 5810
rect 15194 5776 15228 5810
rect 15264 5776 15298 5810
rect 15334 5776 15368 5810
rect 15404 5776 15438 5810
rect 15474 5776 15508 5810
rect 15544 5776 15578 5810
rect 15614 5776 15648 5810
rect 15684 5776 15718 5810
rect 15754 5776 15788 5810
rect 15824 5776 15858 5810
rect 15894 5776 15928 5810
rect 15964 5776 15998 5810
rect 11506 5710 11540 5744
rect 11506 5641 11540 5675
rect 14774 5707 14808 5741
rect 14844 5707 14878 5741
rect 14914 5707 14948 5741
rect 14984 5707 15018 5741
rect 15054 5707 15088 5741
rect 15124 5707 15158 5741
rect 15194 5707 15228 5741
rect 15264 5707 15298 5741
rect 15334 5707 15368 5741
rect 15404 5707 15438 5741
rect 15474 5707 15508 5741
rect 15544 5707 15578 5741
rect 15614 5707 15648 5741
rect 15684 5707 15718 5741
rect 15754 5707 15788 5741
rect 15824 5707 15858 5741
rect 15894 5707 15928 5741
rect 15964 5707 15998 5741
rect 14774 5638 14808 5672
rect 14844 5638 14878 5672
rect 14914 5638 14948 5672
rect 14984 5638 15018 5672
rect 15054 5638 15088 5672
rect 15124 5638 15158 5672
rect 15194 5638 15228 5672
rect 15264 5638 15298 5672
rect 15334 5638 15368 5672
rect 15404 5638 15438 5672
rect 15474 5638 15508 5672
rect 15544 5638 15578 5672
rect 15614 5638 15648 5672
rect 15684 5638 15718 5672
rect 15754 5638 15788 5672
rect 15824 5638 15858 5672
rect 15894 5638 15928 5672
rect 15964 5638 15998 5672
rect 11506 5572 11540 5606
rect 11506 5503 11540 5537
rect 14774 5569 14808 5603
rect 14844 5569 14878 5603
rect 14914 5569 14948 5603
rect 14984 5569 15018 5603
rect 15054 5569 15088 5603
rect 15124 5569 15158 5603
rect 15194 5569 15228 5603
rect 15264 5569 15298 5603
rect 15334 5569 15368 5603
rect 15404 5569 15438 5603
rect 15474 5569 15508 5603
rect 15544 5569 15578 5603
rect 15614 5569 15648 5603
rect 15684 5569 15718 5603
rect 15754 5569 15788 5603
rect 15824 5569 15858 5603
rect 15894 5569 15928 5603
rect 15964 5569 15998 5603
rect 11506 5434 11540 5468
rect 14774 5500 14808 5534
rect 14844 5500 14878 5534
rect 14914 5500 14948 5534
rect 14984 5500 15018 5534
rect 15054 5500 15088 5534
rect 15124 5500 15158 5534
rect 15194 5500 15228 5534
rect 15264 5500 15298 5534
rect 15334 5500 15368 5534
rect 15404 5500 15438 5534
rect 15474 5500 15508 5534
rect 15544 5500 15578 5534
rect 15614 5500 15648 5534
rect 15684 5500 15718 5534
rect 15754 5500 15788 5534
rect 15824 5500 15858 5534
rect 15894 5500 15928 5534
rect 15964 5500 15998 5534
rect 11506 5365 11540 5399
rect 14774 5431 14808 5465
rect 14844 5431 14878 5465
rect 14914 5431 14948 5465
rect 14984 5431 15018 5465
rect 15054 5431 15088 5465
rect 15124 5431 15158 5465
rect 15194 5431 15228 5465
rect 15264 5431 15298 5465
rect 15334 5431 15368 5465
rect 15404 5431 15438 5465
rect 15474 5431 15508 5465
rect 15544 5431 15578 5465
rect 15614 5431 15648 5465
rect 15684 5431 15718 5465
rect 15754 5431 15788 5465
rect 15824 5431 15858 5465
rect 15894 5431 15928 5465
rect 15964 5431 15998 5465
rect 14774 5362 14808 5396
rect 14844 5362 14878 5396
rect 14914 5362 14948 5396
rect 14984 5362 15018 5396
rect 15054 5362 15088 5396
rect 15124 5362 15158 5396
rect 15194 5362 15228 5396
rect 15264 5362 15298 5396
rect 15334 5362 15368 5396
rect 15404 5362 15438 5396
rect 15474 5362 15508 5396
rect 15544 5362 15578 5396
rect 15614 5362 15648 5396
rect 15684 5362 15718 5396
rect 15754 5362 15788 5396
rect 15824 5362 15858 5396
rect 15894 5362 15928 5396
rect 15964 5362 15998 5396
rect 11506 5296 11540 5330
rect 11506 5227 11540 5261
rect 14774 5293 14808 5327
rect 14844 5293 14878 5327
rect 14914 5293 14948 5327
rect 14984 5293 15018 5327
rect 15054 5293 15088 5327
rect 15124 5293 15158 5327
rect 15194 5293 15228 5327
rect 15264 5293 15298 5327
rect 15334 5293 15368 5327
rect 15404 5293 15438 5327
rect 15474 5293 15508 5327
rect 15544 5293 15578 5327
rect 15614 5293 15648 5327
rect 15684 5293 15718 5327
rect 15754 5293 15788 5327
rect 15824 5293 15858 5327
rect 15894 5293 15928 5327
rect 15964 5293 15998 5327
rect 14774 5224 14808 5258
rect 14844 5224 14878 5258
rect 14914 5224 14948 5258
rect 14984 5224 15018 5258
rect 15054 5224 15088 5258
rect 15124 5224 15158 5258
rect 15194 5224 15228 5258
rect 15264 5224 15298 5258
rect 15334 5224 15368 5258
rect 15404 5224 15438 5258
rect 15474 5224 15508 5258
rect 15544 5224 15578 5258
rect 15614 5224 15648 5258
rect 15684 5224 15718 5258
rect 15754 5224 15788 5258
rect 15824 5224 15858 5258
rect 15894 5224 15928 5258
rect 15964 5224 15998 5258
rect 11506 5158 11540 5192
rect 14774 5156 14808 5190
rect 14844 5156 14878 5190
rect 14914 5156 14948 5190
rect 14984 5156 15018 5190
rect 15054 5156 15088 5190
rect 15124 5156 15158 5190
rect 15194 5156 15228 5190
rect 15264 5156 15298 5190
rect 15334 5156 15368 5190
rect 15404 5156 15438 5190
rect 15474 5156 15508 5190
rect 15544 5156 15578 5190
rect 15614 5156 15648 5190
rect 15684 5156 15718 5190
rect 15754 5156 15788 5190
rect 15824 5156 15858 5190
rect 15894 5156 15928 5190
rect 15964 5156 15998 5190
rect 11506 5089 11540 5123
rect 11506 5020 11540 5054
rect 14774 5088 14808 5122
rect 14844 5088 14878 5122
rect 14914 5088 14948 5122
rect 14984 5088 15018 5122
rect 15054 5088 15088 5122
rect 15124 5088 15158 5122
rect 15194 5088 15228 5122
rect 15264 5088 15298 5122
rect 15334 5088 15368 5122
rect 15404 5088 15438 5122
rect 15474 5088 15508 5122
rect 15544 5088 15578 5122
rect 15614 5088 15648 5122
rect 15684 5088 15718 5122
rect 15754 5088 15788 5122
rect 15824 5088 15858 5122
rect 15894 5088 15928 5122
rect 15964 5088 15998 5122
rect 14774 5020 14808 5054
rect 14844 5020 14878 5054
rect 14914 5020 14948 5054
rect 14984 5020 15018 5054
rect 15054 5020 15088 5054
rect 15124 5020 15158 5054
rect 15194 5020 15228 5054
rect 15264 5020 15298 5054
rect 15334 5020 15368 5054
rect 15404 5020 15438 5054
rect 15474 5020 15508 5054
rect 15544 5020 15578 5054
rect 15614 5020 15648 5054
rect 15684 5020 15718 5054
rect 15754 5020 15788 5054
rect 15824 5020 15858 5054
rect 15894 5020 15928 5054
rect 15964 5020 15998 5054
rect 11506 4951 11540 4985
rect 11506 4882 11540 4916
rect 14774 4952 14808 4986
rect 14844 4952 14878 4986
rect 14914 4952 14948 4986
rect 14984 4952 15018 4986
rect 15054 4952 15088 4986
rect 15124 4952 15158 4986
rect 15194 4952 15228 4986
rect 15264 4952 15298 4986
rect 15334 4952 15368 4986
rect 15404 4952 15438 4986
rect 15474 4952 15508 4986
rect 15544 4952 15578 4986
rect 15614 4952 15648 4986
rect 15684 4952 15718 4986
rect 15754 4952 15788 4986
rect 15824 4952 15858 4986
rect 15894 4952 15928 4986
rect 15964 4952 15998 4986
rect 11506 4813 11540 4847
rect 14774 4884 14808 4918
rect 14844 4884 14878 4918
rect 14914 4884 14948 4918
rect 14984 4884 15018 4918
rect 15054 4884 15088 4918
rect 15124 4884 15158 4918
rect 15194 4884 15228 4918
rect 15264 4884 15298 4918
rect 15334 4884 15368 4918
rect 15404 4884 15438 4918
rect 15474 4884 15508 4918
rect 15544 4884 15578 4918
rect 15614 4884 15648 4918
rect 15684 4884 15718 4918
rect 15754 4884 15788 4918
rect 15824 4884 15858 4918
rect 15894 4884 15928 4918
rect 15964 4884 15998 4918
rect 11506 4744 11540 4778
rect 14774 4816 14808 4850
rect 14844 4816 14878 4850
rect 14914 4816 14948 4850
rect 14984 4816 15018 4850
rect 15054 4816 15088 4850
rect 15124 4816 15158 4850
rect 15194 4816 15228 4850
rect 15264 4816 15298 4850
rect 15334 4816 15368 4850
rect 15404 4816 15438 4850
rect 15474 4816 15508 4850
rect 15544 4816 15578 4850
rect 15614 4816 15648 4850
rect 15684 4816 15718 4850
rect 15754 4816 15788 4850
rect 15824 4816 15858 4850
rect 15894 4816 15928 4850
rect 15964 4816 15998 4850
rect 14774 4748 14808 4782
rect 14844 4748 14878 4782
rect 14914 4748 14948 4782
rect 14984 4748 15018 4782
rect 15054 4748 15088 4782
rect 15124 4748 15158 4782
rect 15194 4748 15228 4782
rect 15264 4748 15298 4782
rect 15334 4748 15368 4782
rect 15404 4748 15438 4782
rect 15474 4748 15508 4782
rect 15544 4748 15578 4782
rect 15614 4748 15648 4782
rect 15684 4748 15718 4782
rect 15754 4748 15788 4782
rect 15824 4748 15858 4782
rect 15894 4748 15928 4782
rect 15964 4748 15998 4782
rect 11506 4675 11540 4709
rect 11506 4606 11540 4640
rect 14774 4680 14808 4714
rect 14844 4680 14878 4714
rect 14914 4680 14948 4714
rect 14984 4680 15018 4714
rect 15054 4680 15088 4714
rect 15124 4680 15158 4714
rect 15194 4680 15228 4714
rect 15264 4680 15298 4714
rect 15334 4680 15368 4714
rect 15404 4680 15438 4714
rect 15474 4680 15508 4714
rect 15544 4680 15578 4714
rect 15614 4680 15648 4714
rect 15684 4680 15718 4714
rect 15754 4680 15788 4714
rect 15824 4680 15858 4714
rect 15894 4680 15928 4714
rect 15964 4680 15998 4714
rect 14774 4612 14808 4646
rect 14844 4612 14878 4646
rect 14914 4612 14948 4646
rect 14984 4612 15018 4646
rect 15054 4612 15088 4646
rect 15124 4612 15158 4646
rect 15194 4612 15228 4646
rect 15264 4612 15298 4646
rect 15334 4612 15368 4646
rect 15404 4612 15438 4646
rect 15474 4612 15508 4646
rect 15544 4612 15578 4646
rect 15614 4612 15648 4646
rect 15684 4612 15718 4646
rect 15754 4612 15788 4646
rect 15824 4612 15858 4646
rect 15894 4612 15928 4646
rect 15964 4612 15998 4646
rect 11506 4537 11540 4571
rect 14774 4544 14808 4578
rect 14844 4544 14878 4578
rect 14914 4544 14948 4578
rect 14984 4544 15018 4578
rect 15054 4544 15088 4578
rect 15124 4544 15158 4578
rect 15194 4544 15228 4578
rect 15264 4544 15298 4578
rect 15334 4544 15368 4578
rect 15404 4544 15438 4578
rect 15474 4544 15508 4578
rect 15544 4544 15578 4578
rect 15614 4544 15648 4578
rect 15684 4544 15718 4578
rect 15754 4544 15788 4578
rect 15824 4544 15858 4578
rect 15894 4544 15928 4578
rect 15964 4544 15998 4578
rect 11506 4468 11540 4502
rect 14774 4476 14808 4510
rect 14844 4476 14878 4510
rect 14914 4476 14948 4510
rect 14984 4476 15018 4510
rect 15054 4476 15088 4510
rect 15124 4476 15158 4510
rect 15194 4476 15228 4510
rect 15264 4476 15298 4510
rect 15334 4476 15368 4510
rect 15404 4476 15438 4510
rect 15474 4476 15508 4510
rect 15544 4476 15578 4510
rect 15614 4476 15648 4510
rect 15684 4476 15718 4510
rect 15754 4476 15788 4510
rect 15824 4476 15858 4510
rect 15894 4476 15928 4510
rect 15964 4476 15998 4510
rect 11506 4399 11540 4433
rect 14774 4408 14808 4442
rect 14844 4408 14878 4442
rect 14914 4408 14948 4442
rect 14984 4408 15018 4442
rect 15054 4408 15088 4442
rect 15124 4408 15158 4442
rect 15194 4408 15228 4442
rect 15264 4408 15298 4442
rect 15334 4408 15368 4442
rect 15404 4408 15438 4442
rect 15474 4408 15508 4442
rect 15544 4408 15578 4442
rect 15614 4408 15648 4442
rect 15684 4408 15718 4442
rect 15754 4408 15788 4442
rect 15824 4408 15858 4442
rect 15894 4408 15928 4442
rect 15964 4408 15998 4442
rect 11506 4330 11540 4364
rect 11506 4261 11540 4295
rect 14774 4340 14808 4374
rect 14844 4340 14878 4374
rect 14914 4340 14948 4374
rect 14984 4340 15018 4374
rect 15054 4340 15088 4374
rect 15124 4340 15158 4374
rect 15194 4340 15228 4374
rect 15264 4340 15298 4374
rect 15334 4340 15368 4374
rect 15404 4340 15438 4374
rect 15474 4340 15508 4374
rect 15544 4340 15578 4374
rect 15614 4340 15648 4374
rect 15684 4340 15718 4374
rect 15754 4340 15788 4374
rect 15824 4340 15858 4374
rect 15894 4340 15928 4374
rect 15964 4340 15998 4374
rect 14774 4272 14808 4306
rect 14844 4272 14878 4306
rect 14914 4272 14948 4306
rect 14984 4272 15018 4306
rect 15054 4272 15088 4306
rect 15124 4272 15158 4306
rect 15194 4272 15228 4306
rect 15264 4272 15298 4306
rect 15334 4272 15368 4306
rect 15404 4272 15438 4306
rect 15474 4272 15508 4306
rect 15544 4272 15578 4306
rect 15614 4272 15648 4306
rect 15684 4272 15718 4306
rect 15754 4272 15788 4306
rect 15824 4272 15858 4306
rect 15894 4272 15928 4306
rect 15964 4272 15998 4306
rect 11506 4192 11540 4226
rect 11506 4123 11540 4157
rect 14774 4204 14808 4238
rect 14844 4204 14878 4238
rect 14914 4204 14948 4238
rect 14984 4204 15018 4238
rect 15054 4204 15088 4238
rect 15124 4204 15158 4238
rect 15194 4204 15228 4238
rect 15264 4204 15298 4238
rect 15334 4204 15368 4238
rect 15404 4204 15438 4238
rect 15474 4204 15508 4238
rect 15544 4204 15578 4238
rect 15614 4204 15648 4238
rect 15684 4204 15718 4238
rect 15754 4204 15788 4238
rect 15824 4204 15858 4238
rect 15894 4204 15928 4238
rect 15964 4204 15998 4238
rect 14774 4136 14808 4170
rect 14844 4136 14878 4170
rect 14914 4136 14948 4170
rect 14984 4136 15018 4170
rect 15054 4136 15088 4170
rect 15124 4136 15158 4170
rect 15194 4136 15228 4170
rect 15264 4136 15298 4170
rect 15334 4136 15368 4170
rect 15404 4136 15438 4170
rect 15474 4136 15508 4170
rect 15544 4136 15578 4170
rect 15614 4136 15648 4170
rect 15684 4136 15718 4170
rect 15754 4136 15788 4170
rect 15824 4136 15858 4170
rect 15894 4136 15928 4170
rect 15964 4136 15998 4170
rect 11506 4054 11540 4088
rect 14774 4068 14808 4102
rect 14844 4068 14878 4102
rect 14914 4068 14948 4102
rect 14984 4068 15018 4102
rect 15054 4068 15088 4102
rect 15124 4068 15158 4102
rect 15194 4068 15228 4102
rect 15264 4068 15298 4102
rect 15334 4068 15368 4102
rect 15404 4068 15438 4102
rect 15474 4068 15508 4102
rect 15544 4068 15578 4102
rect 15614 4068 15648 4102
rect 15684 4068 15718 4102
rect 15754 4068 15788 4102
rect 15824 4068 15858 4102
rect 15894 4068 15928 4102
rect 15964 4068 15998 4102
rect 11506 3985 11540 4019
rect 11588 4017 11622 4051
rect 11657 4017 11691 4051
rect 11726 4017 11760 4051
rect 11795 4017 11829 4051
rect 11864 4017 11898 4051
rect 11933 4017 11967 4051
rect 12002 4017 12036 4051
rect 12071 4017 12105 4051
rect 12140 4017 12174 4051
rect 12209 4017 12243 4051
rect 12278 4017 12312 4051
rect 12347 4017 12381 4051
rect 12416 4017 12450 4051
rect 12485 4017 12519 4051
rect 12554 4017 12588 4051
rect 12623 4017 12657 4051
rect 12692 4017 12726 4051
rect 12761 4017 12795 4051
rect 12830 4017 12864 4051
rect 12899 4017 12933 4051
rect 12968 4017 13002 4051
rect 13037 4017 13071 4051
rect 13106 4017 13140 4051
rect 13175 4017 13209 4051
rect 13244 4017 13278 4051
rect 13313 4017 13347 4051
rect 13382 4017 13416 4051
rect 13451 4017 13485 4051
rect 13520 4017 13554 4051
rect 13589 4017 13623 4051
rect 13658 4017 13692 4051
rect 13727 4017 13761 4051
rect 13796 4017 13830 4051
rect 13865 4017 13899 4051
rect 13934 4017 13968 4051
rect 14002 4017 14036 4051
rect 14070 4017 14104 4051
rect 14138 4017 14172 4051
rect 14206 4017 14240 4051
rect 14274 4017 14308 4051
rect 14342 4017 14376 4051
rect 14410 4017 14444 4051
rect 14478 4017 14512 4051
rect 14546 4017 14580 4051
rect 14614 4017 14648 4051
rect 14682 4017 14716 4051
rect 11506 3916 11540 3950
rect 14774 4000 14808 4034
rect 14844 4000 14878 4034
rect 14914 4000 14948 4034
rect 14984 4000 15018 4034
rect 15054 4000 15088 4034
rect 15124 4000 15158 4034
rect 15194 4000 15228 4034
rect 15264 4000 15298 4034
rect 15334 4000 15368 4034
rect 15404 4000 15438 4034
rect 15474 4000 15508 4034
rect 15544 4000 15578 4034
rect 15614 4000 15648 4034
rect 15684 4000 15718 4034
rect 15754 4000 15788 4034
rect 15824 4000 15858 4034
rect 15894 4000 15928 4034
rect 15964 4000 15998 4034
rect 11506 3847 11540 3881
rect 14774 3932 14808 3966
rect 14844 3932 14878 3966
rect 14914 3932 14948 3966
rect 14984 3932 15018 3966
rect 15054 3932 15088 3966
rect 15124 3932 15158 3966
rect 15194 3932 15228 3966
rect 15264 3932 15298 3966
rect 15334 3932 15368 3966
rect 15404 3932 15438 3966
rect 15474 3932 15508 3966
rect 15544 3932 15578 3966
rect 15614 3932 15648 3966
rect 15684 3932 15718 3966
rect 15754 3932 15788 3966
rect 15824 3932 15858 3966
rect 15894 3932 15928 3966
rect 15964 3932 15998 3966
rect 14774 3864 14808 3898
rect 14844 3864 14878 3898
rect 14914 3864 14948 3898
rect 14984 3864 15018 3898
rect 15054 3864 15088 3898
rect 15124 3864 15158 3898
rect 15194 3864 15228 3898
rect 15264 3864 15298 3898
rect 15334 3864 15368 3898
rect 15404 3864 15438 3898
rect 15474 3864 15508 3898
rect 15544 3864 15578 3898
rect 15614 3864 15648 3898
rect 15684 3864 15718 3898
rect 15754 3864 15788 3898
rect 15824 3864 15858 3898
rect 15894 3864 15928 3898
rect 15964 3864 15998 3898
rect 11506 3778 11540 3812
rect 14774 3796 14808 3830
rect 14844 3796 14878 3830
rect 14914 3796 14948 3830
rect 14984 3796 15018 3830
rect 15054 3796 15088 3830
rect 15124 3796 15158 3830
rect 15194 3796 15228 3830
rect 15264 3796 15298 3830
rect 15334 3796 15368 3830
rect 15404 3796 15438 3830
rect 15474 3796 15508 3830
rect 15544 3796 15578 3830
rect 15614 3796 15648 3830
rect 15684 3796 15718 3830
rect 15754 3796 15788 3830
rect 15824 3796 15858 3830
rect 15894 3796 15928 3830
rect 15964 3796 15998 3830
rect 11506 3709 11540 3743
rect 14774 3728 14808 3762
rect 14844 3728 14878 3762
rect 14914 3728 14948 3762
rect 14984 3728 15018 3762
rect 15054 3728 15088 3762
rect 15124 3728 15158 3762
rect 15194 3728 15228 3762
rect 15264 3728 15298 3762
rect 15334 3728 15368 3762
rect 15404 3728 15438 3762
rect 15474 3728 15508 3762
rect 15544 3728 15578 3762
rect 15614 3728 15648 3762
rect 15684 3728 15718 3762
rect 15754 3728 15788 3762
rect 15824 3728 15858 3762
rect 15894 3728 15928 3762
rect 15964 3728 15998 3762
rect 11506 3640 11540 3674
rect 14774 3660 14808 3694
rect 14844 3660 14878 3694
rect 14914 3660 14948 3694
rect 14984 3660 15018 3694
rect 15054 3660 15088 3694
rect 15124 3660 15158 3694
rect 15194 3660 15228 3694
rect 15264 3660 15298 3694
rect 15334 3660 15368 3694
rect 15404 3660 15438 3694
rect 15474 3660 15508 3694
rect 15544 3660 15578 3694
rect 15614 3660 15648 3694
rect 15684 3660 15718 3694
rect 15754 3660 15788 3694
rect 15824 3660 15858 3694
rect 15894 3660 15928 3694
rect 15964 3660 15998 3694
rect 11506 3571 11540 3605
rect 11506 3502 11540 3536
rect 14774 3592 14808 3626
rect 14844 3592 14878 3626
rect 14914 3592 14948 3626
rect 14984 3592 15018 3626
rect 15054 3592 15088 3626
rect 15124 3592 15158 3626
rect 15194 3592 15228 3626
rect 15264 3592 15298 3626
rect 15334 3592 15368 3626
rect 15404 3592 15438 3626
rect 15474 3592 15508 3626
rect 15544 3592 15578 3626
rect 15614 3592 15648 3626
rect 15684 3592 15718 3626
rect 15754 3592 15788 3626
rect 15824 3592 15858 3626
rect 15894 3592 15928 3626
rect 15964 3592 15998 3626
rect 14774 3524 14808 3558
rect 14844 3524 14878 3558
rect 14914 3524 14948 3558
rect 14984 3524 15018 3558
rect 15054 3524 15088 3558
rect 15124 3524 15158 3558
rect 15194 3524 15228 3558
rect 15264 3524 15298 3558
rect 15334 3524 15368 3558
rect 15404 3524 15438 3558
rect 15474 3524 15508 3558
rect 15544 3524 15578 3558
rect 15614 3524 15648 3558
rect 15684 3524 15718 3558
rect 15754 3524 15788 3558
rect 15824 3524 15858 3558
rect 15894 3524 15928 3558
rect 15964 3524 15998 3558
rect 11506 3433 11540 3467
rect 11506 3364 11540 3398
rect 14774 3456 14808 3490
rect 14844 3456 14878 3490
rect 14914 3456 14948 3490
rect 14984 3456 15018 3490
rect 15054 3456 15088 3490
rect 15124 3456 15158 3490
rect 15194 3456 15228 3490
rect 15264 3456 15298 3490
rect 15334 3456 15368 3490
rect 15404 3456 15438 3490
rect 15474 3456 15508 3490
rect 15544 3456 15578 3490
rect 15614 3456 15648 3490
rect 15684 3456 15718 3490
rect 15754 3456 15788 3490
rect 15824 3456 15858 3490
rect 15894 3456 15928 3490
rect 15964 3456 15998 3490
rect 14774 3388 14808 3422
rect 14844 3388 14878 3422
rect 14914 3388 14948 3422
rect 14984 3388 15018 3422
rect 15054 3388 15088 3422
rect 15124 3388 15158 3422
rect 15194 3388 15228 3422
rect 15264 3388 15298 3422
rect 15334 3388 15368 3422
rect 15404 3388 15438 3422
rect 15474 3388 15508 3422
rect 15544 3388 15578 3422
rect 15614 3388 15648 3422
rect 15684 3388 15718 3422
rect 15754 3388 15788 3422
rect 15824 3388 15858 3422
rect 15894 3388 15928 3422
rect 15964 3388 15998 3422
rect 11506 3295 11540 3329
rect 11506 3226 11540 3260
rect 14774 3320 14808 3354
rect 14844 3320 14878 3354
rect 14914 3320 14948 3354
rect 14984 3320 15018 3354
rect 15054 3320 15088 3354
rect 15124 3320 15158 3354
rect 15194 3320 15228 3354
rect 15264 3320 15298 3354
rect 15334 3320 15368 3354
rect 15404 3320 15438 3354
rect 15474 3320 15508 3354
rect 15544 3320 15578 3354
rect 15614 3320 15648 3354
rect 15684 3320 15718 3354
rect 15754 3320 15788 3354
rect 15824 3320 15858 3354
rect 15894 3320 15928 3354
rect 15964 3320 15998 3354
rect 14774 3252 14808 3286
rect 14844 3252 14878 3286
rect 14914 3252 14948 3286
rect 14984 3252 15018 3286
rect 15054 3252 15088 3286
rect 15124 3252 15158 3286
rect 15194 3252 15228 3286
rect 15264 3252 15298 3286
rect 15334 3252 15368 3286
rect 15404 3252 15438 3286
rect 15474 3252 15508 3286
rect 15544 3252 15578 3286
rect 15614 3252 15648 3286
rect 15684 3252 15718 3286
rect 15754 3252 15788 3286
rect 15824 3252 15858 3286
rect 15894 3252 15928 3286
rect 15964 3252 15998 3286
rect 11506 3157 11540 3191
rect 14774 3184 14808 3218
rect 14844 3184 14878 3218
rect 14914 3184 14948 3218
rect 14984 3184 15018 3218
rect 15054 3184 15088 3218
rect 15124 3184 15158 3218
rect 15194 3184 15228 3218
rect 15264 3184 15298 3218
rect 15334 3184 15368 3218
rect 15404 3184 15438 3218
rect 15474 3184 15508 3218
rect 15544 3184 15578 3218
rect 15614 3184 15648 3218
rect 15684 3184 15718 3218
rect 15754 3184 15788 3218
rect 15824 3184 15858 3218
rect 15894 3184 15928 3218
rect 15964 3184 15998 3218
rect 11506 3088 11540 3122
rect 14774 3116 14808 3150
rect 14844 3116 14878 3150
rect 14914 3116 14948 3150
rect 14984 3116 15018 3150
rect 15054 3116 15088 3150
rect 15124 3116 15158 3150
rect 15194 3116 15228 3150
rect 15264 3116 15298 3150
rect 15334 3116 15368 3150
rect 15404 3116 15438 3150
rect 15474 3116 15508 3150
rect 15544 3116 15578 3150
rect 15614 3116 15648 3150
rect 15684 3116 15718 3150
rect 15754 3116 15788 3150
rect 15824 3116 15858 3150
rect 15894 3116 15928 3150
rect 15964 3116 15998 3150
rect 11506 3019 11540 3053
rect 14774 3048 14808 3082
rect 14844 3048 14878 3082
rect 14914 3048 14948 3082
rect 14984 3048 15018 3082
rect 15054 3048 15088 3082
rect 15124 3048 15158 3082
rect 15194 3048 15228 3082
rect 15264 3048 15298 3082
rect 15334 3048 15368 3082
rect 15404 3048 15438 3082
rect 15474 3048 15508 3082
rect 15544 3048 15578 3082
rect 15614 3048 15648 3082
rect 15684 3048 15718 3082
rect 15754 3048 15788 3082
rect 15824 3048 15858 3082
rect 15894 3048 15928 3082
rect 15964 3048 15998 3082
rect 11506 2950 11540 2984
rect 14774 2980 14808 3014
rect 14844 2980 14878 3014
rect 14914 2980 14948 3014
rect 14984 2980 15018 3014
rect 15054 2980 15088 3014
rect 15124 2980 15158 3014
rect 15194 2980 15228 3014
rect 15264 2980 15298 3014
rect 15334 2980 15368 3014
rect 15404 2980 15438 3014
rect 15474 2980 15508 3014
rect 15544 2980 15578 3014
rect 15614 2980 15648 3014
rect 15684 2980 15718 3014
rect 15754 2980 15788 3014
rect 15824 2980 15858 3014
rect 15894 2980 15928 3014
rect 15964 2980 15998 3014
rect 11506 2881 11540 2915
rect 14774 2912 14808 2946
rect 14844 2912 14878 2946
rect 14914 2912 14948 2946
rect 14984 2912 15018 2946
rect 15054 2912 15088 2946
rect 15124 2912 15158 2946
rect 15194 2912 15228 2946
rect 15264 2912 15298 2946
rect 15334 2912 15368 2946
rect 15404 2912 15438 2946
rect 15474 2912 15508 2946
rect 15544 2912 15578 2946
rect 15614 2912 15648 2946
rect 15684 2912 15718 2946
rect 15754 2912 15788 2946
rect 15824 2912 15858 2946
rect 15894 2912 15928 2946
rect 15964 2912 15998 2946
rect 11506 2812 11540 2846
rect 11506 2743 11540 2777
rect 14774 2844 14808 2878
rect 14844 2844 14878 2878
rect 14914 2844 14948 2878
rect 14984 2844 15018 2878
rect 15054 2844 15088 2878
rect 15124 2844 15158 2878
rect 15194 2844 15228 2878
rect 15264 2844 15298 2878
rect 15334 2844 15368 2878
rect 15404 2844 15438 2878
rect 15474 2844 15508 2878
rect 15544 2844 15578 2878
rect 15614 2844 15648 2878
rect 15684 2844 15718 2878
rect 15754 2844 15788 2878
rect 15824 2844 15858 2878
rect 15894 2844 15928 2878
rect 15964 2844 15998 2878
rect 14774 2776 14808 2810
rect 14844 2776 14878 2810
rect 14914 2776 14948 2810
rect 14984 2776 15018 2810
rect 15054 2776 15088 2810
rect 15124 2776 15158 2810
rect 15194 2776 15228 2810
rect 15264 2776 15298 2810
rect 15334 2776 15368 2810
rect 15404 2776 15438 2810
rect 15474 2776 15508 2810
rect 15544 2776 15578 2810
rect 15614 2776 15648 2810
rect 15684 2776 15718 2810
rect 15754 2776 15788 2810
rect 15824 2776 15858 2810
rect 15894 2776 15928 2810
rect 15964 2776 15998 2810
rect 11506 2674 11540 2708
rect 11506 2605 11540 2639
rect 14774 2708 14808 2742
rect 14844 2708 14878 2742
rect 14914 2708 14948 2742
rect 14984 2708 15018 2742
rect 15054 2708 15088 2742
rect 15124 2708 15158 2742
rect 15194 2708 15228 2742
rect 15264 2708 15298 2742
rect 15334 2708 15368 2742
rect 15404 2708 15438 2742
rect 15474 2708 15508 2742
rect 15544 2708 15578 2742
rect 15614 2708 15648 2742
rect 15684 2708 15718 2742
rect 15754 2708 15788 2742
rect 15824 2708 15858 2742
rect 15894 2708 15928 2742
rect 15964 2708 15998 2742
rect 14774 2640 14808 2674
rect 14844 2640 14878 2674
rect 14914 2640 14948 2674
rect 14984 2640 15018 2674
rect 15054 2640 15088 2674
rect 15124 2640 15158 2674
rect 15194 2640 15228 2674
rect 15264 2640 15298 2674
rect 15334 2640 15368 2674
rect 15404 2640 15438 2674
rect 15474 2640 15508 2674
rect 15544 2640 15578 2674
rect 15614 2640 15648 2674
rect 15684 2640 15718 2674
rect 15754 2640 15788 2674
rect 15824 2640 15858 2674
rect 15894 2640 15928 2674
rect 15964 2640 15998 2674
rect 11506 2536 11540 2570
rect 14774 2572 14808 2606
rect 14844 2572 14878 2606
rect 14914 2572 14948 2606
rect 14984 2572 15018 2606
rect 15054 2572 15088 2606
rect 15124 2572 15158 2606
rect 15194 2572 15228 2606
rect 15264 2572 15298 2606
rect 15334 2572 15368 2606
rect 15404 2572 15438 2606
rect 15474 2572 15508 2606
rect 15544 2572 15578 2606
rect 15614 2572 15648 2606
rect 15684 2572 15718 2606
rect 15754 2572 15788 2606
rect 15824 2572 15858 2606
rect 15894 2572 15928 2606
rect 15964 2572 15998 2606
rect 11506 2467 11540 2501
rect 14774 2504 14808 2538
rect 14844 2504 14878 2538
rect 14914 2504 14948 2538
rect 14984 2504 15018 2538
rect 15054 2504 15088 2538
rect 15124 2504 15158 2538
rect 15194 2504 15228 2538
rect 15264 2504 15298 2538
rect 15334 2504 15368 2538
rect 15404 2504 15438 2538
rect 15474 2504 15508 2538
rect 15544 2504 15578 2538
rect 15614 2504 15648 2538
rect 15684 2504 15718 2538
rect 15754 2504 15788 2538
rect 15824 2504 15858 2538
rect 15894 2504 15928 2538
rect 15964 2504 15998 2538
rect 11506 2397 11540 2431
rect 14774 2436 14808 2470
rect 14844 2436 14878 2470
rect 14914 2436 14948 2470
rect 14984 2436 15018 2470
rect 15054 2436 15088 2470
rect 15124 2436 15158 2470
rect 15194 2436 15228 2470
rect 15264 2436 15298 2470
rect 15334 2436 15368 2470
rect 15404 2436 15438 2470
rect 15474 2436 15508 2470
rect 15544 2436 15578 2470
rect 15614 2436 15648 2470
rect 15684 2436 15718 2470
rect 15754 2436 15788 2470
rect 15824 2436 15858 2470
rect 15894 2436 15928 2470
rect 15964 2436 15998 2470
rect 11506 2327 11540 2361
rect 14774 2368 14808 2402
rect 14844 2368 14878 2402
rect 14914 2368 14948 2402
rect 14984 2368 15018 2402
rect 15054 2368 15088 2402
rect 15124 2368 15158 2402
rect 15194 2368 15228 2402
rect 15264 2368 15298 2402
rect 15334 2368 15368 2402
rect 15404 2368 15438 2402
rect 15474 2368 15508 2402
rect 15544 2368 15578 2402
rect 15614 2368 15648 2402
rect 15684 2368 15718 2402
rect 15754 2368 15788 2402
rect 15824 2368 15858 2402
rect 15894 2368 15928 2402
rect 15964 2368 15998 2402
rect 11506 2257 11540 2291
rect 14774 2300 14808 2334
rect 14844 2300 14878 2334
rect 14914 2300 14948 2334
rect 14984 2300 15018 2334
rect 15054 2300 15088 2334
rect 15124 2300 15158 2334
rect 15194 2300 15228 2334
rect 15264 2300 15298 2334
rect 15334 2300 15368 2334
rect 15404 2300 15438 2334
rect 15474 2300 15508 2334
rect 15544 2300 15578 2334
rect 15614 2300 15648 2334
rect 15684 2300 15718 2334
rect 15754 2300 15788 2334
rect 15824 2300 15858 2334
rect 15894 2300 15928 2334
rect 15964 2300 15998 2334
rect 11506 2187 11540 2221
rect 11506 2117 11540 2151
rect 14774 2232 14808 2266
rect 14844 2232 14878 2266
rect 14914 2232 14948 2266
rect 14984 2232 15018 2266
rect 15054 2232 15088 2266
rect 15124 2232 15158 2266
rect 15194 2232 15228 2266
rect 15264 2232 15298 2266
rect 15334 2232 15368 2266
rect 15404 2232 15438 2266
rect 15474 2232 15508 2266
rect 15544 2232 15578 2266
rect 15614 2232 15648 2266
rect 15684 2232 15718 2266
rect 15754 2232 15788 2266
rect 15824 2232 15858 2266
rect 15894 2232 15928 2266
rect 15964 2232 15998 2266
rect 14774 2164 14808 2198
rect 14844 2164 14878 2198
rect 14914 2164 14948 2198
rect 14984 2164 15018 2198
rect 15054 2164 15088 2198
rect 15124 2164 15158 2198
rect 15194 2164 15228 2198
rect 15264 2164 15298 2198
rect 15334 2164 15368 2198
rect 15404 2164 15438 2198
rect 15474 2164 15508 2198
rect 15544 2164 15578 2198
rect 15614 2164 15648 2198
rect 15684 2164 15718 2198
rect 15754 2164 15788 2198
rect 15824 2164 15858 2198
rect 15894 2164 15928 2198
rect 15964 2164 15998 2198
rect 14774 2096 14808 2130
rect 14844 2096 14878 2130
rect 14914 2096 14948 2130
rect 14984 2096 15018 2130
rect 15054 2096 15088 2130
rect 15124 2096 15158 2130
rect 15194 2096 15228 2130
rect 15264 2096 15298 2130
rect 15334 2096 15368 2130
rect 15404 2096 15438 2130
rect 15474 2096 15508 2130
rect 15544 2096 15578 2130
rect 15614 2096 15648 2130
rect 15684 2096 15718 2130
rect 15754 2096 15788 2130
rect 15824 2096 15858 2130
rect 15894 2096 15928 2130
rect 15964 2096 15998 2130
rect 336 2035 370 2069
rect 405 2035 439 2069
rect 474 2035 508 2069
rect 543 2035 577 2069
rect 612 2035 646 2069
rect 681 2035 715 2069
rect 750 2035 784 2069
rect 819 2035 853 2069
rect 888 2035 922 2069
rect 957 2035 991 2069
rect 1026 2035 1060 2069
rect 1095 2035 1129 2069
rect 1164 2035 1198 2069
rect 1233 2035 1267 2069
rect 1302 2035 1336 2069
rect 1371 2035 1405 2069
rect 1440 2035 1474 2069
rect 1509 2035 1543 2069
rect 1578 2035 1612 2069
rect 1647 2035 1681 2069
rect 1716 2035 1750 2069
rect 1785 2035 1819 2069
rect 1854 2035 1888 2069
rect 1923 2035 1957 2069
rect 1992 2035 2026 2069
rect 2061 2035 2095 2069
rect 2130 2035 2164 2069
rect 2199 2035 2233 2069
rect 2268 2035 2302 2069
rect 2337 2035 2371 2069
rect 2406 2035 2440 2069
rect 2475 2035 2509 2069
rect 2544 2035 2578 2069
rect 2613 2035 2647 2069
rect 2682 2035 2716 2069
rect 2751 2035 2785 2069
rect 2820 2035 2854 2069
rect 2889 2035 2923 2069
rect 2958 2035 2992 2069
rect 3027 2035 3061 2069
rect 3096 2035 3130 2069
rect 3165 2035 3199 2069
rect 3234 2035 3268 2069
rect 3303 2035 3337 2069
rect 3372 2035 3406 2069
rect 3441 2035 3475 2069
rect 3510 2035 3544 2069
rect 3579 2035 3613 2069
rect 3648 2035 3682 2069
rect 3717 2035 3751 2069
rect 3786 2035 3820 2069
rect 3855 2035 3889 2069
rect 3924 2035 3958 2069
rect 3993 2035 4027 2069
rect 4062 2035 4096 2069
rect 4131 2035 4165 2069
rect 4200 2035 4234 2069
rect 4269 2035 4303 2069
rect 4338 2035 4372 2069
rect 4407 2035 4441 2069
rect 4475 2035 4509 2069
rect 4543 2035 4577 2069
rect 4611 2035 4645 2069
rect 4679 2035 4713 2069
rect 4747 2035 4781 2069
rect 4815 2035 4849 2069
rect 4883 2035 4917 2069
rect 4951 2035 4985 2069
rect 5019 2035 5053 2069
rect 5087 2035 5121 2069
rect 5155 2035 5189 2069
rect 5223 2035 5257 2069
rect 5291 2035 5325 2069
rect 5359 2035 5393 2069
rect 5427 2035 5461 2069
rect 5495 2035 5529 2069
rect 5563 2035 5597 2069
rect 5631 2035 5665 2069
rect 5699 2035 5733 2069
rect 5767 2035 5801 2069
rect 5835 2035 5869 2069
rect 5903 2035 5937 2069
rect 5971 2035 6005 2069
rect 6039 2035 6073 2069
rect 6107 2035 6141 2069
rect 6175 2035 6209 2069
rect 6243 2035 6277 2069
rect 6311 2035 6345 2069
rect 6379 2035 6413 2069
rect 6447 2035 6481 2069
rect 6515 2035 6549 2069
rect 6583 2035 6617 2069
rect 6651 2035 6685 2069
rect 6719 2035 6753 2069
rect 6787 2035 6821 2069
rect 6855 2035 6889 2069
rect 6923 2035 6957 2069
rect 6991 2035 7025 2069
rect 7059 2035 7093 2069
rect 7127 2035 7161 2069
rect 7195 2035 7229 2069
rect 7263 2035 7297 2069
rect 7331 2035 7365 2069
rect 7399 2035 7433 2069
rect 7467 2035 7501 2069
rect 7535 2035 7569 2069
rect 7603 2035 7637 2069
rect 7671 2035 7705 2069
rect 7739 2035 7773 2069
rect 7807 2035 7841 2069
rect 7875 2035 7909 2069
rect 7943 2035 7977 2069
rect 8011 2035 8045 2069
rect 8079 2035 8113 2069
rect 8147 2035 8181 2069
rect 8215 2035 8249 2069
rect 8283 2035 8317 2069
rect 8351 2035 8385 2069
rect 8419 2035 8453 2069
rect 8487 2035 8521 2069
rect 8555 2035 8589 2069
rect 8623 2035 8657 2069
rect 8691 2035 8725 2069
rect 8759 2035 8793 2069
rect 8827 2035 8861 2069
rect 8895 2035 8929 2069
rect 8963 2035 8997 2069
rect 9031 2035 9065 2069
rect 9099 2035 9133 2069
rect 9167 2035 9201 2069
rect 9235 2035 9269 2069
rect 9303 2035 9337 2069
rect 9371 2035 9405 2069
rect 9439 2035 9473 2069
rect 9507 2035 9541 2069
rect 9575 2035 9609 2069
rect 9643 2035 9677 2069
rect 9711 2035 9745 2069
rect 9779 2035 9813 2069
rect 9847 2035 9881 2069
rect 9915 2035 9949 2069
rect 9983 2035 10017 2069
rect 10051 2035 10085 2069
rect 10119 2035 10153 2069
rect 10187 2035 10221 2069
rect 10255 2035 10289 2069
rect 10323 2035 10357 2069
rect 10391 2035 10425 2069
rect 10459 2035 10493 2069
rect 10527 2035 10561 2069
rect 10595 2035 10629 2069
rect 10663 2035 10697 2069
rect 10731 2035 10765 2069
rect 10799 2035 10833 2069
rect 10867 2035 10901 2069
rect 10935 2035 10969 2069
rect 11003 2035 11037 2069
rect 11071 2035 11105 2069
rect 11139 2035 11173 2069
rect 11207 2035 11241 2069
rect 11275 2035 11309 2069
rect 11343 2035 11377 2069
rect 11411 2035 11445 2069
rect 11479 2035 11513 2069
rect 11547 2035 11581 2069
rect 11615 2035 11649 2069
rect 11683 2035 11717 2069
rect 11751 2035 11785 2069
rect 11819 2035 11853 2069
rect 11887 2035 11921 2069
rect 11955 2035 11989 2069
rect 12023 2035 12057 2069
rect 12091 2035 12125 2069
rect 12159 2035 12193 2069
rect 12227 2035 12261 2069
rect 12295 2035 12329 2069
rect 12363 2035 12397 2069
rect 12431 2035 12465 2069
rect 12499 2035 12533 2069
rect 12567 2035 12601 2069
rect 12635 2035 12669 2069
rect 12703 2035 12737 2069
rect 12771 2035 12805 2069
rect 12839 2035 12873 2069
rect 12907 2035 12941 2069
rect 12975 2035 13009 2069
rect 13043 2035 13077 2069
rect 13111 2035 13145 2069
rect 13179 2035 13213 2069
rect 13247 2035 13281 2069
rect 13315 2035 13349 2069
rect 13383 2035 13417 2069
rect 13451 2035 13485 2069
rect 13519 2035 13553 2069
rect 13587 2035 13621 2069
rect 13655 2035 13689 2069
rect 13723 2035 13757 2069
rect 13791 2035 13825 2069
rect 13859 2035 13893 2069
rect 13927 2035 13961 2069
rect 13995 2035 14029 2069
rect 14063 2035 14097 2069
rect 14131 2035 14165 2069
rect 14199 2035 14233 2069
rect 14267 2035 14301 2069
rect 14335 2035 14369 2069
rect 14403 2035 14437 2069
rect 14471 2035 14505 2069
rect 14539 2035 14573 2069
rect 14607 2035 14641 2069
rect 14675 2035 14709 2069
rect 14774 2028 14808 2062
rect 14844 2028 14878 2062
rect 14914 2028 14948 2062
rect 14984 2028 15018 2062
rect 15054 2028 15088 2062
rect 15124 2028 15158 2062
rect 15194 2028 15228 2062
rect 15264 2028 15298 2062
rect 15334 2028 15368 2062
rect 15404 2028 15438 2062
rect 15474 2028 15508 2062
rect 15544 2028 15578 2062
rect 15614 2028 15648 2062
rect 15684 2028 15718 2062
rect 15754 2028 15788 2062
rect 15824 2028 15858 2062
rect 15894 2028 15928 2062
rect 15964 2028 15998 2062
rect 360 1925 394 1959
rect 13194 1967 13228 2001
rect 13264 1967 13298 2001
rect 13334 1967 13368 2001
rect 13404 1967 13438 2001
rect 13474 1967 13508 2001
rect 13544 1967 13578 2001
rect 13614 1967 13648 2001
rect 13684 1967 13718 2001
rect 13754 1967 13788 2001
rect 13824 1967 13858 2001
rect 13894 1967 13928 2001
rect 13964 1967 13998 2001
rect 14034 1967 14068 2001
rect 14104 1967 14138 2001
rect 14174 1967 14208 2001
rect 14244 1967 14278 2001
rect 14314 1967 14348 2001
rect 14384 1967 14418 2001
rect 14454 1967 14488 2001
rect 14524 1967 14558 2001
rect 14594 1967 14628 2001
rect 14664 1967 14698 2001
rect 14774 1960 14808 1994
rect 14844 1960 14878 1994
rect 14914 1960 14948 1994
rect 14984 1960 15018 1994
rect 15054 1960 15088 1994
rect 15124 1960 15158 1994
rect 15194 1960 15228 1994
rect 15264 1960 15298 1994
rect 15334 1960 15368 1994
rect 15404 1960 15438 1994
rect 15474 1960 15508 1994
rect 15544 1960 15578 1994
rect 15614 1960 15648 1994
rect 15684 1960 15718 1994
rect 15754 1960 15788 1994
rect 15824 1960 15858 1994
rect 15894 1960 15928 1994
rect 15964 1960 15998 1994
rect 360 1855 394 1889
rect 13194 1897 13228 1931
rect 13264 1897 13298 1931
rect 13334 1897 13368 1931
rect 13404 1897 13438 1931
rect 13474 1897 13508 1931
rect 13544 1897 13578 1931
rect 13614 1897 13648 1931
rect 13684 1897 13718 1931
rect 13754 1897 13788 1931
rect 13824 1897 13858 1931
rect 13894 1897 13928 1931
rect 13964 1897 13998 1931
rect 14034 1897 14068 1931
rect 14104 1897 14138 1931
rect 14174 1897 14208 1931
rect 14244 1897 14278 1931
rect 14314 1897 14348 1931
rect 14384 1897 14418 1931
rect 14454 1897 14488 1931
rect 14524 1897 14558 1931
rect 14594 1897 14628 1931
rect 14664 1897 14698 1931
rect 14774 1892 14808 1926
rect 14844 1892 14878 1926
rect 14914 1892 14948 1926
rect 14984 1892 15018 1926
rect 15054 1892 15088 1926
rect 15124 1892 15158 1926
rect 15194 1892 15228 1926
rect 15264 1892 15298 1926
rect 15334 1892 15368 1926
rect 15404 1892 15438 1926
rect 15474 1892 15508 1926
rect 15544 1892 15578 1926
rect 15614 1892 15648 1926
rect 15684 1892 15718 1926
rect 15754 1892 15788 1926
rect 15824 1892 15858 1926
rect 15894 1892 15928 1926
rect 15964 1892 15998 1926
rect 360 1785 394 1819
rect 13194 1827 13228 1861
rect 13264 1827 13298 1861
rect 13334 1827 13368 1861
rect 13404 1827 13438 1861
rect 13474 1827 13508 1861
rect 13544 1827 13578 1861
rect 13614 1827 13648 1861
rect 13684 1827 13718 1861
rect 13754 1827 13788 1861
rect 13824 1827 13858 1861
rect 13894 1827 13928 1861
rect 13964 1827 13998 1861
rect 14034 1827 14068 1861
rect 14104 1827 14138 1861
rect 14174 1827 14208 1861
rect 14244 1827 14278 1861
rect 14314 1827 14348 1861
rect 14384 1827 14418 1861
rect 14454 1827 14488 1861
rect 14524 1827 14558 1861
rect 14594 1827 14628 1861
rect 14664 1827 14698 1861
rect 14774 1824 14808 1858
rect 14844 1824 14878 1858
rect 14914 1824 14948 1858
rect 14984 1824 15018 1858
rect 15054 1824 15088 1858
rect 15124 1824 15158 1858
rect 15194 1824 15228 1858
rect 15264 1824 15298 1858
rect 15334 1824 15368 1858
rect 15404 1824 15438 1858
rect 15474 1824 15508 1858
rect 15544 1824 15578 1858
rect 15614 1824 15648 1858
rect 15684 1824 15718 1858
rect 15754 1824 15788 1858
rect 15824 1824 15858 1858
rect 15894 1824 15928 1858
rect 15964 1824 15998 1858
rect 360 1715 394 1749
rect 13194 1757 13228 1791
rect 13264 1757 13298 1791
rect 13334 1757 13368 1791
rect 13404 1757 13438 1791
rect 13474 1757 13508 1791
rect 13544 1757 13578 1791
rect 13614 1757 13648 1791
rect 13684 1757 13718 1791
rect 13754 1757 13788 1791
rect 13824 1757 13858 1791
rect 13894 1757 13928 1791
rect 13964 1757 13998 1791
rect 14034 1757 14068 1791
rect 14104 1757 14138 1791
rect 14174 1757 14208 1791
rect 14244 1757 14278 1791
rect 14314 1757 14348 1791
rect 14384 1757 14418 1791
rect 14454 1757 14488 1791
rect 14524 1757 14558 1791
rect 14594 1757 14628 1791
rect 14664 1757 14698 1791
rect 14774 1756 14808 1790
rect 14844 1756 14878 1790
rect 14914 1756 14948 1790
rect 14984 1756 15018 1790
rect 15054 1756 15088 1790
rect 15124 1756 15158 1790
rect 15194 1756 15228 1790
rect 15264 1756 15298 1790
rect 15334 1756 15368 1790
rect 15404 1756 15438 1790
rect 15474 1756 15508 1790
rect 15544 1756 15578 1790
rect 15614 1756 15648 1790
rect 15684 1756 15718 1790
rect 15754 1756 15788 1790
rect 15824 1756 15858 1790
rect 15894 1756 15928 1790
rect 15964 1756 15998 1790
rect 360 1645 394 1679
rect 13194 1687 13228 1721
rect 13264 1687 13298 1721
rect 13334 1687 13368 1721
rect 13404 1687 13438 1721
rect 13474 1687 13508 1721
rect 13544 1687 13578 1721
rect 13614 1687 13648 1721
rect 13684 1687 13718 1721
rect 13754 1687 13788 1721
rect 13824 1687 13858 1721
rect 13894 1687 13928 1721
rect 13964 1687 13998 1721
rect 14034 1687 14068 1721
rect 14104 1687 14138 1721
rect 14174 1687 14208 1721
rect 14244 1687 14278 1721
rect 14314 1687 14348 1721
rect 14384 1687 14418 1721
rect 14454 1687 14488 1721
rect 14524 1687 14558 1721
rect 14594 1687 14628 1721
rect 14664 1687 14698 1721
rect 14774 1688 14808 1722
rect 14844 1688 14878 1722
rect 14914 1688 14948 1722
rect 14984 1688 15018 1722
rect 15054 1688 15088 1722
rect 15124 1688 15158 1722
rect 15194 1688 15228 1722
rect 15264 1688 15298 1722
rect 15334 1688 15368 1722
rect 15404 1688 15438 1722
rect 15474 1688 15508 1722
rect 15544 1688 15578 1722
rect 15614 1688 15648 1722
rect 15684 1688 15718 1722
rect 15754 1688 15788 1722
rect 15824 1688 15858 1722
rect 15894 1688 15928 1722
rect 15964 1688 15998 1722
rect 360 1575 394 1609
rect 13194 1617 13228 1651
rect 13264 1617 13298 1651
rect 13334 1617 13368 1651
rect 13404 1617 13438 1651
rect 13474 1617 13508 1651
rect 13544 1617 13578 1651
rect 13614 1617 13648 1651
rect 13684 1617 13718 1651
rect 13754 1617 13788 1651
rect 13824 1617 13858 1651
rect 13894 1617 13928 1651
rect 13964 1617 13998 1651
rect 14034 1617 14068 1651
rect 14104 1617 14138 1651
rect 14174 1617 14208 1651
rect 14244 1617 14278 1651
rect 14314 1617 14348 1651
rect 14384 1617 14418 1651
rect 14454 1617 14488 1651
rect 14524 1617 14558 1651
rect 14594 1617 14628 1651
rect 14664 1617 14698 1651
rect 14774 1620 14808 1654
rect 14844 1620 14878 1654
rect 14914 1620 14948 1654
rect 14984 1620 15018 1654
rect 15054 1620 15088 1654
rect 15124 1620 15158 1654
rect 15194 1620 15228 1654
rect 15264 1620 15298 1654
rect 15334 1620 15368 1654
rect 15404 1620 15438 1654
rect 15474 1620 15508 1654
rect 15544 1620 15578 1654
rect 15614 1620 15648 1654
rect 15684 1620 15718 1654
rect 15754 1620 15788 1654
rect 15824 1620 15858 1654
rect 15894 1620 15928 1654
rect 15964 1620 15998 1654
rect 360 1505 394 1539
rect 13194 1547 13228 1581
rect 13264 1547 13298 1581
rect 13334 1547 13368 1581
rect 13404 1547 13438 1581
rect 13474 1547 13508 1581
rect 13544 1547 13578 1581
rect 13614 1547 13648 1581
rect 13684 1547 13718 1581
rect 13754 1547 13788 1581
rect 13824 1547 13858 1581
rect 13894 1547 13928 1581
rect 13964 1547 13998 1581
rect 14034 1547 14068 1581
rect 14104 1547 14138 1581
rect 14174 1547 14208 1581
rect 14244 1547 14278 1581
rect 14314 1547 14348 1581
rect 14384 1547 14418 1581
rect 14454 1547 14488 1581
rect 14524 1547 14558 1581
rect 14594 1547 14628 1581
rect 14664 1547 14698 1581
rect 14774 1552 14808 1586
rect 14844 1552 14878 1586
rect 14914 1552 14948 1586
rect 14984 1552 15018 1586
rect 15054 1552 15088 1586
rect 15124 1552 15158 1586
rect 15194 1552 15228 1586
rect 15264 1552 15298 1586
rect 15334 1552 15368 1586
rect 15404 1552 15438 1586
rect 15474 1552 15508 1586
rect 15544 1552 15578 1586
rect 15614 1552 15648 1586
rect 15684 1552 15718 1586
rect 15754 1552 15788 1586
rect 15824 1552 15858 1586
rect 15894 1552 15928 1586
rect 15964 1552 15998 1586
rect 360 1435 394 1469
rect 360 1365 394 1399
rect 13194 1477 13228 1511
rect 13264 1477 13298 1511
rect 13334 1477 13368 1511
rect 13404 1477 13438 1511
rect 13474 1477 13508 1511
rect 13544 1477 13578 1511
rect 13614 1477 13648 1511
rect 13684 1477 13718 1511
rect 13754 1477 13788 1511
rect 13824 1477 13858 1511
rect 13894 1477 13928 1511
rect 13964 1477 13998 1511
rect 14034 1477 14068 1511
rect 14104 1477 14138 1511
rect 14174 1477 14208 1511
rect 14244 1477 14278 1511
rect 14314 1477 14348 1511
rect 14384 1477 14418 1511
rect 14454 1477 14488 1511
rect 14524 1477 14558 1511
rect 14594 1477 14628 1511
rect 14664 1477 14698 1511
rect 14774 1484 14808 1518
rect 14844 1484 14878 1518
rect 14914 1484 14948 1518
rect 14984 1484 15018 1518
rect 15054 1484 15088 1518
rect 15124 1484 15158 1518
rect 15194 1484 15228 1518
rect 15264 1484 15298 1518
rect 15334 1484 15368 1518
rect 15404 1484 15438 1518
rect 15474 1484 15508 1518
rect 15544 1484 15578 1518
rect 15614 1484 15648 1518
rect 15684 1484 15718 1518
rect 15754 1484 15788 1518
rect 15824 1484 15858 1518
rect 15894 1484 15928 1518
rect 15964 1484 15998 1518
rect 13194 1407 13228 1441
rect 13264 1407 13298 1441
rect 13334 1407 13368 1441
rect 13404 1407 13438 1441
rect 13474 1407 13508 1441
rect 13544 1407 13578 1441
rect 13614 1407 13648 1441
rect 13684 1407 13718 1441
rect 13754 1407 13788 1441
rect 13824 1407 13858 1441
rect 13894 1407 13928 1441
rect 13964 1407 13998 1441
rect 14034 1407 14068 1441
rect 14104 1407 14138 1441
rect 14174 1407 14208 1441
rect 14244 1407 14278 1441
rect 14314 1407 14348 1441
rect 14384 1407 14418 1441
rect 14454 1407 14488 1441
rect 14524 1407 14558 1441
rect 14594 1407 14628 1441
rect 14664 1407 14698 1441
rect 14774 1416 14808 1450
rect 14844 1416 14878 1450
rect 14914 1416 14948 1450
rect 14984 1416 15018 1450
rect 15054 1416 15088 1450
rect 15124 1416 15158 1450
rect 15194 1416 15228 1450
rect 15264 1416 15298 1450
rect 15334 1416 15368 1450
rect 15404 1416 15438 1450
rect 15474 1416 15508 1450
rect 15544 1416 15578 1450
rect 15614 1416 15648 1450
rect 15684 1416 15718 1450
rect 15754 1416 15788 1450
rect 15824 1416 15858 1450
rect 15894 1416 15928 1450
rect 15964 1416 15998 1450
rect 360 1295 394 1329
rect 360 1225 394 1259
rect 13194 1337 13228 1371
rect 13264 1337 13298 1371
rect 13334 1337 13368 1371
rect 13404 1337 13438 1371
rect 13474 1337 13508 1371
rect 13544 1337 13578 1371
rect 13614 1337 13648 1371
rect 13684 1337 13718 1371
rect 13754 1337 13788 1371
rect 13824 1337 13858 1371
rect 13894 1337 13928 1371
rect 13964 1337 13998 1371
rect 14034 1337 14068 1371
rect 14104 1337 14138 1371
rect 14174 1337 14208 1371
rect 14244 1337 14278 1371
rect 14314 1337 14348 1371
rect 14384 1337 14418 1371
rect 14454 1337 14488 1371
rect 14524 1337 14558 1371
rect 14594 1337 14628 1371
rect 14664 1337 14698 1371
rect 14774 1348 14808 1382
rect 14844 1348 14878 1382
rect 14914 1348 14948 1382
rect 14984 1348 15018 1382
rect 15054 1348 15088 1382
rect 15124 1348 15158 1382
rect 15194 1348 15228 1382
rect 15264 1348 15298 1382
rect 15334 1348 15368 1382
rect 15404 1348 15438 1382
rect 15474 1348 15508 1382
rect 15544 1348 15578 1382
rect 15614 1348 15648 1382
rect 15684 1348 15718 1382
rect 15754 1348 15788 1382
rect 15824 1348 15858 1382
rect 15894 1348 15928 1382
rect 15964 1348 15998 1382
rect 13194 1267 13228 1301
rect 13264 1267 13298 1301
rect 13334 1267 13368 1301
rect 13404 1267 13438 1301
rect 13474 1267 13508 1301
rect 13544 1267 13578 1301
rect 13614 1267 13648 1301
rect 13684 1267 13718 1301
rect 13754 1267 13788 1301
rect 13824 1267 13858 1301
rect 13894 1267 13928 1301
rect 13964 1267 13998 1301
rect 14034 1267 14068 1301
rect 14104 1267 14138 1301
rect 14174 1267 14208 1301
rect 14244 1267 14278 1301
rect 14314 1267 14348 1301
rect 14384 1267 14418 1301
rect 14454 1267 14488 1301
rect 14524 1267 14558 1301
rect 14594 1267 14628 1301
rect 14664 1267 14698 1301
rect 14774 1280 14808 1314
rect 14844 1280 14878 1314
rect 14914 1280 14948 1314
rect 14984 1280 15018 1314
rect 15054 1280 15088 1314
rect 15124 1280 15158 1314
rect 15194 1280 15228 1314
rect 15264 1280 15298 1314
rect 15334 1280 15368 1314
rect 15404 1280 15438 1314
rect 15474 1280 15508 1314
rect 15544 1280 15578 1314
rect 15614 1280 15648 1314
rect 15684 1280 15718 1314
rect 15754 1280 15788 1314
rect 15824 1280 15858 1314
rect 15894 1280 15928 1314
rect 15964 1280 15998 1314
rect 360 1155 394 1189
rect 13194 1197 13228 1231
rect 13264 1197 13298 1231
rect 13334 1197 13368 1231
rect 13404 1197 13438 1231
rect 13474 1197 13508 1231
rect 13544 1197 13578 1231
rect 13614 1197 13648 1231
rect 13684 1197 13718 1231
rect 13754 1197 13788 1231
rect 13824 1197 13858 1231
rect 13894 1197 13928 1231
rect 13964 1197 13998 1231
rect 14034 1197 14068 1231
rect 14104 1197 14138 1231
rect 14174 1197 14208 1231
rect 14244 1197 14278 1231
rect 14314 1197 14348 1231
rect 14384 1197 14418 1231
rect 14454 1197 14488 1231
rect 14524 1197 14558 1231
rect 14594 1197 14628 1231
rect 14664 1197 14698 1231
rect 14774 1212 14808 1246
rect 14844 1212 14878 1246
rect 14914 1212 14948 1246
rect 14984 1212 15018 1246
rect 15054 1212 15088 1246
rect 15124 1212 15158 1246
rect 15194 1212 15228 1246
rect 15264 1212 15298 1246
rect 15334 1212 15368 1246
rect 15404 1212 15438 1246
rect 15474 1212 15508 1246
rect 15544 1212 15578 1246
rect 15614 1212 15648 1246
rect 15684 1212 15718 1246
rect 15754 1212 15788 1246
rect 15824 1212 15858 1246
rect 15894 1212 15928 1246
rect 15964 1212 15998 1246
rect 360 1085 394 1119
rect 13194 1127 13228 1161
rect 13264 1127 13298 1161
rect 13334 1127 13368 1161
rect 13404 1127 13438 1161
rect 13474 1127 13508 1161
rect 13544 1127 13578 1161
rect 13614 1127 13648 1161
rect 13684 1127 13718 1161
rect 13754 1127 13788 1161
rect 13824 1127 13858 1161
rect 13894 1127 13928 1161
rect 13964 1127 13998 1161
rect 14034 1127 14068 1161
rect 14104 1127 14138 1161
rect 14174 1127 14208 1161
rect 14244 1127 14278 1161
rect 14314 1127 14348 1161
rect 14384 1127 14418 1161
rect 14454 1127 14488 1161
rect 14524 1127 14558 1161
rect 14594 1127 14628 1161
rect 14664 1127 14698 1161
rect 14774 1144 14808 1178
rect 14844 1144 14878 1178
rect 14914 1144 14948 1178
rect 14984 1144 15018 1178
rect 15054 1144 15088 1178
rect 15124 1144 15158 1178
rect 15194 1144 15228 1178
rect 15264 1144 15298 1178
rect 15334 1144 15368 1178
rect 15404 1144 15438 1178
rect 15474 1144 15508 1178
rect 15544 1144 15578 1178
rect 15614 1144 15648 1178
rect 15684 1144 15718 1178
rect 15754 1144 15788 1178
rect 15824 1144 15858 1178
rect 15894 1144 15928 1178
rect 15964 1144 15998 1178
rect 360 1016 394 1050
rect 13194 1057 13228 1091
rect 13264 1057 13298 1091
rect 13334 1057 13368 1091
rect 13404 1057 13438 1091
rect 13474 1057 13508 1091
rect 13544 1057 13578 1091
rect 13614 1057 13648 1091
rect 13684 1057 13718 1091
rect 13754 1057 13788 1091
rect 13824 1057 13858 1091
rect 13894 1057 13928 1091
rect 13964 1057 13998 1091
rect 14034 1057 14068 1091
rect 14104 1057 14138 1091
rect 14174 1057 14208 1091
rect 14244 1057 14278 1091
rect 14314 1057 14348 1091
rect 14384 1057 14418 1091
rect 14454 1057 14488 1091
rect 14524 1057 14558 1091
rect 14594 1057 14628 1091
rect 14664 1057 14698 1091
rect 14774 1076 14808 1110
rect 14844 1076 14878 1110
rect 14914 1076 14948 1110
rect 14984 1076 15018 1110
rect 15054 1076 15088 1110
rect 15124 1076 15158 1110
rect 15194 1076 15228 1110
rect 15264 1076 15298 1110
rect 15334 1076 15368 1110
rect 15404 1076 15438 1110
rect 15474 1076 15508 1110
rect 15544 1076 15578 1110
rect 15614 1076 15648 1110
rect 15684 1076 15718 1110
rect 15754 1076 15788 1110
rect 15824 1076 15858 1110
rect 15894 1076 15928 1110
rect 15964 1076 15998 1110
rect 360 947 394 981
rect 13194 987 13228 1021
rect 13264 987 13298 1021
rect 13334 987 13368 1021
rect 13404 987 13438 1021
rect 13474 987 13508 1021
rect 13544 987 13578 1021
rect 13614 987 13648 1021
rect 13684 987 13718 1021
rect 13754 987 13788 1021
rect 13824 987 13858 1021
rect 13894 987 13928 1021
rect 13964 987 13998 1021
rect 14034 987 14068 1021
rect 14104 987 14138 1021
rect 14174 987 14208 1021
rect 14244 987 14278 1021
rect 14314 987 14348 1021
rect 14384 987 14418 1021
rect 14454 987 14488 1021
rect 14524 987 14558 1021
rect 14594 987 14628 1021
rect 14664 987 14698 1021
rect 14774 1008 14808 1042
rect 14844 1008 14878 1042
rect 14914 1008 14948 1042
rect 14984 1008 15018 1042
rect 15054 1008 15088 1042
rect 15124 1008 15158 1042
rect 15194 1008 15228 1042
rect 15264 1008 15298 1042
rect 15334 1008 15368 1042
rect 15404 1008 15438 1042
rect 15474 1008 15508 1042
rect 15544 1008 15578 1042
rect 15614 1008 15648 1042
rect 15684 1008 15718 1042
rect 15754 1008 15788 1042
rect 15824 1008 15858 1042
rect 15894 1008 15928 1042
rect 15964 1008 15998 1042
rect 360 878 394 912
rect 13194 917 13228 951
rect 13264 917 13298 951
rect 13334 917 13368 951
rect 13404 917 13438 951
rect 13474 917 13508 951
rect 13544 917 13578 951
rect 13614 917 13648 951
rect 13684 917 13718 951
rect 13754 917 13788 951
rect 13824 917 13858 951
rect 13894 917 13928 951
rect 13964 917 13998 951
rect 14034 917 14068 951
rect 14104 917 14138 951
rect 14174 917 14208 951
rect 14244 917 14278 951
rect 14314 917 14348 951
rect 14384 917 14418 951
rect 14454 917 14488 951
rect 14524 917 14558 951
rect 14594 917 14628 951
rect 14664 917 14698 951
rect 14774 940 14808 974
rect 14844 940 14878 974
rect 14914 940 14948 974
rect 14984 940 15018 974
rect 15054 940 15088 974
rect 15124 940 15158 974
rect 15194 940 15228 974
rect 15264 940 15298 974
rect 15334 940 15368 974
rect 15404 940 15438 974
rect 15474 940 15508 974
rect 15544 940 15578 974
rect 15614 940 15648 974
rect 15684 940 15718 974
rect 15754 940 15788 974
rect 15824 940 15858 974
rect 15894 940 15928 974
rect 15964 940 15998 974
rect 360 809 394 843
rect 13194 847 13228 881
rect 13264 847 13298 881
rect 13334 847 13368 881
rect 13404 847 13438 881
rect 13474 847 13508 881
rect 13544 847 13578 881
rect 13614 847 13648 881
rect 13684 847 13718 881
rect 13754 847 13788 881
rect 13824 847 13858 881
rect 13894 847 13928 881
rect 13964 847 13998 881
rect 14034 847 14068 881
rect 14104 847 14138 881
rect 14174 847 14208 881
rect 14244 847 14278 881
rect 14314 847 14348 881
rect 14384 847 14418 881
rect 14454 847 14488 881
rect 14524 847 14558 881
rect 14594 847 14628 881
rect 14664 847 14698 881
rect 14774 872 14808 906
rect 14844 872 14878 906
rect 14914 872 14948 906
rect 14984 872 15018 906
rect 15054 872 15088 906
rect 15124 872 15158 906
rect 15194 872 15228 906
rect 15264 872 15298 906
rect 15334 872 15368 906
rect 15404 872 15438 906
rect 15474 872 15508 906
rect 15544 872 15578 906
rect 15614 872 15648 906
rect 15684 872 15718 906
rect 15754 872 15788 906
rect 15824 872 15858 906
rect 15894 872 15928 906
rect 15964 872 15998 906
rect 360 740 394 774
rect 13194 777 13228 811
rect 13264 777 13298 811
rect 13334 777 13368 811
rect 13404 777 13438 811
rect 13474 777 13508 811
rect 13544 777 13578 811
rect 13614 777 13648 811
rect 13684 777 13718 811
rect 13754 777 13788 811
rect 13824 777 13858 811
rect 13894 777 13928 811
rect 13964 777 13998 811
rect 14034 777 14068 811
rect 14104 777 14138 811
rect 14174 777 14208 811
rect 14244 777 14278 811
rect 14314 777 14348 811
rect 14384 777 14418 811
rect 14454 777 14488 811
rect 14524 777 14558 811
rect 14594 777 14628 811
rect 14664 777 14698 811
rect 14774 804 14808 838
rect 14844 804 14878 838
rect 14914 804 14948 838
rect 14984 804 15018 838
rect 15054 804 15088 838
rect 15124 804 15158 838
rect 15194 804 15228 838
rect 15264 804 15298 838
rect 15334 804 15368 838
rect 15404 804 15438 838
rect 15474 804 15508 838
rect 15544 804 15578 838
rect 15614 804 15648 838
rect 15684 804 15718 838
rect 15754 804 15788 838
rect 15824 804 15858 838
rect 15894 804 15928 838
rect 15964 804 15998 838
rect 360 671 394 705
rect 360 602 394 636
rect 13194 707 13228 741
rect 13264 707 13298 741
rect 13334 707 13368 741
rect 13404 707 13438 741
rect 13474 707 13508 741
rect 13544 707 13578 741
rect 13614 707 13648 741
rect 13684 707 13718 741
rect 13754 707 13788 741
rect 13824 707 13858 741
rect 13894 707 13928 741
rect 13964 707 13998 741
rect 14034 707 14068 741
rect 14104 707 14138 741
rect 14174 707 14208 741
rect 14244 707 14278 741
rect 14314 707 14348 741
rect 14384 707 14418 741
rect 14454 707 14488 741
rect 14524 707 14558 741
rect 14594 707 14628 741
rect 14664 707 14698 741
rect 14774 736 14808 770
rect 14844 736 14878 770
rect 14914 736 14948 770
rect 14984 736 15018 770
rect 15054 736 15088 770
rect 15124 736 15158 770
rect 15194 736 15228 770
rect 15264 736 15298 770
rect 15334 736 15368 770
rect 15404 736 15438 770
rect 15474 736 15508 770
rect 15544 736 15578 770
rect 15614 736 15648 770
rect 15684 736 15718 770
rect 15754 736 15788 770
rect 15824 736 15858 770
rect 15894 736 15928 770
rect 15964 736 15998 770
rect 13194 637 13228 671
rect 13264 637 13298 671
rect 13334 637 13368 671
rect 13404 637 13438 671
rect 13474 637 13508 671
rect 13544 637 13578 671
rect 13614 637 13648 671
rect 13684 637 13718 671
rect 13754 637 13788 671
rect 13824 637 13858 671
rect 13894 637 13928 671
rect 13964 637 13998 671
rect 14034 637 14068 671
rect 14104 637 14138 671
rect 14174 637 14208 671
rect 14244 637 14278 671
rect 14314 637 14348 671
rect 14384 637 14418 671
rect 14454 637 14488 671
rect 14524 637 14558 671
rect 14594 637 14628 671
rect 14664 637 14698 671
rect 14774 668 14808 702
rect 14844 668 14878 702
rect 14914 668 14948 702
rect 14984 668 15018 702
rect 15054 668 15088 702
rect 15124 668 15158 702
rect 15194 668 15228 702
rect 15264 668 15298 702
rect 15334 668 15368 702
rect 15404 668 15438 702
rect 15474 668 15508 702
rect 15544 668 15578 702
rect 15614 668 15648 702
rect 15684 668 15718 702
rect 15754 668 15788 702
rect 15824 668 15858 702
rect 15894 668 15928 702
rect 15964 668 15998 702
rect 360 533 394 567
rect 360 464 394 498
rect 13194 567 13228 601
rect 13264 567 13298 601
rect 13334 567 13368 601
rect 13404 567 13438 601
rect 13474 567 13508 601
rect 13544 567 13578 601
rect 13614 567 13648 601
rect 13684 567 13718 601
rect 13754 567 13788 601
rect 13824 567 13858 601
rect 13894 567 13928 601
rect 13964 567 13998 601
rect 14034 567 14068 601
rect 14104 567 14138 601
rect 14174 567 14208 601
rect 14244 567 14278 601
rect 14314 567 14348 601
rect 14384 567 14418 601
rect 14454 567 14488 601
rect 14524 567 14558 601
rect 14594 567 14628 601
rect 14664 567 14698 601
rect 14774 600 14808 634
rect 14844 600 14878 634
rect 14914 600 14948 634
rect 14984 600 15018 634
rect 15054 600 15088 634
rect 15124 600 15158 634
rect 15194 600 15228 634
rect 15264 600 15298 634
rect 15334 600 15368 634
rect 15404 600 15438 634
rect 15474 600 15508 634
rect 15544 600 15578 634
rect 15614 600 15648 634
rect 15684 600 15718 634
rect 15754 600 15788 634
rect 15824 600 15858 634
rect 15894 600 15928 634
rect 15964 600 15998 634
rect 14774 532 14808 566
rect 14844 532 14878 566
rect 14914 532 14948 566
rect 14984 532 15018 566
rect 15054 532 15088 566
rect 15124 532 15158 566
rect 15194 532 15228 566
rect 15264 532 15298 566
rect 15334 532 15368 566
rect 15404 532 15438 566
rect 15474 532 15508 566
rect 15544 532 15578 566
rect 15614 532 15648 566
rect 15684 532 15718 566
rect 15754 532 15788 566
rect 15824 532 15858 566
rect 15894 532 15928 566
rect 15964 532 15998 566
rect 13194 497 13228 531
rect 13264 497 13298 531
rect 13334 497 13368 531
rect 13404 497 13438 531
rect 13474 497 13508 531
rect 13544 497 13578 531
rect 13614 497 13648 531
rect 13684 497 13718 531
rect 13754 497 13788 531
rect 13824 497 13858 531
rect 13894 497 13928 531
rect 13964 497 13998 531
rect 14034 497 14068 531
rect 14104 497 14138 531
rect 14174 497 14208 531
rect 14244 497 14278 531
rect 14314 497 14348 531
rect 14384 497 14418 531
rect 14454 497 14488 531
rect 14524 497 14558 531
rect 14594 497 14628 531
rect 14664 497 14698 531
rect 360 395 394 429
rect 14774 464 14808 498
rect 14844 464 14878 498
rect 14914 464 14948 498
rect 14984 464 15018 498
rect 15054 464 15088 498
rect 15124 464 15158 498
rect 15194 464 15228 498
rect 15264 464 15298 498
rect 15334 464 15368 498
rect 15404 464 15438 498
rect 15474 464 15508 498
rect 15544 464 15578 498
rect 15614 464 15648 498
rect 15684 464 15718 498
rect 15754 464 15788 498
rect 15824 464 15858 498
rect 15894 464 15928 498
rect 15964 464 15998 498
rect 13194 427 13228 461
rect 13264 427 13298 461
rect 13334 427 13368 461
rect 13404 427 13438 461
rect 13474 427 13508 461
rect 13544 427 13578 461
rect 13614 427 13648 461
rect 13684 427 13718 461
rect 13754 427 13788 461
rect 13824 427 13858 461
rect 13894 427 13928 461
rect 13964 427 13998 461
rect 14034 427 14068 461
rect 14104 427 14138 461
rect 14174 427 14208 461
rect 14244 427 14278 461
rect 14314 427 14348 461
rect 14384 427 14418 461
rect 14454 427 14488 461
rect 14524 427 14558 461
rect 14594 427 14628 461
rect 14664 427 14698 461
rect 360 326 394 360
rect 14774 396 14808 430
rect 14844 396 14878 430
rect 14914 396 14948 430
rect 14984 396 15018 430
rect 15054 396 15088 430
rect 15124 396 15158 430
rect 15194 396 15228 430
rect 15264 396 15298 430
rect 15334 396 15368 430
rect 15404 396 15438 430
rect 15474 396 15508 430
rect 15544 396 15578 430
rect 15614 396 15648 430
rect 15684 396 15718 430
rect 15754 396 15788 430
rect 15824 396 15858 430
rect 15894 396 15928 430
rect 15964 396 15998 430
rect 13194 357 13228 391
rect 13264 357 13298 391
rect 13334 357 13368 391
rect 13404 357 13438 391
rect 13474 357 13508 391
rect 13544 357 13578 391
rect 13614 357 13648 391
rect 13684 357 13718 391
rect 13754 357 13788 391
rect 13824 357 13858 391
rect 13894 357 13928 391
rect 13964 357 13998 391
rect 14034 357 14068 391
rect 14104 357 14138 391
rect 14174 357 14208 391
rect 14244 357 14278 391
rect 14314 357 14348 391
rect 14384 357 14418 391
rect 14454 357 14488 391
rect 14524 357 14558 391
rect 14594 357 14628 391
rect 14664 357 14698 391
rect 14774 328 14808 362
rect 14844 328 14878 362
rect 14914 328 14948 362
rect 14984 328 15018 362
rect 15054 328 15088 362
rect 15124 328 15158 362
rect 15194 328 15228 362
rect 15264 328 15298 362
rect 15334 328 15368 362
rect 15404 328 15438 362
rect 15474 328 15508 362
rect 15544 328 15578 362
rect 15614 328 15648 362
rect 15684 328 15718 362
rect 15754 328 15788 362
rect 15824 328 15858 362
rect 15894 328 15928 362
rect 15964 328 15998 362
rect 360 257 394 291
rect 13194 287 13228 321
rect 13264 287 13298 321
rect 13334 287 13368 321
rect 13404 287 13438 321
rect 13474 287 13508 321
rect 13544 287 13578 321
rect 13614 287 13648 321
rect 13684 287 13718 321
rect 13754 287 13788 321
rect 13824 287 13858 321
rect 13894 287 13928 321
rect 13964 287 13998 321
rect 14034 287 14068 321
rect 14104 287 14138 321
rect 14174 287 14208 321
rect 14244 287 14278 321
rect 14314 287 14348 321
rect 14384 287 14418 321
rect 14454 287 14488 321
rect 14524 287 14558 321
rect 14594 287 14628 321
rect 14664 287 14698 321
rect 360 188 394 222
rect 14774 260 14808 294
rect 14844 260 14878 294
rect 14914 260 14948 294
rect 14984 260 15018 294
rect 15054 260 15088 294
rect 15124 260 15158 294
rect 15194 260 15228 294
rect 15264 260 15298 294
rect 15334 260 15368 294
rect 15404 260 15438 294
rect 15474 260 15508 294
rect 15544 260 15578 294
rect 15614 260 15648 294
rect 15684 260 15718 294
rect 15754 260 15788 294
rect 15824 260 15858 294
rect 15894 260 15928 294
rect 15964 260 15998 294
rect 13194 217 13228 251
rect 13264 217 13298 251
rect 13334 217 13368 251
rect 13404 217 13438 251
rect 13474 217 13508 251
rect 13544 217 13578 251
rect 13614 217 13648 251
rect 13684 217 13718 251
rect 13754 217 13788 251
rect 13824 217 13858 251
rect 13894 217 13928 251
rect 13964 217 13998 251
rect 14034 217 14068 251
rect 14104 217 14138 251
rect 14174 217 14208 251
rect 14244 217 14278 251
rect 14314 217 14348 251
rect 14384 217 14418 251
rect 14454 217 14488 251
rect 14524 217 14558 251
rect 14594 217 14628 251
rect 14664 217 14698 251
rect 14774 192 14808 226
rect 14844 192 14878 226
rect 14914 192 14948 226
rect 14984 192 15018 226
rect 15054 192 15088 226
rect 15124 192 15158 226
rect 15194 192 15228 226
rect 15264 192 15298 226
rect 15334 192 15368 226
rect 15404 192 15438 226
rect 15474 192 15508 226
rect 15544 192 15578 226
rect 15614 192 15648 226
rect 15684 192 15718 226
rect 15754 192 15788 226
rect 15824 192 15858 226
rect 15894 192 15928 226
rect 15964 192 15998 226
rect 360 119 394 153
rect 13194 147 13228 181
rect 13264 147 13298 181
rect 13334 147 13368 181
rect 13404 147 13438 181
rect 13474 147 13508 181
rect 13544 147 13578 181
rect 13614 147 13648 181
rect 13684 147 13718 181
rect 13754 147 13788 181
rect 13824 147 13858 181
rect 13894 147 13928 181
rect 13964 147 13998 181
rect 14034 147 14068 181
rect 14104 147 14138 181
rect 14174 147 14208 181
rect 14244 147 14278 181
rect 14314 147 14348 181
rect 14384 147 14418 181
rect 14454 147 14488 181
rect 14524 147 14558 181
rect 14594 147 14628 181
rect 14664 147 14698 181
rect 14774 124 14808 158
rect 14844 124 14878 158
rect 14914 124 14948 158
rect 14984 124 15018 158
rect 15054 124 15088 158
rect 15124 124 15158 158
rect 15194 124 15228 158
rect 15264 124 15298 158
rect 15334 124 15368 158
rect 15404 124 15438 158
rect 15474 124 15508 158
rect 15544 124 15578 158
rect 15614 124 15648 158
rect 15684 124 15718 158
rect 15754 124 15788 158
rect 15824 124 15858 158
rect 15894 124 15928 158
rect 15964 124 15998 158
rect 360 50 394 84
rect 429 50 463 84
rect 498 50 532 84
rect 567 50 601 84
rect 636 50 670 84
rect 705 50 739 84
rect 774 50 808 84
rect 843 50 877 84
rect 912 50 946 84
rect 981 50 1015 84
rect 1050 50 1084 84
rect 1119 50 1153 84
rect 1188 50 1222 84
rect 1257 50 1291 84
rect 1326 50 1360 84
rect 1395 50 1429 84
rect 1464 50 1498 84
rect 1533 50 1567 84
rect 1602 50 1636 84
rect 1671 50 1705 84
rect 1740 50 1774 84
rect 1809 50 1843 84
rect 1878 50 1912 84
rect 1947 50 1981 84
rect 2016 50 2050 84
rect 2085 50 2119 84
rect 2154 50 2188 84
rect 2223 50 2257 84
rect 2292 50 2326 84
rect 2361 50 2395 84
rect 2430 50 2464 84
rect 2499 50 2533 84
rect 2568 50 2602 84
rect 2637 50 2671 84
rect 2706 50 2740 84
rect 2775 50 2809 84
rect 2844 50 2878 84
rect 2913 50 2947 84
rect 2982 50 3016 84
rect 3051 50 3085 84
rect 3120 50 3154 84
rect 3189 50 3223 84
rect 3258 50 3292 84
rect 3327 50 3361 84
rect 3396 50 3430 84
rect 3465 50 3499 84
rect 3534 50 3568 84
rect 3603 50 3637 84
rect 3672 50 3706 84
rect 3741 50 3775 84
rect 3810 50 3844 84
rect 3879 50 3913 84
rect 3948 50 3982 84
rect 4017 50 4051 84
rect 4086 50 4120 84
rect 4155 50 4189 84
rect 4224 50 4258 84
rect 4293 50 4327 84
rect 4362 50 4396 84
rect 4431 50 4465 84
rect 4500 50 4534 84
rect 4569 50 4603 84
rect 4638 50 4672 84
rect 4707 50 4741 84
rect 4776 50 4810 84
rect 4845 50 4879 84
rect 4914 50 4948 84
rect 4982 50 5016 84
rect 5050 50 5084 84
rect 5118 50 5152 84
rect 5186 50 5220 84
rect 5254 50 5288 84
rect 5322 50 5356 84
rect 5390 50 5424 84
rect 5458 50 5492 84
rect 5526 50 5560 84
rect 5594 50 5628 84
rect 5662 50 5696 84
rect 5730 50 5764 84
rect 5798 50 5832 84
rect 5866 50 5900 84
rect 5934 50 5968 84
rect 6002 50 6036 84
rect 6070 50 6104 84
rect 6138 50 6172 84
rect 6206 50 6240 84
rect 6274 50 6308 84
rect 6342 50 6376 84
rect 6410 50 6444 84
rect 6478 50 6512 84
rect 6546 50 6580 84
rect 6614 50 6648 84
rect 6682 50 6716 84
rect 6750 50 6784 84
rect 6818 50 6852 84
rect 6886 50 6920 84
rect 6954 50 6988 84
rect 7022 50 7056 84
rect 7090 50 7124 84
rect 7158 50 7192 84
rect 7226 50 7260 84
rect 7294 50 7328 84
rect 7362 50 7396 84
rect 7430 50 7464 84
rect 7498 50 7532 84
rect 7566 50 7600 84
rect 7634 50 7668 84
rect 7702 50 7736 84
rect 7770 50 7804 84
rect 7838 50 7872 84
rect 7906 50 7940 84
rect 7974 50 8008 84
rect 8042 50 8076 84
rect 8110 50 8144 84
rect 8178 50 8212 84
rect 8246 50 8280 84
rect 8314 50 8348 84
rect 8382 50 8416 84
rect 8450 50 8484 84
rect 8518 50 8552 84
rect 8586 50 8620 84
rect 8654 50 8688 84
rect 8722 50 8756 84
rect 8790 50 8824 84
rect 8858 50 8892 84
rect 8926 50 8960 84
rect 8994 50 9028 84
rect 9062 50 9096 84
rect 9130 50 9164 84
rect 9198 50 9232 84
rect 9266 50 9300 84
rect 9334 50 9368 84
rect 9402 50 9436 84
rect 9470 50 9504 84
rect 9538 50 9572 84
rect 9606 50 9640 84
rect 9674 50 9708 84
rect 9742 50 9776 84
rect 9810 50 9844 84
rect 9878 50 9912 84
rect 9946 50 9980 84
rect 10014 50 10048 84
rect 10082 50 10116 84
rect 10150 50 10184 84
rect 10218 50 10252 84
rect 10286 50 10320 84
rect 10354 50 10388 84
rect 10422 50 10456 84
rect 10490 50 10524 84
rect 10558 50 10592 84
rect 10626 50 10660 84
rect 10694 50 10728 84
rect 10762 50 10796 84
rect 10830 50 10864 84
rect 10898 50 10932 84
rect 10966 50 11000 84
rect 11034 50 11068 84
rect 11102 50 11136 84
rect 11170 50 11204 84
rect 11238 50 11272 84
rect 11306 50 11340 84
rect 11374 50 11408 84
rect 11442 50 11476 84
rect 11510 50 11544 84
rect 11578 50 11612 84
rect 11646 50 11680 84
rect 11714 50 11748 84
rect 11782 50 11816 84
rect 11850 50 11884 84
rect 11918 50 11952 84
rect 11986 50 12020 84
rect 12054 50 12088 84
rect 12122 50 12156 84
rect 12190 50 12224 84
rect 12258 50 12292 84
rect 12326 50 12360 84
rect 12394 50 12428 84
rect 12462 50 12496 84
rect 12530 50 12564 84
rect 12598 50 12632 84
rect 12666 50 12700 84
rect 12734 50 12768 84
rect 12802 50 12836 84
rect 12870 50 12904 84
rect 12938 50 12972 84
rect 13006 50 13040 84
rect 13074 50 13108 84
rect 13142 50 13176 84
rect 13210 50 13244 84
rect 13278 50 13312 84
rect 13346 50 13380 84
rect 13414 50 13448 84
rect 13482 50 13516 84
rect 13550 50 13584 84
rect 13618 50 13652 84
rect 13686 50 13720 84
rect 13754 50 13788 84
rect 13822 50 13856 84
rect 13890 50 13924 84
rect 13958 50 13992 84
rect 14026 50 14060 84
rect 14094 50 14128 84
rect 14162 50 14196 84
rect 14230 50 14264 84
rect 14298 50 14332 84
rect 14366 50 14400 84
rect 14434 50 14468 84
rect 14502 50 14536 84
rect 14570 50 14604 84
rect 14638 50 14672 84
rect 14706 50 14740 84
rect 14774 50 14808 84
rect 14842 50 14876 84
rect 14910 50 14944 84
rect 14978 50 15012 84
rect 15046 50 15080 84
rect 15114 50 15148 84
rect 15182 50 15216 84
rect 15250 50 15284 84
rect 15318 50 15352 84
rect 15386 50 15420 84
rect 15454 50 15488 84
rect 15522 50 15556 84
rect 15590 50 15624 84
rect 15658 50 15692 84
rect 15726 50 15760 84
rect 15794 50 15828 84
rect 15862 50 15896 84
rect 15930 50 15964 84
rect 15998 50 16032 84
<< mvpsubdiffcont >>
rect 360 3872 394 3906
rect 470 3875 504 3909
rect 538 3875 572 3909
rect 606 3875 640 3909
rect 674 3875 708 3909
rect 742 3875 776 3909
rect 810 3875 844 3909
rect 878 3875 912 3909
rect 946 3875 980 3909
rect 1014 3875 1048 3909
rect 1082 3875 1116 3909
rect 1150 3875 1184 3909
rect 1218 3875 1252 3909
rect 1286 3875 1320 3909
rect 1354 3875 1388 3909
rect 1422 3875 1456 3909
rect 1490 3875 1524 3909
rect 1558 3875 1592 3909
rect 1626 3875 1660 3909
rect 1694 3875 1728 3909
rect 1762 3875 1796 3909
rect 1830 3875 1864 3909
rect 1898 3875 1932 3909
rect 1966 3875 2000 3909
rect 2034 3875 2068 3909
rect 2102 3875 2136 3909
rect 2170 3875 2204 3909
rect 2238 3875 2272 3909
rect 2306 3875 2340 3909
rect 2374 3875 2408 3909
rect 2442 3875 2476 3909
rect 2510 3875 2544 3909
rect 2578 3875 2612 3909
rect 2646 3875 2680 3909
rect 2714 3875 2748 3909
rect 2782 3875 2816 3909
rect 2850 3875 2884 3909
rect 2918 3875 2952 3909
rect 2986 3875 3020 3909
rect 3054 3875 3088 3909
rect 3122 3875 3156 3909
rect 3190 3875 3224 3909
rect 3258 3875 3292 3909
rect 3326 3875 3360 3909
rect 3394 3875 3428 3909
rect 3462 3875 3496 3909
rect 3530 3875 3564 3909
rect 3598 3875 3632 3909
rect 3666 3875 3700 3909
rect 3734 3875 3768 3909
rect 3802 3875 3836 3909
rect 3870 3875 3904 3909
rect 3938 3875 3972 3909
rect 4006 3875 4040 3909
rect 4074 3875 4108 3909
rect 4142 3875 4176 3909
rect 4210 3875 4244 3909
rect 4278 3875 4312 3909
rect 4346 3875 4380 3909
rect 4414 3875 4448 3909
rect 4482 3875 4516 3909
rect 4550 3875 4584 3909
rect 4618 3875 4652 3909
rect 4686 3875 4720 3909
rect 4754 3875 4788 3909
rect 4822 3875 4856 3909
rect 4890 3875 4924 3909
rect 4958 3875 4992 3909
rect 5026 3875 5060 3909
rect 5094 3875 5128 3909
rect 5162 3875 5196 3909
rect 5230 3875 5264 3909
rect 5298 3875 5332 3909
rect 5366 3875 5400 3909
rect 5434 3875 5468 3909
rect 5502 3875 5536 3909
rect 5570 3875 5604 3909
rect 5638 3875 5672 3909
rect 5706 3875 5740 3909
rect 5774 3875 5808 3909
rect 5842 3875 5876 3909
rect 5910 3875 5944 3909
rect 5978 3875 6012 3909
rect 6046 3875 6080 3909
rect 6114 3875 6148 3909
rect 6182 3875 6216 3909
rect 6250 3875 6284 3909
rect 6318 3875 6352 3909
rect 6386 3875 6420 3909
rect 6454 3875 6488 3909
rect 6522 3875 6556 3909
rect 6590 3875 6624 3909
rect 6658 3875 6692 3909
rect 6726 3875 6760 3909
rect 6794 3875 6828 3909
rect 6862 3875 6896 3909
rect 6930 3875 6964 3909
rect 6998 3875 7032 3909
rect 7066 3875 7100 3909
rect 7134 3875 7168 3909
rect 7202 3875 7236 3909
rect 7270 3875 7304 3909
rect 7338 3875 7372 3909
rect 7406 3875 7440 3909
rect 7474 3875 7508 3909
rect 7542 3875 7576 3909
rect 7610 3875 7644 3909
rect 7678 3875 7712 3909
rect 7746 3875 7780 3909
rect 7814 3875 7848 3909
rect 7882 3875 7916 3909
rect 7950 3875 7984 3909
rect 8018 3875 8052 3909
rect 8086 3875 8120 3909
rect 8154 3875 8188 3909
rect 8222 3875 8256 3909
rect 8290 3875 8324 3909
rect 8359 3875 8393 3909
rect 8428 3875 8462 3909
rect 8497 3875 8531 3909
rect 8566 3875 8600 3909
rect 8635 3875 8669 3909
rect 8704 3875 8738 3909
rect 8773 3875 8807 3909
rect 8842 3875 8876 3909
rect 8911 3875 8945 3909
rect 8980 3875 9014 3909
rect 9049 3875 9083 3909
rect 9118 3875 9152 3909
rect 9187 3875 9221 3909
rect 9256 3875 9290 3909
rect 9325 3875 9359 3909
rect 9394 3875 9428 3909
rect 9463 3875 9497 3909
rect 9532 3875 9566 3909
rect 9601 3875 9635 3909
rect 9670 3875 9704 3909
rect 9739 3875 9773 3909
rect 9808 3875 9842 3909
rect 9877 3875 9911 3909
rect 9946 3875 9980 3909
rect 10015 3875 10049 3909
rect 10084 3875 10118 3909
rect 10153 3875 10187 3909
rect 10222 3875 10256 3909
rect 10291 3875 10325 3909
rect 10360 3875 10394 3909
rect 10429 3875 10463 3909
rect 10498 3875 10532 3909
rect 10567 3875 10601 3909
rect 10636 3875 10670 3909
rect 10705 3875 10739 3909
rect 10774 3875 10808 3909
rect 10843 3875 10877 3909
rect 10912 3875 10946 3909
rect 360 3801 394 3835
rect 360 3730 394 3764
rect 10912 3805 10946 3839
rect 10912 3735 10946 3769
rect 360 3659 394 3693
rect 360 3589 394 3623
rect 360 3519 394 3553
rect 360 3449 394 3483
rect 360 3379 394 3413
rect 360 3309 394 3343
rect 360 3239 394 3273
rect 360 3169 394 3203
rect 360 3099 394 3133
rect 360 3029 394 3063
rect 360 2959 394 2993
rect 360 2889 394 2923
rect 360 2819 394 2853
rect 360 2749 394 2783
rect 360 2679 394 2713
rect 360 2609 394 2643
rect 360 2539 394 2573
rect 360 2469 394 2503
rect 360 2399 394 2433
rect 360 2329 394 2363
rect 10912 3665 10946 3699
rect 10912 3595 10946 3629
rect 10912 3525 10946 3559
rect 10912 3455 10946 3489
rect 10912 3385 10946 3419
rect 10912 3315 10946 3349
rect 10912 3245 10946 3279
rect 10912 3175 10946 3209
rect 10912 3105 10946 3139
rect 10912 3035 10946 3069
rect 10912 2965 10946 2999
rect 10912 2895 10946 2929
rect 10912 2825 10946 2859
rect 10912 2755 10946 2789
rect 10912 2685 10946 2719
rect 10912 2615 10946 2649
rect 10912 2544 10946 2578
rect 10912 2473 10946 2507
rect 10912 2402 10946 2436
rect 10912 2331 10946 2365
rect 360 2259 394 2293
rect 10912 2260 10946 2294
rect 360 2189 394 2223
rect 429 2189 463 2223
rect 498 2189 532 2223
rect 567 2189 601 2223
rect 636 2189 670 2223
rect 705 2189 739 2223
rect 774 2189 808 2223
rect 843 2189 877 2223
rect 912 2189 946 2223
rect 981 2189 1015 2223
rect 1050 2189 1084 2223
rect 1119 2189 1153 2223
rect 1188 2189 1222 2223
rect 1256 2189 1290 2223
rect 1324 2189 1358 2223
rect 1392 2189 1426 2223
rect 1460 2189 1494 2223
rect 1528 2189 1562 2223
rect 1596 2189 1630 2223
rect 1664 2189 1698 2223
rect 1732 2189 1766 2223
rect 1800 2189 1834 2223
rect 1868 2189 1902 2223
rect 1936 2189 1970 2223
rect 2004 2189 2038 2223
rect 2072 2189 2106 2223
rect 2140 2189 2174 2223
rect 2208 2189 2242 2223
rect 2276 2189 2310 2223
rect 2344 2189 2378 2223
rect 2412 2189 2446 2223
rect 2480 2189 2514 2223
rect 2548 2189 2582 2223
rect 2616 2189 2650 2223
rect 2684 2189 2718 2223
rect 2752 2189 2786 2223
rect 2820 2189 2854 2223
rect 2888 2189 2922 2223
rect 2956 2189 2990 2223
rect 3024 2189 3058 2223
rect 3092 2189 3126 2223
rect 3160 2189 3194 2223
rect 3228 2189 3262 2223
rect 3296 2189 3330 2223
rect 3364 2189 3398 2223
rect 3432 2189 3466 2223
rect 3500 2189 3534 2223
rect 3568 2189 3602 2223
rect 3636 2189 3670 2223
rect 3704 2189 3738 2223
rect 3772 2189 3806 2223
rect 3840 2189 3874 2223
rect 3908 2189 3942 2223
rect 3976 2189 4010 2223
rect 4044 2189 4078 2223
rect 4112 2189 4146 2223
rect 4180 2189 4214 2223
rect 4248 2189 4282 2223
rect 4316 2189 4350 2223
rect 4384 2189 4418 2223
rect 4452 2189 4486 2223
rect 4520 2189 4554 2223
rect 4588 2189 4622 2223
rect 4656 2189 4690 2223
rect 4724 2189 4758 2223
rect 4792 2189 4826 2223
rect 4860 2189 4894 2223
rect 4928 2189 4962 2223
rect 4996 2189 5030 2223
rect 5064 2189 5098 2223
rect 5132 2189 5166 2223
rect 5200 2189 5234 2223
rect 5268 2189 5302 2223
rect 5336 2189 5370 2223
rect 5404 2189 5438 2223
rect 5472 2189 5506 2223
rect 5540 2189 5574 2223
rect 5608 2189 5642 2223
rect 5676 2189 5710 2223
rect 5744 2189 5778 2223
rect 5812 2189 5846 2223
rect 5880 2189 5914 2223
rect 5948 2189 5982 2223
rect 6016 2189 6050 2223
rect 6084 2189 6118 2223
rect 6152 2189 6186 2223
rect 6220 2189 6254 2223
rect 6288 2189 6322 2223
rect 6356 2189 6390 2223
rect 6424 2189 6458 2223
rect 6492 2189 6526 2223
rect 6560 2189 6594 2223
rect 6628 2189 6662 2223
rect 6696 2189 6730 2223
rect 6764 2189 6798 2223
rect 6832 2189 6866 2223
rect 6900 2189 6934 2223
rect 6968 2189 7002 2223
rect 7036 2189 7070 2223
rect 7104 2189 7138 2223
rect 7172 2189 7206 2223
rect 7240 2189 7274 2223
rect 7308 2189 7342 2223
rect 7376 2189 7410 2223
rect 7444 2189 7478 2223
rect 7512 2189 7546 2223
rect 7580 2189 7614 2223
rect 7648 2189 7682 2223
rect 7716 2189 7750 2223
rect 7784 2189 7818 2223
rect 7852 2189 7886 2223
rect 7920 2189 7954 2223
rect 7988 2189 8022 2223
rect 8056 2189 8090 2223
rect 8124 2189 8158 2223
rect 8192 2189 8226 2223
rect 8260 2189 8294 2223
rect 8328 2189 8362 2223
rect 8396 2189 8430 2223
rect 8464 2189 8498 2223
rect 8532 2189 8566 2223
rect 8600 2189 8634 2223
rect 8668 2189 8702 2223
rect 8736 2189 8770 2223
rect 8804 2189 8838 2223
rect 8872 2189 8906 2223
rect 8940 2189 8974 2223
rect 9008 2189 9042 2223
rect 9076 2189 9110 2223
rect 9144 2189 9178 2223
rect 9212 2189 9246 2223
rect 9280 2189 9314 2223
rect 9348 2189 9382 2223
rect 9416 2189 9450 2223
rect 9484 2189 9518 2223
rect 9552 2189 9586 2223
rect 9620 2189 9654 2223
rect 9688 2189 9722 2223
rect 9756 2189 9790 2223
rect 9824 2189 9858 2223
rect 9892 2189 9926 2223
rect 9960 2189 9994 2223
rect 10028 2189 10062 2223
rect 10096 2189 10130 2223
rect 10164 2189 10198 2223
rect 10232 2189 10266 2223
rect 10300 2189 10334 2223
rect 10368 2189 10402 2223
rect 10436 2189 10470 2223
rect 10504 2189 10538 2223
rect 10572 2189 10606 2223
rect 10640 2189 10674 2223
rect 10708 2189 10742 2223
rect 10776 2189 10810 2223
rect 10844 2189 10878 2223
rect 10912 2189 10946 2223
<< mvnsubdiffcont >>
rect 360 5765 394 5799
rect 428 5765 462 5799
rect 496 5765 530 5799
rect 564 5765 598 5799
rect 632 5765 666 5799
rect 700 5765 734 5799
rect 768 5765 802 5799
rect 836 5765 870 5799
rect 904 5765 938 5799
rect 972 5765 1006 5799
rect 1040 5765 1074 5799
rect 1108 5765 1142 5799
rect 1176 5765 1210 5799
rect 1244 5765 1278 5799
rect 1312 5765 1346 5799
rect 1380 5765 1414 5799
rect 1448 5765 1482 5799
rect 1516 5765 1550 5799
rect 1584 5765 1618 5799
rect 1652 5765 1686 5799
rect 1720 5765 1754 5799
rect 1788 5765 1822 5799
rect 1856 5765 1890 5799
rect 1924 5765 1958 5799
rect 1992 5765 2026 5799
rect 2060 5765 2094 5799
rect 2128 5765 2162 5799
rect 2196 5765 2230 5799
rect 2264 5765 2298 5799
rect 2332 5765 2366 5799
rect 2400 5765 2434 5799
rect 2468 5765 2502 5799
rect 2536 5765 2570 5799
rect 2604 5765 2638 5799
rect 2672 5765 2706 5799
rect 2740 5765 2774 5799
rect 2808 5765 2842 5799
rect 2876 5765 2910 5799
rect 2944 5765 2978 5799
rect 3012 5765 3046 5799
rect 3080 5765 3114 5799
rect 3148 5765 3182 5799
rect 3216 5765 3250 5799
rect 3284 5765 3318 5799
rect 3352 5765 3386 5799
rect 3420 5765 3454 5799
rect 3488 5765 3522 5799
rect 3556 5765 3590 5799
rect 3624 5765 3658 5799
rect 3692 5765 3726 5799
rect 3760 5765 3794 5799
rect 3828 5765 3862 5799
rect 3896 5765 3930 5799
rect 3964 5765 3998 5799
rect 4032 5765 4066 5799
rect 4100 5765 4134 5799
rect 4168 5765 4202 5799
rect 4236 5765 4270 5799
rect 4304 5765 4338 5799
rect 4372 5765 4406 5799
rect 4440 5765 4474 5799
rect 4508 5765 4542 5799
rect 4576 5765 4610 5799
rect 4644 5765 4678 5799
rect 4712 5765 4746 5799
rect 4780 5765 4814 5799
rect 4848 5765 4882 5799
rect 4916 5765 4950 5799
rect 4984 5765 5018 5799
rect 5052 5765 5086 5799
rect 5120 5765 5154 5799
rect 5188 5765 5222 5799
rect 5256 5765 5290 5799
rect 5324 5765 5358 5799
rect 5392 5765 5426 5799
rect 5460 5765 5494 5799
rect 5528 5765 5562 5799
rect 5596 5765 5630 5799
rect 5664 5765 5698 5799
rect 5732 5765 5766 5799
rect 5800 5765 5834 5799
rect 5868 5765 5902 5799
rect 5936 5765 5970 5799
rect 6004 5765 6038 5799
rect 6072 5765 6106 5799
rect 6140 5765 6174 5799
rect 6208 5765 6242 5799
rect 6276 5765 6310 5799
rect 6344 5765 6378 5799
rect 6412 5765 6446 5799
rect 6480 5765 6514 5799
rect 6548 5765 6582 5799
rect 6616 5765 6650 5799
rect 6684 5765 6718 5799
rect 6752 5765 6786 5799
rect 6820 5765 6854 5799
rect 6888 5765 6922 5799
rect 6956 5765 6990 5799
rect 7024 5765 7058 5799
rect 7092 5765 7126 5799
rect 7160 5765 7194 5799
rect 7228 5765 7262 5799
rect 7296 5765 7330 5799
rect 7364 5765 7398 5799
rect 7432 5765 7466 5799
rect 7500 5765 7534 5799
rect 7568 5765 7602 5799
rect 7636 5765 7670 5799
rect 7704 5765 7738 5799
rect 7772 5765 7806 5799
rect 7840 5765 7874 5799
rect 7908 5765 7942 5799
rect 7976 5765 8010 5799
rect 8044 5765 8078 5799
rect 8112 5765 8146 5799
rect 8181 5765 8215 5799
rect 8250 5765 8284 5799
rect 8319 5765 8353 5799
rect 8388 5765 8422 5799
rect 8457 5765 8491 5799
rect 8526 5765 8560 5799
rect 8595 5765 8629 5799
rect 8664 5765 8698 5799
rect 8733 5765 8767 5799
rect 8802 5765 8836 5799
rect 8871 5765 8905 5799
rect 8940 5765 8974 5799
rect 9009 5765 9043 5799
rect 9078 5765 9112 5799
rect 9147 5765 9181 5799
rect 9216 5765 9250 5799
rect 9285 5765 9319 5799
rect 9354 5765 9388 5799
rect 9423 5765 9457 5799
rect 9492 5765 9526 5799
rect 9561 5765 9595 5799
rect 9630 5765 9664 5799
rect 9699 5765 9733 5799
rect 9768 5765 9802 5799
rect 9837 5765 9871 5799
rect 9906 5765 9940 5799
rect 9975 5765 10009 5799
rect 10044 5765 10078 5799
rect 10113 5765 10147 5799
rect 10182 5765 10216 5799
rect 10251 5765 10285 5799
rect 10320 5765 10354 5799
rect 10389 5765 10423 5799
rect 10458 5765 10492 5799
rect 10527 5765 10561 5799
rect 10596 5765 10630 5799
rect 10665 5765 10699 5799
rect 10734 5765 10768 5799
rect 10803 5765 10837 5799
rect 10872 5765 10906 5799
rect 360 5690 394 5724
rect 10872 5696 10906 5730
rect 360 5615 394 5649
rect 360 5541 394 5575
rect 360 5467 394 5501
rect 360 5393 394 5427
rect 360 5287 394 5321
rect 360 5217 394 5251
rect 360 5147 394 5181
rect 360 5077 394 5111
rect 360 5007 394 5041
rect 360 4937 394 4971
rect 360 4868 394 4902
rect 360 4799 394 4833
rect 360 4730 394 4764
rect 360 4661 394 4695
rect 360 4592 394 4626
rect 360 4523 394 4557
rect 360 4454 394 4488
rect 360 4385 394 4419
rect 360 4316 394 4350
rect 10872 5627 10906 5661
rect 10872 5558 10906 5592
rect 10872 5489 10906 5523
rect 10872 5420 10906 5454
rect 10872 5351 10906 5385
rect 10872 5282 10906 5316
rect 10872 5213 10906 5247
rect 10872 5144 10906 5178
rect 10872 5075 10906 5109
rect 10872 5006 10906 5040
rect 10872 4937 10906 4971
rect 10872 4868 10906 4902
rect 10872 4799 10906 4833
rect 10872 4730 10906 4764
rect 10872 4661 10906 4695
rect 10872 4592 10906 4626
rect 10872 4523 10906 4557
rect 10872 4454 10906 4488
rect 10872 4385 10906 4419
rect 10872 4316 10906 4350
rect 360 4247 394 4281
rect 360 4178 394 4212
rect 10872 4247 10906 4281
rect 10872 4178 10906 4212
rect 360 4109 394 4143
rect 429 4109 463 4143
rect 498 4109 532 4143
rect 567 4109 601 4143
rect 636 4109 670 4143
rect 705 4109 739 4143
rect 774 4109 808 4143
rect 843 4109 877 4143
rect 912 4109 946 4143
rect 981 4109 1015 4143
rect 1050 4109 1084 4143
rect 1119 4109 1153 4143
rect 1188 4109 1222 4143
rect 1257 4109 1291 4143
rect 1326 4109 1360 4143
rect 1395 4109 1429 4143
rect 1464 4109 1498 4143
rect 1533 4109 1567 4143
rect 1602 4109 1636 4143
rect 1671 4109 1705 4143
rect 1740 4109 1774 4143
rect 1809 4109 1843 4143
rect 1878 4109 1912 4143
rect 1947 4109 1981 4143
rect 2016 4109 2050 4143
rect 2085 4109 2119 4143
rect 2154 4109 2188 4143
rect 2223 4109 2257 4143
rect 2292 4109 2326 4143
rect 2361 4109 2395 4143
rect 2430 4109 2464 4143
rect 2499 4109 2533 4143
rect 2568 4109 2602 4143
rect 2637 4109 2671 4143
rect 2706 4109 2740 4143
rect 2775 4109 2809 4143
rect 2844 4109 2878 4143
rect 2913 4109 2947 4143
rect 2982 4109 3016 4143
rect 3051 4109 3085 4143
rect 3120 4109 3154 4143
rect 3188 4109 3222 4143
rect 3256 4109 3290 4143
rect 3324 4109 3358 4143
rect 3392 4109 3426 4143
rect 3460 4109 3494 4143
rect 3528 4109 3562 4143
rect 3596 4109 3630 4143
rect 3664 4109 3698 4143
rect 3732 4109 3766 4143
rect 3800 4109 3834 4143
rect 3868 4109 3902 4143
rect 3936 4109 3970 4143
rect 4004 4109 4038 4143
rect 4072 4109 4106 4143
rect 4140 4109 4174 4143
rect 4208 4109 4242 4143
rect 4276 4109 4310 4143
rect 4344 4109 4378 4143
rect 4412 4109 4446 4143
rect 4480 4109 4514 4143
rect 4548 4109 4582 4143
rect 4616 4109 4650 4143
rect 4684 4109 4718 4143
rect 4752 4109 4786 4143
rect 4820 4109 4854 4143
rect 4888 4109 4922 4143
rect 4956 4109 4990 4143
rect 5024 4109 5058 4143
rect 5092 4109 5126 4143
rect 5160 4109 5194 4143
rect 5228 4109 5262 4143
rect 5296 4109 5330 4143
rect 5364 4109 5398 4143
rect 5432 4109 5466 4143
rect 5500 4109 5534 4143
rect 5568 4109 5602 4143
rect 5636 4109 5670 4143
rect 5704 4109 5738 4143
rect 5772 4109 5806 4143
rect 5840 4109 5874 4143
rect 5908 4109 5942 4143
rect 5976 4109 6010 4143
rect 6044 4109 6078 4143
rect 6112 4109 6146 4143
rect 6180 4109 6214 4143
rect 6248 4109 6282 4143
rect 6316 4109 6350 4143
rect 6384 4109 6418 4143
rect 6452 4109 6486 4143
rect 6520 4109 6554 4143
rect 6588 4109 6622 4143
rect 6656 4109 6690 4143
rect 6724 4109 6758 4143
rect 6792 4109 6826 4143
rect 6860 4109 6894 4143
rect 6928 4109 6962 4143
rect 6996 4109 7030 4143
rect 7064 4109 7098 4143
rect 7132 4109 7166 4143
rect 7200 4109 7234 4143
rect 7268 4109 7302 4143
rect 7336 4109 7370 4143
rect 7404 4109 7438 4143
rect 7472 4109 7506 4143
rect 7540 4109 7574 4143
rect 7608 4109 7642 4143
rect 7676 4109 7710 4143
rect 7744 4109 7778 4143
rect 7812 4109 7846 4143
rect 7880 4109 7914 4143
rect 7948 4109 7982 4143
rect 8016 4109 8050 4143
rect 8084 4109 8118 4143
rect 8152 4109 8186 4143
rect 8220 4109 8254 4143
rect 8288 4109 8322 4143
rect 8356 4109 8390 4143
rect 8424 4109 8458 4143
rect 8492 4109 8526 4143
rect 8560 4109 8594 4143
rect 8628 4109 8662 4143
rect 8696 4109 8730 4143
rect 8764 4109 8798 4143
rect 8832 4109 8866 4143
rect 8900 4109 8934 4143
rect 8968 4109 9002 4143
rect 9036 4109 9070 4143
rect 9104 4109 9138 4143
rect 9172 4109 9206 4143
rect 9240 4109 9274 4143
rect 9308 4109 9342 4143
rect 9376 4109 9410 4143
rect 9444 4109 9478 4143
rect 9512 4109 9546 4143
rect 9580 4109 9614 4143
rect 9648 4109 9682 4143
rect 9716 4109 9750 4143
rect 9784 4109 9818 4143
rect 9852 4109 9886 4143
rect 9920 4109 9954 4143
rect 9988 4109 10022 4143
rect 10056 4109 10090 4143
rect 10124 4109 10158 4143
rect 10192 4109 10226 4143
rect 10260 4109 10294 4143
rect 10328 4109 10362 4143
rect 10396 4109 10430 4143
rect 10464 4109 10498 4143
rect 10532 4109 10566 4143
rect 10600 4109 10634 4143
rect 10668 4109 10702 4143
rect 10736 4109 10770 4143
rect 10804 4109 10838 4143
rect 10872 4109 10906 4143
<< poly >>
rect 525 5687 1325 5713
rect 1381 5687 2181 5713
rect 2237 5687 3037 5713
rect 3093 5687 3893 5713
rect 3949 5687 4749 5713
rect 4805 5687 5605 5713
rect 5661 5687 6461 5713
rect 6517 5687 7317 5713
rect 7373 5687 8173 5713
rect 8229 5687 9029 5713
rect 9085 5687 9885 5713
rect 9941 5687 10741 5713
rect 525 4239 1325 4287
rect 525 4205 568 4239
rect 602 4205 636 4239
rect 670 4205 704 4239
rect 738 4205 772 4239
rect 806 4205 840 4239
rect 874 4205 908 4239
rect 942 4205 976 4239
rect 1010 4205 1044 4239
rect 1078 4205 1112 4239
rect 1146 4205 1180 4239
rect 1214 4205 1248 4239
rect 1282 4205 1325 4239
rect 525 4189 1325 4205
rect 1381 4239 2181 4287
rect 1381 4205 1424 4239
rect 1458 4205 1492 4239
rect 1526 4205 1560 4239
rect 1594 4205 1628 4239
rect 1662 4205 1696 4239
rect 1730 4205 1764 4239
rect 1798 4205 1832 4239
rect 1866 4205 1900 4239
rect 1934 4205 1968 4239
rect 2002 4205 2036 4239
rect 2070 4205 2104 4239
rect 2138 4205 2181 4239
rect 1381 4189 2181 4205
rect 2237 4239 3037 4287
rect 2237 4205 2280 4239
rect 2314 4205 2348 4239
rect 2382 4205 2416 4239
rect 2450 4205 2484 4239
rect 2518 4205 2552 4239
rect 2586 4205 2620 4239
rect 2654 4205 2688 4239
rect 2722 4205 2756 4239
rect 2790 4205 2824 4239
rect 2858 4205 2892 4239
rect 2926 4205 2960 4239
rect 2994 4205 3037 4239
rect 2237 4189 3037 4205
rect 3093 4239 3893 4287
rect 3093 4205 3136 4239
rect 3170 4205 3204 4239
rect 3238 4205 3272 4239
rect 3306 4205 3340 4239
rect 3374 4205 3408 4239
rect 3442 4205 3476 4239
rect 3510 4205 3544 4239
rect 3578 4205 3612 4239
rect 3646 4205 3680 4239
rect 3714 4205 3748 4239
rect 3782 4205 3816 4239
rect 3850 4205 3893 4239
rect 3093 4189 3893 4205
rect 3949 4239 4749 4287
rect 3949 4205 3992 4239
rect 4026 4205 4060 4239
rect 4094 4205 4128 4239
rect 4162 4205 4196 4239
rect 4230 4205 4264 4239
rect 4298 4205 4332 4239
rect 4366 4205 4400 4239
rect 4434 4205 4468 4239
rect 4502 4205 4536 4239
rect 4570 4205 4604 4239
rect 4638 4205 4672 4239
rect 4706 4205 4749 4239
rect 3949 4189 4749 4205
rect 4805 4239 5605 4287
rect 4805 4205 4848 4239
rect 4882 4205 4916 4239
rect 4950 4205 4984 4239
rect 5018 4205 5052 4239
rect 5086 4205 5120 4239
rect 5154 4205 5188 4239
rect 5222 4205 5256 4239
rect 5290 4205 5324 4239
rect 5358 4205 5392 4239
rect 5426 4205 5460 4239
rect 5494 4205 5528 4239
rect 5562 4205 5605 4239
rect 4805 4189 5605 4205
rect 5661 4239 6461 4287
rect 5661 4205 5704 4239
rect 5738 4205 5772 4239
rect 5806 4205 5840 4239
rect 5874 4205 5908 4239
rect 5942 4205 5976 4239
rect 6010 4205 6044 4239
rect 6078 4205 6112 4239
rect 6146 4205 6180 4239
rect 6214 4205 6248 4239
rect 6282 4205 6316 4239
rect 6350 4205 6384 4239
rect 6418 4205 6461 4239
rect 5661 4189 6461 4205
rect 6517 4239 7317 4287
rect 6517 4205 6560 4239
rect 6594 4205 6628 4239
rect 6662 4205 6696 4239
rect 6730 4205 6764 4239
rect 6798 4205 6832 4239
rect 6866 4205 6900 4239
rect 6934 4205 6968 4239
rect 7002 4205 7036 4239
rect 7070 4205 7104 4239
rect 7138 4205 7172 4239
rect 7206 4205 7240 4239
rect 7274 4205 7317 4239
rect 6517 4189 7317 4205
rect 7373 4239 8173 4287
rect 7373 4205 7416 4239
rect 7450 4205 7484 4239
rect 7518 4205 7552 4239
rect 7586 4205 7620 4239
rect 7654 4205 7688 4239
rect 7722 4205 7756 4239
rect 7790 4205 7824 4239
rect 7858 4205 7892 4239
rect 7926 4205 7960 4239
rect 7994 4205 8028 4239
rect 8062 4205 8096 4239
rect 8130 4205 8173 4239
rect 7373 4189 8173 4205
rect 8229 4239 9029 4287
rect 8229 4205 8272 4239
rect 8306 4205 8340 4239
rect 8374 4205 8408 4239
rect 8442 4205 8476 4239
rect 8510 4205 8544 4239
rect 8578 4205 8612 4239
rect 8646 4205 8680 4239
rect 8714 4205 8748 4239
rect 8782 4205 8816 4239
rect 8850 4205 8884 4239
rect 8918 4205 8952 4239
rect 8986 4205 9029 4239
rect 8229 4189 9029 4205
rect 9085 4239 9885 4287
rect 9085 4205 9128 4239
rect 9162 4205 9196 4239
rect 9230 4205 9264 4239
rect 9298 4205 9332 4239
rect 9366 4205 9400 4239
rect 9434 4205 9468 4239
rect 9502 4205 9536 4239
rect 9570 4205 9604 4239
rect 9638 4205 9672 4239
rect 9706 4205 9740 4239
rect 9774 4205 9808 4239
rect 9842 4205 9885 4239
rect 9085 4189 9885 4205
rect 9941 4239 10741 4287
rect 9941 4205 9984 4239
rect 10018 4205 10052 4239
rect 10086 4205 10120 4239
rect 10154 4205 10188 4239
rect 10222 4205 10256 4239
rect 10290 4205 10324 4239
rect 10358 4205 10392 4239
rect 10426 4205 10460 4239
rect 10494 4205 10528 4239
rect 10562 4205 10596 4239
rect 10630 4205 10664 4239
rect 10698 4205 10741 4239
rect 9941 4189 10741 4205
rect 545 3803 1345 3819
rect 545 3769 588 3803
rect 622 3769 656 3803
rect 690 3769 724 3803
rect 758 3769 792 3803
rect 826 3769 860 3803
rect 894 3769 928 3803
rect 962 3769 996 3803
rect 1030 3769 1064 3803
rect 1098 3769 1132 3803
rect 1166 3769 1200 3803
rect 1234 3769 1268 3803
rect 1302 3769 1345 3803
rect 545 3721 1345 3769
rect 1401 3803 2201 3819
rect 1401 3769 1444 3803
rect 1478 3769 1512 3803
rect 1546 3769 1580 3803
rect 1614 3769 1648 3803
rect 1682 3769 1716 3803
rect 1750 3769 1784 3803
rect 1818 3769 1852 3803
rect 1886 3769 1920 3803
rect 1954 3769 1988 3803
rect 2022 3769 2056 3803
rect 2090 3769 2124 3803
rect 2158 3769 2201 3803
rect 1401 3721 2201 3769
rect 2257 3803 3057 3819
rect 2257 3769 2300 3803
rect 2334 3769 2368 3803
rect 2402 3769 2436 3803
rect 2470 3769 2504 3803
rect 2538 3769 2572 3803
rect 2606 3769 2640 3803
rect 2674 3769 2708 3803
rect 2742 3769 2776 3803
rect 2810 3769 2844 3803
rect 2878 3769 2912 3803
rect 2946 3769 2980 3803
rect 3014 3769 3057 3803
rect 2257 3721 3057 3769
rect 3113 3803 3913 3819
rect 3113 3769 3156 3803
rect 3190 3769 3224 3803
rect 3258 3769 3292 3803
rect 3326 3769 3360 3803
rect 3394 3769 3428 3803
rect 3462 3769 3496 3803
rect 3530 3769 3564 3803
rect 3598 3769 3632 3803
rect 3666 3769 3700 3803
rect 3734 3769 3768 3803
rect 3802 3769 3836 3803
rect 3870 3769 3913 3803
rect 3113 3721 3913 3769
rect 3969 3803 4769 3819
rect 3969 3769 4012 3803
rect 4046 3769 4080 3803
rect 4114 3769 4148 3803
rect 4182 3769 4216 3803
rect 4250 3769 4284 3803
rect 4318 3769 4352 3803
rect 4386 3769 4420 3803
rect 4454 3769 4488 3803
rect 4522 3769 4556 3803
rect 4590 3769 4624 3803
rect 4658 3769 4692 3803
rect 4726 3769 4769 3803
rect 3969 3721 4769 3769
rect 4825 3803 5625 3819
rect 4825 3769 4868 3803
rect 4902 3769 4936 3803
rect 4970 3769 5004 3803
rect 5038 3769 5072 3803
rect 5106 3769 5140 3803
rect 5174 3769 5208 3803
rect 5242 3769 5276 3803
rect 5310 3769 5344 3803
rect 5378 3769 5412 3803
rect 5446 3769 5480 3803
rect 5514 3769 5548 3803
rect 5582 3769 5625 3803
rect 4825 3721 5625 3769
rect 5681 3803 6481 3819
rect 5681 3769 5724 3803
rect 5758 3769 5792 3803
rect 5826 3769 5860 3803
rect 5894 3769 5928 3803
rect 5962 3769 5996 3803
rect 6030 3769 6064 3803
rect 6098 3769 6132 3803
rect 6166 3769 6200 3803
rect 6234 3769 6268 3803
rect 6302 3769 6336 3803
rect 6370 3769 6404 3803
rect 6438 3769 6481 3803
rect 5681 3721 6481 3769
rect 6537 3803 7337 3819
rect 6537 3769 6580 3803
rect 6614 3769 6648 3803
rect 6682 3769 6716 3803
rect 6750 3769 6784 3803
rect 6818 3769 6852 3803
rect 6886 3769 6920 3803
rect 6954 3769 6988 3803
rect 7022 3769 7056 3803
rect 7090 3769 7124 3803
rect 7158 3769 7192 3803
rect 7226 3769 7260 3803
rect 7294 3769 7337 3803
rect 6537 3721 7337 3769
rect 7393 3803 8193 3819
rect 7393 3769 7436 3803
rect 7470 3769 7504 3803
rect 7538 3769 7572 3803
rect 7606 3769 7640 3803
rect 7674 3769 7708 3803
rect 7742 3769 7776 3803
rect 7810 3769 7844 3803
rect 7878 3769 7912 3803
rect 7946 3769 7980 3803
rect 8014 3769 8048 3803
rect 8082 3769 8116 3803
rect 8150 3769 8193 3803
rect 7393 3721 8193 3769
rect 8249 3803 9049 3819
rect 8249 3769 8292 3803
rect 8326 3769 8360 3803
rect 8394 3769 8428 3803
rect 8462 3769 8496 3803
rect 8530 3769 8564 3803
rect 8598 3769 8632 3803
rect 8666 3769 8700 3803
rect 8734 3769 8768 3803
rect 8802 3769 8836 3803
rect 8870 3769 8904 3803
rect 8938 3769 8972 3803
rect 9006 3769 9049 3803
rect 8249 3721 9049 3769
rect 9105 3803 9905 3819
rect 9105 3769 9148 3803
rect 9182 3769 9216 3803
rect 9250 3769 9284 3803
rect 9318 3769 9352 3803
rect 9386 3769 9420 3803
rect 9454 3769 9488 3803
rect 9522 3769 9556 3803
rect 9590 3769 9624 3803
rect 9658 3769 9692 3803
rect 9726 3769 9760 3803
rect 9794 3769 9828 3803
rect 9862 3769 9905 3803
rect 9105 3721 9905 3769
rect 9961 3803 10761 3819
rect 9961 3769 10004 3803
rect 10038 3769 10072 3803
rect 10106 3769 10140 3803
rect 10174 3769 10208 3803
rect 10242 3769 10276 3803
rect 10310 3769 10344 3803
rect 10378 3769 10412 3803
rect 10446 3769 10480 3803
rect 10514 3769 10548 3803
rect 10582 3769 10616 3803
rect 10650 3769 10684 3803
rect 10718 3769 10761 3803
rect 9961 3721 10761 3769
rect 545 2295 1345 2321
rect 1401 2295 2201 2321
rect 2257 2295 3057 2321
rect 3113 2295 3913 2321
rect 3969 2295 4769 2321
rect 4825 2295 5625 2321
rect 5681 2295 6481 2321
rect 6537 2295 7337 2321
rect 7393 2295 8193 2321
rect 8249 2295 9049 2321
rect 9105 2295 9905 2321
rect 9961 2295 10761 2321
<< polycont >>
rect 568 4205 602 4239
rect 636 4205 670 4239
rect 704 4205 738 4239
rect 772 4205 806 4239
rect 840 4205 874 4239
rect 908 4205 942 4239
rect 976 4205 1010 4239
rect 1044 4205 1078 4239
rect 1112 4205 1146 4239
rect 1180 4205 1214 4239
rect 1248 4205 1282 4239
rect 1424 4205 1458 4239
rect 1492 4205 1526 4239
rect 1560 4205 1594 4239
rect 1628 4205 1662 4239
rect 1696 4205 1730 4239
rect 1764 4205 1798 4239
rect 1832 4205 1866 4239
rect 1900 4205 1934 4239
rect 1968 4205 2002 4239
rect 2036 4205 2070 4239
rect 2104 4205 2138 4239
rect 2280 4205 2314 4239
rect 2348 4205 2382 4239
rect 2416 4205 2450 4239
rect 2484 4205 2518 4239
rect 2552 4205 2586 4239
rect 2620 4205 2654 4239
rect 2688 4205 2722 4239
rect 2756 4205 2790 4239
rect 2824 4205 2858 4239
rect 2892 4205 2926 4239
rect 2960 4205 2994 4239
rect 3136 4205 3170 4239
rect 3204 4205 3238 4239
rect 3272 4205 3306 4239
rect 3340 4205 3374 4239
rect 3408 4205 3442 4239
rect 3476 4205 3510 4239
rect 3544 4205 3578 4239
rect 3612 4205 3646 4239
rect 3680 4205 3714 4239
rect 3748 4205 3782 4239
rect 3816 4205 3850 4239
rect 3992 4205 4026 4239
rect 4060 4205 4094 4239
rect 4128 4205 4162 4239
rect 4196 4205 4230 4239
rect 4264 4205 4298 4239
rect 4332 4205 4366 4239
rect 4400 4205 4434 4239
rect 4468 4205 4502 4239
rect 4536 4205 4570 4239
rect 4604 4205 4638 4239
rect 4672 4205 4706 4239
rect 4848 4205 4882 4239
rect 4916 4205 4950 4239
rect 4984 4205 5018 4239
rect 5052 4205 5086 4239
rect 5120 4205 5154 4239
rect 5188 4205 5222 4239
rect 5256 4205 5290 4239
rect 5324 4205 5358 4239
rect 5392 4205 5426 4239
rect 5460 4205 5494 4239
rect 5528 4205 5562 4239
rect 5704 4205 5738 4239
rect 5772 4205 5806 4239
rect 5840 4205 5874 4239
rect 5908 4205 5942 4239
rect 5976 4205 6010 4239
rect 6044 4205 6078 4239
rect 6112 4205 6146 4239
rect 6180 4205 6214 4239
rect 6248 4205 6282 4239
rect 6316 4205 6350 4239
rect 6384 4205 6418 4239
rect 6560 4205 6594 4239
rect 6628 4205 6662 4239
rect 6696 4205 6730 4239
rect 6764 4205 6798 4239
rect 6832 4205 6866 4239
rect 6900 4205 6934 4239
rect 6968 4205 7002 4239
rect 7036 4205 7070 4239
rect 7104 4205 7138 4239
rect 7172 4205 7206 4239
rect 7240 4205 7274 4239
rect 7416 4205 7450 4239
rect 7484 4205 7518 4239
rect 7552 4205 7586 4239
rect 7620 4205 7654 4239
rect 7688 4205 7722 4239
rect 7756 4205 7790 4239
rect 7824 4205 7858 4239
rect 7892 4205 7926 4239
rect 7960 4205 7994 4239
rect 8028 4205 8062 4239
rect 8096 4205 8130 4239
rect 8272 4205 8306 4239
rect 8340 4205 8374 4239
rect 8408 4205 8442 4239
rect 8476 4205 8510 4239
rect 8544 4205 8578 4239
rect 8612 4205 8646 4239
rect 8680 4205 8714 4239
rect 8748 4205 8782 4239
rect 8816 4205 8850 4239
rect 8884 4205 8918 4239
rect 8952 4205 8986 4239
rect 9128 4205 9162 4239
rect 9196 4205 9230 4239
rect 9264 4205 9298 4239
rect 9332 4205 9366 4239
rect 9400 4205 9434 4239
rect 9468 4205 9502 4239
rect 9536 4205 9570 4239
rect 9604 4205 9638 4239
rect 9672 4205 9706 4239
rect 9740 4205 9774 4239
rect 9808 4205 9842 4239
rect 9984 4205 10018 4239
rect 10052 4205 10086 4239
rect 10120 4205 10154 4239
rect 10188 4205 10222 4239
rect 10256 4205 10290 4239
rect 10324 4205 10358 4239
rect 10392 4205 10426 4239
rect 10460 4205 10494 4239
rect 10528 4205 10562 4239
rect 10596 4205 10630 4239
rect 10664 4205 10698 4239
rect 588 3769 622 3803
rect 656 3769 690 3803
rect 724 3769 758 3803
rect 792 3769 826 3803
rect 860 3769 894 3803
rect 928 3769 962 3803
rect 996 3769 1030 3803
rect 1064 3769 1098 3803
rect 1132 3769 1166 3803
rect 1200 3769 1234 3803
rect 1268 3769 1302 3803
rect 1444 3769 1478 3803
rect 1512 3769 1546 3803
rect 1580 3769 1614 3803
rect 1648 3769 1682 3803
rect 1716 3769 1750 3803
rect 1784 3769 1818 3803
rect 1852 3769 1886 3803
rect 1920 3769 1954 3803
rect 1988 3769 2022 3803
rect 2056 3769 2090 3803
rect 2124 3769 2158 3803
rect 2300 3769 2334 3803
rect 2368 3769 2402 3803
rect 2436 3769 2470 3803
rect 2504 3769 2538 3803
rect 2572 3769 2606 3803
rect 2640 3769 2674 3803
rect 2708 3769 2742 3803
rect 2776 3769 2810 3803
rect 2844 3769 2878 3803
rect 2912 3769 2946 3803
rect 2980 3769 3014 3803
rect 3156 3769 3190 3803
rect 3224 3769 3258 3803
rect 3292 3769 3326 3803
rect 3360 3769 3394 3803
rect 3428 3769 3462 3803
rect 3496 3769 3530 3803
rect 3564 3769 3598 3803
rect 3632 3769 3666 3803
rect 3700 3769 3734 3803
rect 3768 3769 3802 3803
rect 3836 3769 3870 3803
rect 4012 3769 4046 3803
rect 4080 3769 4114 3803
rect 4148 3769 4182 3803
rect 4216 3769 4250 3803
rect 4284 3769 4318 3803
rect 4352 3769 4386 3803
rect 4420 3769 4454 3803
rect 4488 3769 4522 3803
rect 4556 3769 4590 3803
rect 4624 3769 4658 3803
rect 4692 3769 4726 3803
rect 4868 3769 4902 3803
rect 4936 3769 4970 3803
rect 5004 3769 5038 3803
rect 5072 3769 5106 3803
rect 5140 3769 5174 3803
rect 5208 3769 5242 3803
rect 5276 3769 5310 3803
rect 5344 3769 5378 3803
rect 5412 3769 5446 3803
rect 5480 3769 5514 3803
rect 5548 3769 5582 3803
rect 5724 3769 5758 3803
rect 5792 3769 5826 3803
rect 5860 3769 5894 3803
rect 5928 3769 5962 3803
rect 5996 3769 6030 3803
rect 6064 3769 6098 3803
rect 6132 3769 6166 3803
rect 6200 3769 6234 3803
rect 6268 3769 6302 3803
rect 6336 3769 6370 3803
rect 6404 3769 6438 3803
rect 6580 3769 6614 3803
rect 6648 3769 6682 3803
rect 6716 3769 6750 3803
rect 6784 3769 6818 3803
rect 6852 3769 6886 3803
rect 6920 3769 6954 3803
rect 6988 3769 7022 3803
rect 7056 3769 7090 3803
rect 7124 3769 7158 3803
rect 7192 3769 7226 3803
rect 7260 3769 7294 3803
rect 7436 3769 7470 3803
rect 7504 3769 7538 3803
rect 7572 3769 7606 3803
rect 7640 3769 7674 3803
rect 7708 3769 7742 3803
rect 7776 3769 7810 3803
rect 7844 3769 7878 3803
rect 7912 3769 7946 3803
rect 7980 3769 8014 3803
rect 8048 3769 8082 3803
rect 8116 3769 8150 3803
rect 8292 3769 8326 3803
rect 8360 3769 8394 3803
rect 8428 3769 8462 3803
rect 8496 3769 8530 3803
rect 8564 3769 8598 3803
rect 8632 3769 8666 3803
rect 8700 3769 8734 3803
rect 8768 3769 8802 3803
rect 8836 3769 8870 3803
rect 8904 3769 8938 3803
rect 8972 3769 9006 3803
rect 9148 3769 9182 3803
rect 9216 3769 9250 3803
rect 9284 3769 9318 3803
rect 9352 3769 9386 3803
rect 9420 3769 9454 3803
rect 9488 3769 9522 3803
rect 9556 3769 9590 3803
rect 9624 3769 9658 3803
rect 9692 3769 9726 3803
rect 9760 3769 9794 3803
rect 9828 3769 9862 3803
rect 10004 3769 10038 3803
rect 10072 3769 10106 3803
rect 10140 3769 10174 3803
rect 10208 3769 10242 3803
rect 10276 3769 10310 3803
rect 10344 3769 10378 3803
rect 10412 3769 10446 3803
rect 10480 3769 10514 3803
rect 10548 3769 10582 3803
rect 10616 3769 10650 3803
rect 10684 3769 10718 3803
<< ndiffres >>
rect 582 7806 3382 7906
rect 3484 7806 12884 7906
rect 582 7652 3382 7752
rect 3484 7652 12884 7752
rect 582 7498 3382 7598
rect 3484 7498 12884 7598
rect 582 7344 3382 7444
rect 3484 7344 12884 7444
rect 582 7190 3382 7290
rect 3484 7190 12884 7290
rect 582 7036 3382 7136
rect 3484 7036 12884 7136
rect 582 6882 3382 6982
rect 3484 6882 12884 6982
rect 582 6728 3382 6828
rect 3484 6728 12884 6828
rect 582 6574 3382 6674
rect 3484 6574 12884 6674
rect 582 6420 3382 6520
rect 3484 6420 12884 6520
rect 582 6266 3382 6366
rect 3484 6266 12884 6366
rect 582 6112 3382 6212
rect 3484 6112 12884 6212
rect 11728 5821 14528 5921
rect 11728 5667 14528 5767
rect 11728 5513 14528 5613
rect 11728 5359 14528 5459
rect 11728 5205 14528 5305
rect 11728 5051 14528 5151
rect 11728 4897 14528 4997
rect 11728 4743 14528 4843
rect 11728 4589 14528 4689
rect 11728 4435 14528 4535
rect 11728 4281 14528 4381
rect 11728 4127 14528 4227
rect 11728 3841 14528 3941
rect 11728 3687 14528 3787
rect 11728 3533 14528 3633
rect 11728 3379 14528 3479
rect 11728 3225 14528 3325
rect 11728 3071 14528 3171
rect 11728 2917 14528 3017
rect 11728 2763 14528 2863
rect 11728 2609 14528 2709
rect 11728 2455 14528 2555
rect 11728 2301 14528 2401
rect 11728 2147 14528 2247
rect 582 1857 3382 1957
rect 3484 1857 12884 1957
rect 582 1703 3382 1803
rect 3484 1703 12884 1803
rect 582 1549 3382 1649
rect 3484 1549 12884 1649
rect 582 1395 3382 1495
rect 3484 1395 12884 1495
rect 582 1241 3382 1341
rect 3484 1241 12884 1341
rect 582 1087 3382 1187
rect 3484 1087 12884 1187
rect 582 933 3382 1033
rect 3484 933 12884 1033
rect 582 779 3382 879
rect 3484 779 12884 879
rect 582 625 3382 725
rect 3484 625 12884 725
rect 582 471 3382 571
rect 3484 471 12884 571
rect 582 317 3382 417
rect 3484 317 12884 417
rect 582 163 3382 263
rect 3484 163 12884 263
<< locali >>
rect 344 8034 16033 8042
rect 336 8018 16033 8034
rect 370 8000 405 8018
rect 394 7984 405 8000
rect 439 7984 445 8018
rect 508 7984 517 8018
rect 577 7984 589 8018
rect 646 7984 661 8018
rect 715 7984 745 8018
rect 784 7984 819 8018
rect 853 7984 876 8018
rect 922 7984 948 8018
rect 991 7984 1020 8018
rect 1060 7984 1092 8018
rect 1129 7984 1164 8018
rect 1198 7984 1233 8018
rect 1270 7984 1302 8018
rect 1342 7984 1371 8018
rect 1414 7984 1440 8018
rect 1486 7984 1509 8018
rect 1558 7984 1578 8018
rect 1630 7984 1647 8018
rect 1702 7984 1716 8018
rect 1774 7984 1784 8018
rect 1846 7984 1852 8018
rect 1918 7984 1920 8018
rect 1954 7984 1956 8018
rect 2022 7984 2028 8018
rect 2090 7984 2100 8018
rect 2158 7984 2172 8018
rect 2226 7984 2244 8018
rect 2294 7984 2316 8018
rect 2362 7984 2388 8018
rect 2430 7984 2460 8018
rect 2498 7984 2532 8018
rect 2566 7984 2600 8018
rect 2638 7984 2668 8018
rect 2710 7984 2736 8018
rect 2782 7984 2804 8018
rect 2854 7984 2872 8018
rect 2926 7984 2940 8018
rect 2998 7984 3008 8018
rect 3070 7984 3076 8018
rect 3142 7984 3144 8018
rect 3178 7984 3180 8018
rect 3246 7984 3252 8018
rect 3314 7984 3324 8018
rect 3382 7984 3396 8018
rect 3450 7984 3468 8018
rect 3518 7984 3540 8018
rect 3586 7984 3612 8018
rect 3654 7984 3684 8018
rect 3722 7984 3756 8018
rect 3790 7984 3824 8018
rect 3862 7984 3892 8018
rect 3934 7984 3960 8018
rect 4006 7984 4028 8018
rect 4078 7984 4096 8018
rect 4150 7984 4164 8018
rect 4222 7984 4232 8018
rect 4294 7984 4300 8018
rect 4366 7984 4368 8018
rect 4402 7984 4404 8018
rect 4470 7984 4476 8018
rect 4538 7984 4572 8018
rect 4617 7984 4640 8018
rect 4691 7984 4708 8018
rect 4742 7984 4766 8018
rect 4810 7984 4838 8018
rect 4878 7984 4910 8018
rect 4946 7984 4980 8018
rect 5016 7984 5048 8018
rect 5088 7984 5116 8018
rect 5160 7984 5184 8018
rect 5232 7984 5252 8018
rect 5304 7984 5320 8018
rect 5376 7984 5388 8018
rect 5448 7984 5456 8018
rect 5520 7984 5524 8018
rect 5626 7984 5630 8018
rect 5694 7984 5702 8018
rect 5762 7984 5774 8018
rect 5830 7984 5846 8018
rect 5898 7984 5918 8018
rect 5966 7984 5990 8018
rect 6034 7984 6062 8018
rect 6102 7984 6134 8018
rect 6170 7984 6204 8018
rect 6240 7984 6272 8018
rect 6312 7984 6340 8018
rect 6384 7984 6408 8018
rect 6456 7984 6476 8018
rect 6528 7984 6544 8018
rect 6600 7984 6612 8018
rect 6646 7984 6667 8018
rect 6714 7984 6741 8018
rect 6782 7984 6816 8018
rect 6918 7984 6922 8018
rect 6986 7984 6994 8018
rect 7054 7984 7066 8018
rect 7122 7984 7138 8018
rect 7190 7984 7210 8018
rect 7258 7984 7282 8018
rect 7326 7984 7354 8018
rect 7394 7984 7426 8018
rect 7462 7984 7496 8018
rect 7532 7984 7564 8018
rect 7604 7984 7632 8018
rect 7676 7984 7700 8018
rect 7748 7984 7768 8018
rect 7820 7984 7836 8018
rect 7892 7984 7904 8018
rect 7964 7984 7972 8018
rect 8036 7984 8040 8018
rect 8142 7984 8146 8018
rect 8210 7984 8218 8018
rect 8278 7984 8290 8018
rect 8346 7984 8362 8018
rect 8414 7984 8434 8018
rect 8482 7984 8506 8018
rect 8550 7984 8578 8018
rect 8618 7984 8650 8018
rect 8686 7984 8720 8018
rect 8756 7984 8788 8018
rect 8828 7984 8856 8018
rect 8900 7984 8924 8018
rect 8972 7984 8992 8018
rect 9044 7984 9060 8018
rect 9116 7984 9128 8018
rect 9188 7984 9196 8018
rect 9260 7984 9264 8018
rect 9366 7984 9370 8018
rect 9434 7984 9442 8018
rect 9502 7984 9514 8018
rect 9570 7984 9586 8018
rect 9638 7984 9658 8018
rect 9706 7984 9730 8018
rect 9774 7984 9802 8018
rect 9842 7984 9874 8018
rect 9910 7984 9944 8018
rect 9980 7984 10012 8018
rect 10052 7984 10080 8018
rect 10124 7984 10148 8018
rect 10196 7984 10216 8018
rect 10268 7984 10284 8018
rect 10340 7984 10352 8018
rect 10412 7984 10420 8018
rect 10484 7984 10488 8018
rect 10590 7984 10594 8018
rect 10658 7984 10666 8018
rect 10726 7984 10738 8018
rect 10794 7984 10810 8018
rect 10862 7984 10882 8018
rect 10930 7984 10954 8018
rect 10998 7984 11026 8018
rect 11066 7984 11098 8018
rect 11134 7984 11168 8018
rect 11204 7984 11236 8018
rect 11276 7984 11304 8018
rect 11348 7984 11372 8018
rect 11420 7984 11440 8018
rect 11492 7984 11508 8018
rect 11564 7984 11576 8018
rect 11636 7984 11644 8018
rect 11708 7984 11712 8018
rect 11814 7984 11818 8018
rect 11882 7984 11890 8018
rect 11950 7984 11962 8018
rect 12018 7984 12034 8018
rect 12086 7984 12106 8018
rect 12154 7984 12178 8018
rect 12222 7984 12250 8018
rect 12290 7984 12322 8018
rect 12358 7984 12392 8018
rect 12428 7984 12460 8018
rect 12500 7984 12528 8018
rect 12572 7984 12596 8018
rect 12644 7984 12664 8018
rect 12716 7984 12732 8018
rect 12788 7984 12800 8018
rect 12860 7984 12868 8018
rect 12932 7984 12936 8018
rect 13038 7984 13042 8018
rect 13106 7984 13114 8018
rect 13174 7984 13186 8018
rect 13242 7984 13258 8018
rect 13310 7984 13330 8018
rect 13378 7984 13402 8018
rect 13446 7984 13474 8018
rect 13514 7984 13546 8018
rect 13582 7984 13616 8018
rect 13650 7984 13684 8018
rect 13718 7984 13752 8018
rect 13786 7984 13820 8018
rect 13854 7984 13888 8018
rect 13922 7984 13956 8018
rect 13990 7984 14024 8018
rect 14058 7984 14092 8018
rect 14126 7984 14160 8018
rect 14194 7984 14228 8018
rect 14262 7984 14296 8018
rect 14330 7984 14364 8018
rect 14398 7984 14432 8018
rect 14466 7984 14500 8018
rect 14534 7984 14568 8018
rect 14602 7984 14636 8018
rect 14670 7984 14774 8018
rect 14808 7984 14844 8018
rect 14878 7984 14914 8018
rect 14948 7984 14984 8018
rect 15018 7984 15054 8018
rect 15088 7984 15124 8018
rect 15158 7984 15194 8018
rect 15228 7984 15264 8018
rect 15298 7984 15334 8018
rect 15368 7984 15404 8018
rect 15438 7984 15474 8018
rect 15508 7984 15544 8018
rect 15578 7984 15614 8018
rect 15648 7984 15684 8018
rect 15718 8010 15754 8018
rect 15788 8010 15824 8018
rect 15718 7984 15733 8010
rect 15788 7984 15819 8010
rect 15858 7984 15894 8018
rect 15928 8010 15964 8018
rect 15998 8010 16033 8018
rect 15939 7984 15964 8010
rect 336 7968 360 7984
rect 344 7966 360 7968
rect 394 7976 15733 7984
rect 15767 7976 15819 7984
rect 15853 7976 15905 7984
rect 15939 7976 15991 7984
rect 16025 7976 16033 8010
rect 394 7966 16033 7976
rect 344 7960 16033 7966
rect 344 7928 410 7960
rect 344 7874 360 7928
rect 394 7874 410 7928
rect 13152 7949 16033 7960
rect 13152 7928 14774 7949
rect 13152 7894 13194 7928
rect 13228 7894 13264 7928
rect 13298 7894 13334 7928
rect 13368 7894 13404 7928
rect 13438 7894 13474 7928
rect 13508 7894 13544 7928
rect 13578 7894 13614 7928
rect 13648 7894 13684 7928
rect 13718 7894 13754 7928
rect 13788 7894 13824 7928
rect 13858 7894 13894 7928
rect 13928 7894 13964 7928
rect 13998 7894 14034 7928
rect 14068 7894 14104 7928
rect 14138 7894 14174 7928
rect 14208 7894 14244 7928
rect 14278 7894 14314 7928
rect 14348 7894 14384 7928
rect 14418 7894 14454 7928
rect 14488 7894 14524 7928
rect 14558 7894 14594 7928
rect 14628 7894 14664 7928
rect 14698 7915 14774 7928
rect 14808 7915 14844 7949
rect 14878 7915 14914 7949
rect 14948 7915 14984 7949
rect 15018 7915 15054 7949
rect 15088 7915 15124 7949
rect 15158 7915 15194 7949
rect 15228 7915 15264 7949
rect 15298 7915 15334 7949
rect 15368 7915 15404 7949
rect 15438 7915 15474 7949
rect 15508 7915 15544 7949
rect 15578 7915 15614 7949
rect 15648 7915 15684 7949
rect 15718 7938 15754 7949
rect 15788 7938 15824 7949
rect 15718 7915 15733 7938
rect 15788 7915 15819 7938
rect 15858 7915 15894 7949
rect 15928 7938 15964 7949
rect 15998 7938 16033 7949
rect 15939 7915 15964 7938
rect 14698 7904 15733 7915
rect 15767 7904 15819 7915
rect 15853 7904 15905 7915
rect 15939 7904 15991 7915
rect 16025 7904 16033 7938
rect 14698 7894 16033 7904
rect 344 7856 410 7874
rect 480 7873 582 7889
rect 3382 7873 3484 7889
rect 12884 7873 12986 7889
rect 13152 7880 16033 7894
rect 344 7804 360 7856
rect 394 7804 410 7856
rect 514 7839 548 7873
rect 3416 7839 3450 7873
rect 12918 7839 12952 7873
rect 13152 7858 14774 7880
rect 480 7823 582 7839
rect 3382 7823 3484 7839
rect 12884 7823 12986 7839
rect 13152 7824 13194 7858
rect 13228 7824 13264 7858
rect 13298 7824 13334 7858
rect 13368 7824 13404 7858
rect 13438 7824 13474 7858
rect 13508 7824 13544 7858
rect 13578 7824 13614 7858
rect 13648 7824 13684 7858
rect 13718 7824 13754 7858
rect 13788 7824 13824 7858
rect 13858 7824 13894 7858
rect 13928 7824 13964 7858
rect 13998 7824 14034 7858
rect 14068 7824 14104 7858
rect 14138 7824 14174 7858
rect 14208 7824 14244 7858
rect 14278 7824 14314 7858
rect 14348 7824 14384 7858
rect 14418 7824 14454 7858
rect 14488 7824 14524 7858
rect 14558 7824 14594 7858
rect 14628 7824 14664 7858
rect 14698 7846 14774 7858
rect 14808 7846 14844 7880
rect 14878 7846 14914 7880
rect 14948 7846 14984 7880
rect 15018 7846 15054 7880
rect 15088 7846 15124 7880
rect 15158 7846 15194 7880
rect 15228 7846 15264 7880
rect 15298 7846 15334 7880
rect 15368 7846 15404 7880
rect 15438 7846 15474 7880
rect 15508 7846 15544 7880
rect 15578 7846 15614 7880
rect 15648 7846 15684 7880
rect 15718 7866 15754 7880
rect 15788 7866 15824 7880
rect 15718 7846 15733 7866
rect 15788 7846 15819 7866
rect 15858 7846 15894 7880
rect 15928 7866 15964 7880
rect 15998 7866 16033 7880
rect 15939 7846 15964 7866
rect 14698 7832 15733 7846
rect 15767 7832 15819 7846
rect 15853 7832 15905 7846
rect 15939 7832 15991 7846
rect 16025 7832 16033 7866
rect 14698 7824 16033 7832
rect 344 7784 410 7804
rect 344 7734 360 7784
rect 394 7734 410 7784
rect 13152 7811 16033 7824
rect 13152 7788 14774 7811
rect 13152 7754 13194 7788
rect 13228 7754 13264 7788
rect 13298 7754 13334 7788
rect 13368 7754 13404 7788
rect 13438 7754 13474 7788
rect 13508 7754 13544 7788
rect 13578 7754 13614 7788
rect 13648 7754 13684 7788
rect 13718 7754 13754 7788
rect 13788 7754 13824 7788
rect 13858 7754 13894 7788
rect 13928 7754 13964 7788
rect 13998 7754 14034 7788
rect 14068 7754 14104 7788
rect 14138 7754 14174 7788
rect 14208 7754 14244 7788
rect 14278 7754 14314 7788
rect 14348 7754 14384 7788
rect 14418 7754 14454 7788
rect 14488 7754 14524 7788
rect 14558 7754 14594 7788
rect 14628 7754 14664 7788
rect 14698 7777 14774 7788
rect 14808 7777 14844 7811
rect 14878 7777 14914 7811
rect 14948 7777 14984 7811
rect 15018 7777 15054 7811
rect 15088 7777 15124 7811
rect 15158 7777 15194 7811
rect 15228 7777 15264 7811
rect 15298 7777 15334 7811
rect 15368 7777 15404 7811
rect 15438 7777 15474 7811
rect 15508 7777 15544 7811
rect 15578 7777 15614 7811
rect 15648 7777 15684 7811
rect 15718 7794 15754 7811
rect 15788 7794 15824 7811
rect 15718 7777 15733 7794
rect 15788 7777 15819 7794
rect 15858 7777 15894 7811
rect 15928 7794 15964 7811
rect 15998 7794 16033 7811
rect 15939 7777 15964 7794
rect 14698 7760 15733 7777
rect 15767 7760 15819 7777
rect 15853 7760 15905 7777
rect 15939 7760 15991 7777
rect 16025 7760 16033 7794
rect 14698 7754 16033 7760
rect 13152 7742 16033 7754
rect 344 7712 410 7734
rect 480 7719 582 7735
rect 3382 7719 3484 7735
rect 12884 7719 12986 7735
rect 344 7664 360 7712
rect 394 7664 410 7712
rect 514 7685 548 7719
rect 3416 7685 3450 7719
rect 12918 7685 12952 7719
rect 13152 7718 14774 7742
rect 480 7669 582 7685
rect 3382 7669 3484 7685
rect 12884 7669 12986 7685
rect 13152 7684 13194 7718
rect 13228 7684 13264 7718
rect 13298 7684 13334 7718
rect 13368 7684 13404 7718
rect 13438 7684 13474 7718
rect 13508 7684 13544 7718
rect 13578 7684 13614 7718
rect 13648 7684 13684 7718
rect 13718 7684 13754 7718
rect 13788 7684 13824 7718
rect 13858 7684 13894 7718
rect 13928 7684 13964 7718
rect 13998 7684 14034 7718
rect 14068 7684 14104 7718
rect 14138 7684 14174 7718
rect 14208 7684 14244 7718
rect 14278 7684 14314 7718
rect 14348 7684 14384 7718
rect 14418 7684 14454 7718
rect 14488 7684 14524 7718
rect 14558 7684 14594 7718
rect 14628 7684 14664 7718
rect 14698 7708 14774 7718
rect 14808 7708 14844 7742
rect 14878 7708 14914 7742
rect 14948 7708 14984 7742
rect 15018 7708 15054 7742
rect 15088 7708 15124 7742
rect 15158 7708 15194 7742
rect 15228 7708 15264 7742
rect 15298 7708 15334 7742
rect 15368 7708 15404 7742
rect 15438 7708 15474 7742
rect 15508 7708 15544 7742
rect 15578 7708 15614 7742
rect 15648 7708 15684 7742
rect 15718 7722 15754 7742
rect 15788 7722 15824 7742
rect 15718 7708 15733 7722
rect 15788 7708 15819 7722
rect 15858 7708 15894 7742
rect 15928 7722 15964 7742
rect 15998 7722 16033 7742
rect 15939 7708 15964 7722
rect 14698 7688 15733 7708
rect 15767 7688 15819 7708
rect 15853 7688 15905 7708
rect 15939 7688 15991 7708
rect 16025 7688 16033 7722
rect 14698 7684 16033 7688
rect 13152 7673 16033 7684
rect 344 7640 410 7664
rect 344 7594 360 7640
rect 394 7594 410 7640
rect 344 7568 410 7594
rect 13152 7648 14774 7673
rect 13152 7614 13194 7648
rect 13228 7614 13264 7648
rect 13298 7614 13334 7648
rect 13368 7614 13404 7648
rect 13438 7614 13474 7648
rect 13508 7614 13544 7648
rect 13578 7614 13614 7648
rect 13648 7614 13684 7648
rect 13718 7614 13754 7648
rect 13788 7614 13824 7648
rect 13858 7614 13894 7648
rect 13928 7614 13964 7648
rect 13998 7614 14034 7648
rect 14068 7614 14104 7648
rect 14138 7614 14174 7648
rect 14208 7614 14244 7648
rect 14278 7614 14314 7648
rect 14348 7614 14384 7648
rect 14418 7614 14454 7648
rect 14488 7614 14524 7648
rect 14558 7614 14594 7648
rect 14628 7614 14664 7648
rect 14698 7639 14774 7648
rect 14808 7639 14844 7673
rect 14878 7639 14914 7673
rect 14948 7639 14984 7673
rect 15018 7639 15054 7673
rect 15088 7639 15124 7673
rect 15158 7639 15194 7673
rect 15228 7639 15264 7673
rect 15298 7639 15334 7673
rect 15368 7639 15404 7673
rect 15438 7639 15474 7673
rect 15508 7639 15544 7673
rect 15578 7639 15614 7673
rect 15648 7639 15684 7673
rect 15718 7650 15754 7673
rect 15788 7650 15824 7673
rect 15718 7639 15733 7650
rect 15788 7639 15819 7650
rect 15858 7639 15894 7673
rect 15928 7650 15964 7673
rect 15998 7650 16033 7673
rect 15939 7639 15964 7650
rect 14698 7616 15733 7639
rect 15767 7616 15819 7639
rect 15853 7616 15905 7639
rect 15939 7616 15991 7639
rect 16025 7616 16033 7650
rect 14698 7614 16033 7616
rect 13152 7604 16033 7614
rect 344 7524 360 7568
rect 394 7524 410 7568
rect 480 7565 582 7581
rect 3382 7565 3484 7581
rect 12884 7565 12986 7581
rect 13152 7578 14774 7604
rect 514 7531 548 7565
rect 3416 7531 3450 7565
rect 12918 7531 12952 7565
rect 13152 7544 13194 7578
rect 13228 7544 13264 7578
rect 13298 7544 13334 7578
rect 13368 7544 13404 7578
rect 13438 7544 13474 7578
rect 13508 7544 13544 7578
rect 13578 7544 13614 7578
rect 13648 7544 13684 7578
rect 13718 7544 13754 7578
rect 13788 7544 13824 7578
rect 13858 7544 13894 7578
rect 13928 7544 13964 7578
rect 13998 7544 14034 7578
rect 14068 7544 14104 7578
rect 14138 7544 14174 7578
rect 14208 7544 14244 7578
rect 14278 7544 14314 7578
rect 14348 7544 14384 7578
rect 14418 7544 14454 7578
rect 14488 7544 14524 7578
rect 14558 7544 14594 7578
rect 14628 7544 14664 7578
rect 14698 7570 14774 7578
rect 14808 7570 14844 7604
rect 14878 7570 14914 7604
rect 14948 7570 14984 7604
rect 15018 7570 15054 7604
rect 15088 7570 15124 7604
rect 15158 7570 15194 7604
rect 15228 7570 15264 7604
rect 15298 7570 15334 7604
rect 15368 7570 15404 7604
rect 15438 7570 15474 7604
rect 15508 7570 15544 7604
rect 15578 7570 15614 7604
rect 15648 7570 15684 7604
rect 15718 7578 15754 7604
rect 15788 7578 15824 7604
rect 15718 7570 15733 7578
rect 15788 7570 15819 7578
rect 15858 7570 15894 7604
rect 15928 7578 15964 7604
rect 15998 7578 16033 7604
rect 15939 7570 15964 7578
rect 14698 7544 15733 7570
rect 15767 7544 15819 7570
rect 15853 7544 15905 7570
rect 15939 7544 15991 7570
rect 16025 7544 16033 7578
rect 13152 7535 16033 7544
rect 344 7496 410 7524
rect 480 7515 582 7531
rect 3382 7515 3484 7531
rect 12884 7515 12986 7531
rect 344 7454 360 7496
rect 394 7454 410 7496
rect 344 7424 410 7454
rect 13152 7508 14774 7535
rect 13152 7474 13194 7508
rect 13228 7474 13264 7508
rect 13298 7474 13334 7508
rect 13368 7474 13404 7508
rect 13438 7474 13474 7508
rect 13508 7474 13544 7508
rect 13578 7474 13614 7508
rect 13648 7474 13684 7508
rect 13718 7474 13754 7508
rect 13788 7474 13824 7508
rect 13858 7474 13894 7508
rect 13928 7474 13964 7508
rect 13998 7474 14034 7508
rect 14068 7474 14104 7508
rect 14138 7474 14174 7508
rect 14208 7474 14244 7508
rect 14278 7474 14314 7508
rect 14348 7474 14384 7508
rect 14418 7474 14454 7508
rect 14488 7474 14524 7508
rect 14558 7474 14594 7508
rect 14628 7474 14664 7508
rect 14698 7501 14774 7508
rect 14808 7501 14844 7535
rect 14878 7501 14914 7535
rect 14948 7501 14984 7535
rect 15018 7501 15054 7535
rect 15088 7501 15124 7535
rect 15158 7501 15194 7535
rect 15228 7501 15264 7535
rect 15298 7501 15334 7535
rect 15368 7501 15404 7535
rect 15438 7501 15474 7535
rect 15508 7501 15544 7535
rect 15578 7501 15614 7535
rect 15648 7501 15684 7535
rect 15718 7506 15754 7535
rect 15788 7506 15824 7535
rect 15718 7501 15733 7506
rect 15788 7501 15819 7506
rect 15858 7501 15894 7535
rect 15928 7506 15964 7535
rect 15998 7506 16033 7535
rect 15939 7501 15964 7506
rect 14698 7474 15733 7501
rect 13152 7472 15733 7474
rect 15767 7472 15819 7501
rect 15853 7472 15905 7501
rect 15939 7472 15991 7501
rect 16025 7472 16033 7506
rect 13152 7466 16033 7472
rect 13152 7438 14774 7466
rect 344 7384 360 7424
rect 394 7384 410 7424
rect 480 7411 582 7427
rect 3382 7411 3484 7427
rect 12884 7411 12986 7427
rect 344 7352 410 7384
rect 514 7377 548 7411
rect 3416 7377 3450 7411
rect 12918 7377 12952 7411
rect 13152 7404 13194 7438
rect 13228 7404 13264 7438
rect 13298 7404 13334 7438
rect 13368 7404 13404 7438
rect 13438 7404 13474 7438
rect 13508 7404 13544 7438
rect 13578 7404 13614 7438
rect 13648 7404 13684 7438
rect 13718 7404 13754 7438
rect 13788 7404 13824 7438
rect 13858 7404 13894 7438
rect 13928 7404 13964 7438
rect 13998 7404 14034 7438
rect 14068 7404 14104 7438
rect 14138 7404 14174 7438
rect 14208 7404 14244 7438
rect 14278 7404 14314 7438
rect 14348 7404 14384 7438
rect 14418 7404 14454 7438
rect 14488 7404 14524 7438
rect 14558 7404 14594 7438
rect 14628 7404 14664 7438
rect 14698 7432 14774 7438
rect 14808 7432 14844 7466
rect 14878 7432 14914 7466
rect 14948 7432 14984 7466
rect 15018 7432 15054 7466
rect 15088 7432 15124 7466
rect 15158 7432 15194 7466
rect 15228 7432 15264 7466
rect 15298 7432 15334 7466
rect 15368 7432 15404 7466
rect 15438 7432 15474 7466
rect 15508 7432 15544 7466
rect 15578 7432 15614 7466
rect 15648 7432 15684 7466
rect 15718 7434 15754 7466
rect 15788 7434 15824 7466
rect 15718 7432 15733 7434
rect 15788 7432 15819 7434
rect 15858 7432 15894 7466
rect 15928 7434 15964 7466
rect 15998 7434 16033 7466
rect 15939 7432 15964 7434
rect 14698 7404 15733 7432
rect 13152 7400 15733 7404
rect 15767 7400 15819 7432
rect 15853 7400 15905 7432
rect 15939 7400 15991 7432
rect 16025 7400 16033 7434
rect 13152 7397 16033 7400
rect 480 7361 582 7377
rect 3382 7361 3484 7377
rect 12884 7361 12986 7377
rect 13152 7368 14774 7397
rect 344 7314 360 7352
rect 394 7314 410 7352
rect 344 7280 410 7314
rect 344 7244 360 7280
rect 394 7244 410 7280
rect 13152 7334 13194 7368
rect 13228 7334 13264 7368
rect 13298 7334 13334 7368
rect 13368 7334 13404 7368
rect 13438 7334 13474 7368
rect 13508 7334 13544 7368
rect 13578 7334 13614 7368
rect 13648 7334 13684 7368
rect 13718 7334 13754 7368
rect 13788 7334 13824 7368
rect 13858 7334 13894 7368
rect 13928 7334 13964 7368
rect 13998 7334 14034 7368
rect 14068 7334 14104 7368
rect 14138 7334 14174 7368
rect 14208 7334 14244 7368
rect 14278 7334 14314 7368
rect 14348 7334 14384 7368
rect 14418 7334 14454 7368
rect 14488 7334 14524 7368
rect 14558 7334 14594 7368
rect 14628 7334 14664 7368
rect 14698 7363 14774 7368
rect 14808 7363 14844 7397
rect 14878 7363 14914 7397
rect 14948 7363 14984 7397
rect 15018 7363 15054 7397
rect 15088 7363 15124 7397
rect 15158 7363 15194 7397
rect 15228 7363 15264 7397
rect 15298 7363 15334 7397
rect 15368 7363 15404 7397
rect 15438 7363 15474 7397
rect 15508 7363 15544 7397
rect 15578 7363 15614 7397
rect 15648 7363 15684 7397
rect 15718 7363 15754 7397
rect 15788 7363 15824 7397
rect 15858 7363 15894 7397
rect 15928 7363 15964 7397
rect 15998 7363 16033 7397
rect 14698 7362 16033 7363
rect 14698 7334 15733 7362
rect 13152 7328 15733 7334
rect 15767 7328 15819 7362
rect 15853 7328 15905 7362
rect 15939 7328 15991 7362
rect 16025 7328 16033 7362
rect 13152 7298 14774 7328
rect 480 7257 582 7273
rect 3382 7257 3484 7273
rect 12884 7257 12986 7273
rect 13152 7264 13194 7298
rect 13228 7264 13264 7298
rect 13298 7264 13334 7298
rect 13368 7264 13404 7298
rect 13438 7264 13474 7298
rect 13508 7264 13544 7298
rect 13578 7264 13614 7298
rect 13648 7264 13684 7298
rect 13718 7264 13754 7298
rect 13788 7264 13824 7298
rect 13858 7264 13894 7298
rect 13928 7264 13964 7298
rect 13998 7264 14034 7298
rect 14068 7264 14104 7298
rect 14138 7264 14174 7298
rect 14208 7264 14244 7298
rect 14278 7264 14314 7298
rect 14348 7264 14384 7298
rect 14418 7264 14454 7298
rect 14488 7264 14524 7298
rect 14558 7264 14594 7298
rect 14628 7264 14664 7298
rect 14698 7294 14774 7298
rect 14808 7294 14844 7328
rect 14878 7294 14914 7328
rect 14948 7294 14984 7328
rect 15018 7294 15054 7328
rect 15088 7294 15124 7328
rect 15158 7294 15194 7328
rect 15228 7294 15264 7328
rect 15298 7294 15334 7328
rect 15368 7294 15404 7328
rect 15438 7294 15474 7328
rect 15508 7294 15544 7328
rect 15578 7294 15614 7328
rect 15648 7294 15684 7328
rect 15718 7294 15754 7328
rect 15788 7294 15824 7328
rect 15858 7294 15894 7328
rect 15928 7294 15964 7328
rect 15998 7294 16033 7328
rect 14698 7290 16033 7294
rect 14698 7264 15733 7290
rect 13152 7259 15733 7264
rect 15767 7259 15819 7290
rect 15853 7259 15905 7290
rect 15939 7259 15991 7290
rect 344 7208 410 7244
rect 514 7223 548 7257
rect 3416 7223 3450 7257
rect 12918 7223 12952 7257
rect 13152 7228 14774 7259
rect 344 7174 360 7208
rect 394 7174 410 7208
rect 480 7207 582 7223
rect 3382 7207 3484 7223
rect 12884 7207 12986 7223
rect 344 7138 410 7174
rect 344 7102 360 7138
rect 394 7102 410 7138
rect 13152 7194 13194 7228
rect 13228 7194 13264 7228
rect 13298 7194 13334 7228
rect 13368 7194 13404 7228
rect 13438 7194 13474 7228
rect 13508 7194 13544 7228
rect 13578 7194 13614 7228
rect 13648 7194 13684 7228
rect 13718 7194 13754 7228
rect 13788 7194 13824 7228
rect 13858 7194 13894 7228
rect 13928 7194 13964 7228
rect 13998 7194 14034 7228
rect 14068 7194 14104 7228
rect 14138 7194 14174 7228
rect 14208 7194 14244 7228
rect 14278 7194 14314 7228
rect 14348 7194 14384 7228
rect 14418 7194 14454 7228
rect 14488 7194 14524 7228
rect 14558 7194 14594 7228
rect 14628 7194 14664 7228
rect 14698 7225 14774 7228
rect 14808 7225 14844 7259
rect 14878 7225 14914 7259
rect 14948 7225 14984 7259
rect 15018 7225 15054 7259
rect 15088 7225 15124 7259
rect 15158 7225 15194 7259
rect 15228 7225 15264 7259
rect 15298 7225 15334 7259
rect 15368 7225 15404 7259
rect 15438 7225 15474 7259
rect 15508 7225 15544 7259
rect 15578 7225 15614 7259
rect 15648 7225 15684 7259
rect 15718 7256 15733 7259
rect 15788 7256 15819 7259
rect 15718 7225 15754 7256
rect 15788 7225 15824 7256
rect 15858 7225 15894 7259
rect 15939 7256 15964 7259
rect 16025 7256 16033 7290
rect 15928 7225 15964 7256
rect 15998 7225 16033 7256
rect 14698 7218 16033 7225
rect 14698 7194 15733 7218
rect 13152 7190 15733 7194
rect 15767 7190 15819 7218
rect 15853 7190 15905 7218
rect 15939 7190 15991 7218
rect 13152 7158 14774 7190
rect 13152 7124 13194 7158
rect 13228 7124 13264 7158
rect 13298 7124 13334 7158
rect 13368 7124 13404 7158
rect 13438 7124 13474 7158
rect 13508 7124 13544 7158
rect 13578 7124 13614 7158
rect 13648 7124 13684 7158
rect 13718 7124 13754 7158
rect 13788 7124 13824 7158
rect 13858 7124 13894 7158
rect 13928 7124 13964 7158
rect 13998 7124 14034 7158
rect 14068 7124 14104 7158
rect 14138 7124 14174 7158
rect 14208 7124 14244 7158
rect 14278 7124 14314 7158
rect 14348 7124 14384 7158
rect 14418 7124 14454 7158
rect 14488 7124 14524 7158
rect 14558 7124 14594 7158
rect 14628 7124 14664 7158
rect 14698 7156 14774 7158
rect 14808 7156 14844 7190
rect 14878 7156 14914 7190
rect 14948 7156 14984 7190
rect 15018 7156 15054 7190
rect 15088 7156 15124 7190
rect 15158 7156 15194 7190
rect 15228 7156 15264 7190
rect 15298 7156 15334 7190
rect 15368 7156 15404 7190
rect 15438 7156 15474 7190
rect 15508 7156 15544 7190
rect 15578 7156 15614 7190
rect 15648 7156 15684 7190
rect 15718 7184 15733 7190
rect 15788 7184 15819 7190
rect 15718 7156 15754 7184
rect 15788 7156 15824 7184
rect 15858 7156 15894 7190
rect 15939 7184 15964 7190
rect 16025 7184 16033 7218
rect 15928 7156 15964 7184
rect 15998 7156 16033 7184
rect 14698 7146 16033 7156
rect 14698 7124 15733 7146
rect 13152 7121 15733 7124
rect 15767 7121 15819 7146
rect 15853 7121 15905 7146
rect 15939 7121 15991 7146
rect 480 7103 582 7119
rect 3382 7103 3484 7119
rect 12884 7103 12986 7119
rect 344 7068 410 7102
rect 514 7069 548 7103
rect 3416 7069 3450 7103
rect 12918 7069 12952 7103
rect 13152 7088 14774 7121
rect 344 7030 360 7068
rect 394 7030 410 7068
rect 480 7053 582 7069
rect 3382 7053 3484 7069
rect 12884 7053 12986 7069
rect 13152 7054 13194 7088
rect 13228 7054 13264 7088
rect 13298 7054 13334 7088
rect 13368 7054 13404 7088
rect 13438 7054 13474 7088
rect 13508 7054 13544 7088
rect 13578 7054 13614 7088
rect 13648 7054 13684 7088
rect 13718 7054 13754 7088
rect 13788 7054 13824 7088
rect 13858 7054 13894 7088
rect 13928 7054 13964 7088
rect 13998 7054 14034 7088
rect 14068 7054 14104 7088
rect 14138 7054 14174 7088
rect 14208 7054 14244 7088
rect 14278 7054 14314 7088
rect 14348 7054 14384 7088
rect 14418 7054 14454 7088
rect 14488 7054 14524 7088
rect 14558 7054 14594 7088
rect 14628 7054 14664 7088
rect 14698 7087 14774 7088
rect 14808 7087 14844 7121
rect 14878 7087 14914 7121
rect 14948 7087 14984 7121
rect 15018 7087 15054 7121
rect 15088 7087 15124 7121
rect 15158 7087 15194 7121
rect 15228 7087 15264 7121
rect 15298 7087 15334 7121
rect 15368 7087 15404 7121
rect 15438 7087 15474 7121
rect 15508 7087 15544 7121
rect 15578 7087 15614 7121
rect 15648 7087 15684 7121
rect 15718 7112 15733 7121
rect 15788 7112 15819 7121
rect 15718 7087 15754 7112
rect 15788 7087 15824 7112
rect 15858 7087 15894 7121
rect 15939 7112 15964 7121
rect 16025 7112 16033 7146
rect 15928 7087 15964 7112
rect 15998 7087 16033 7112
rect 14698 7074 16033 7087
rect 14698 7054 15733 7074
rect 344 6999 410 7030
rect 344 6958 360 6999
rect 394 6958 410 6999
rect 13152 7052 15733 7054
rect 15767 7052 15819 7074
rect 15853 7052 15905 7074
rect 15939 7052 15991 7074
rect 13152 7018 14774 7052
rect 14808 7018 14844 7052
rect 14878 7018 14914 7052
rect 14948 7018 14984 7052
rect 15018 7018 15054 7052
rect 15088 7018 15124 7052
rect 15158 7018 15194 7052
rect 15228 7018 15264 7052
rect 15298 7018 15334 7052
rect 15368 7018 15404 7052
rect 15438 7018 15474 7052
rect 15508 7018 15544 7052
rect 15578 7018 15614 7052
rect 15648 7018 15684 7052
rect 15718 7040 15733 7052
rect 15788 7040 15819 7052
rect 15718 7018 15754 7040
rect 15788 7018 15824 7040
rect 15858 7018 15894 7052
rect 15939 7040 15964 7052
rect 16025 7040 16033 7074
rect 15928 7018 15964 7040
rect 15998 7018 16033 7040
rect 13152 6984 13194 7018
rect 13228 6984 13264 7018
rect 13298 6984 13334 7018
rect 13368 6984 13404 7018
rect 13438 6984 13474 7018
rect 13508 6984 13544 7018
rect 13578 6984 13614 7018
rect 13648 6984 13684 7018
rect 13718 6984 13754 7018
rect 13788 6984 13824 7018
rect 13858 6984 13894 7018
rect 13928 6984 13964 7018
rect 13998 6984 14034 7018
rect 14068 6984 14104 7018
rect 14138 6984 14174 7018
rect 14208 6984 14244 7018
rect 14278 6984 14314 7018
rect 14348 6984 14384 7018
rect 14418 6984 14454 7018
rect 14488 6984 14524 7018
rect 14558 6984 14594 7018
rect 14628 6984 14664 7018
rect 14698 7002 16033 7018
rect 14698 6984 15733 7002
rect 13152 6983 15733 6984
rect 15767 6983 15819 7002
rect 15853 6983 15905 7002
rect 15939 6983 15991 7002
rect 344 6930 410 6958
rect 480 6949 582 6965
rect 3382 6949 3484 6965
rect 12884 6949 12986 6965
rect 13152 6949 14774 6983
rect 14808 6949 14844 6983
rect 14878 6949 14914 6983
rect 14948 6949 14984 6983
rect 15018 6949 15054 6983
rect 15088 6949 15124 6983
rect 15158 6949 15194 6983
rect 15228 6949 15264 6983
rect 15298 6949 15334 6983
rect 15368 6949 15404 6983
rect 15438 6949 15474 6983
rect 15508 6949 15544 6983
rect 15578 6949 15614 6983
rect 15648 6949 15684 6983
rect 15718 6968 15733 6983
rect 15788 6968 15819 6983
rect 15718 6949 15754 6968
rect 15788 6949 15824 6968
rect 15858 6949 15894 6983
rect 15939 6968 15964 6983
rect 16025 6968 16033 7002
rect 15928 6949 15964 6968
rect 15998 6949 16033 6968
rect 344 6886 360 6930
rect 394 6886 410 6930
rect 514 6915 548 6949
rect 3416 6915 3450 6949
rect 12918 6915 12952 6949
rect 13152 6948 16033 6949
rect 480 6899 582 6915
rect 3382 6899 3484 6915
rect 12884 6899 12986 6915
rect 13152 6914 13194 6948
rect 13228 6914 13264 6948
rect 13298 6914 13334 6948
rect 13368 6914 13404 6948
rect 13438 6914 13474 6948
rect 13508 6914 13544 6948
rect 13578 6914 13614 6948
rect 13648 6914 13684 6948
rect 13718 6914 13754 6948
rect 13788 6914 13824 6948
rect 13858 6914 13894 6948
rect 13928 6914 13964 6948
rect 13998 6914 14034 6948
rect 14068 6914 14104 6948
rect 14138 6914 14174 6948
rect 14208 6914 14244 6948
rect 14278 6914 14314 6948
rect 14348 6914 14384 6948
rect 14418 6914 14454 6948
rect 14488 6914 14524 6948
rect 14558 6914 14594 6948
rect 14628 6914 14664 6948
rect 14698 6930 16033 6948
rect 14698 6914 15733 6930
rect 15767 6914 15819 6930
rect 15853 6914 15905 6930
rect 15939 6914 15991 6930
rect 344 6861 410 6886
rect 344 6814 360 6861
rect 394 6814 410 6861
rect 344 6792 410 6814
rect 13152 6880 14774 6914
rect 14808 6880 14844 6914
rect 14878 6880 14914 6914
rect 14948 6880 14984 6914
rect 15018 6880 15054 6914
rect 15088 6880 15124 6914
rect 15158 6880 15194 6914
rect 15228 6880 15264 6914
rect 15298 6880 15334 6914
rect 15368 6880 15404 6914
rect 15438 6880 15474 6914
rect 15508 6880 15544 6914
rect 15578 6880 15614 6914
rect 15648 6880 15684 6914
rect 15718 6896 15733 6914
rect 15788 6896 15819 6914
rect 15718 6880 15754 6896
rect 15788 6880 15824 6896
rect 15858 6880 15894 6914
rect 15939 6896 15964 6914
rect 16025 6896 16033 6930
rect 15928 6880 15964 6896
rect 15998 6880 16033 6896
rect 13152 6878 16033 6880
rect 13152 6844 13194 6878
rect 13228 6844 13264 6878
rect 13298 6844 13334 6878
rect 13368 6844 13404 6878
rect 13438 6844 13474 6878
rect 13508 6844 13544 6878
rect 13578 6844 13614 6878
rect 13648 6844 13684 6878
rect 13718 6844 13754 6878
rect 13788 6844 13824 6878
rect 13858 6844 13894 6878
rect 13928 6844 13964 6878
rect 13998 6844 14034 6878
rect 14068 6844 14104 6878
rect 14138 6844 14174 6878
rect 14208 6844 14244 6878
rect 14278 6844 14314 6878
rect 14348 6844 14384 6878
rect 14418 6844 14454 6878
rect 14488 6844 14524 6878
rect 14558 6844 14594 6878
rect 14628 6844 14664 6878
rect 14698 6858 16033 6878
rect 14698 6845 15733 6858
rect 15767 6845 15819 6858
rect 15853 6845 15905 6858
rect 15939 6845 15991 6858
rect 14698 6844 14774 6845
rect 13152 6811 14774 6844
rect 14808 6811 14844 6845
rect 14878 6811 14914 6845
rect 14948 6811 14984 6845
rect 15018 6811 15054 6845
rect 15088 6811 15124 6845
rect 15158 6811 15194 6845
rect 15228 6811 15264 6845
rect 15298 6811 15334 6845
rect 15368 6811 15404 6845
rect 15438 6811 15474 6845
rect 15508 6811 15544 6845
rect 15578 6811 15614 6845
rect 15648 6811 15684 6845
rect 15718 6824 15733 6845
rect 15788 6824 15819 6845
rect 15718 6811 15754 6824
rect 15788 6811 15824 6824
rect 15858 6811 15894 6845
rect 15939 6824 15964 6845
rect 16025 6824 16033 6858
rect 15928 6811 15964 6824
rect 15998 6811 16033 6824
rect 480 6795 582 6811
rect 3382 6795 3484 6811
rect 12884 6795 12986 6811
rect 13152 6808 16033 6811
rect 344 6742 360 6792
rect 394 6742 410 6792
rect 514 6761 548 6795
rect 3416 6761 3450 6795
rect 12918 6761 12952 6795
rect 13152 6774 13194 6808
rect 13228 6774 13264 6808
rect 13298 6774 13334 6808
rect 13368 6774 13404 6808
rect 13438 6774 13474 6808
rect 13508 6774 13544 6808
rect 13578 6774 13614 6808
rect 13648 6774 13684 6808
rect 13718 6774 13754 6808
rect 13788 6774 13824 6808
rect 13858 6774 13894 6808
rect 13928 6774 13964 6808
rect 13998 6774 14034 6808
rect 14068 6774 14104 6808
rect 14138 6774 14174 6808
rect 14208 6774 14244 6808
rect 14278 6774 14314 6808
rect 14348 6774 14384 6808
rect 14418 6774 14454 6808
rect 14488 6774 14524 6808
rect 14558 6774 14594 6808
rect 14628 6774 14664 6808
rect 14698 6786 16033 6808
rect 14698 6776 15733 6786
rect 15767 6776 15819 6786
rect 15853 6776 15905 6786
rect 15939 6776 15991 6786
rect 14698 6774 14774 6776
rect 480 6745 582 6761
rect 3382 6745 3484 6761
rect 12884 6745 12986 6761
rect 344 6723 410 6742
rect 344 6670 360 6723
rect 394 6670 410 6723
rect 344 6654 410 6670
rect 13152 6742 14774 6774
rect 14808 6742 14844 6776
rect 14878 6742 14914 6776
rect 14948 6742 14984 6776
rect 15018 6742 15054 6776
rect 15088 6742 15124 6776
rect 15158 6742 15194 6776
rect 15228 6742 15264 6776
rect 15298 6742 15334 6776
rect 15368 6742 15404 6776
rect 15438 6742 15474 6776
rect 15508 6742 15544 6776
rect 15578 6742 15614 6776
rect 15648 6742 15684 6776
rect 15718 6752 15733 6776
rect 15788 6752 15819 6776
rect 15718 6742 15754 6752
rect 15788 6742 15824 6752
rect 15858 6742 15894 6776
rect 15939 6752 15964 6776
rect 16025 6752 16033 6786
rect 15928 6742 15964 6752
rect 15998 6742 16033 6752
rect 13152 6738 16033 6742
rect 13152 6704 13194 6738
rect 13228 6704 13264 6738
rect 13298 6704 13334 6738
rect 13368 6704 13404 6738
rect 13438 6704 13474 6738
rect 13508 6704 13544 6738
rect 13578 6704 13614 6738
rect 13648 6704 13684 6738
rect 13718 6704 13754 6738
rect 13788 6704 13824 6738
rect 13858 6704 13894 6738
rect 13928 6704 13964 6738
rect 13998 6704 14034 6738
rect 14068 6704 14104 6738
rect 14138 6704 14174 6738
rect 14208 6704 14244 6738
rect 14278 6704 14314 6738
rect 14348 6704 14384 6738
rect 14418 6704 14454 6738
rect 14488 6704 14524 6738
rect 14558 6704 14594 6738
rect 14628 6704 14664 6738
rect 14698 6714 16033 6738
rect 14698 6707 15733 6714
rect 15767 6707 15819 6714
rect 15853 6707 15905 6714
rect 15939 6707 15991 6714
rect 14698 6704 14774 6707
rect 13152 6673 14774 6704
rect 14808 6673 14844 6707
rect 14878 6673 14914 6707
rect 14948 6673 14984 6707
rect 15018 6673 15054 6707
rect 15088 6673 15124 6707
rect 15158 6673 15194 6707
rect 15228 6673 15264 6707
rect 15298 6673 15334 6707
rect 15368 6673 15404 6707
rect 15438 6673 15474 6707
rect 15508 6673 15544 6707
rect 15578 6673 15614 6707
rect 15648 6673 15684 6707
rect 15718 6680 15733 6707
rect 15788 6680 15819 6707
rect 15718 6673 15754 6680
rect 15788 6673 15824 6680
rect 15858 6673 15894 6707
rect 15939 6680 15964 6707
rect 16025 6680 16033 6714
rect 15928 6673 15964 6680
rect 15998 6673 16033 6680
rect 13152 6668 16033 6673
rect 344 6598 360 6654
rect 394 6598 410 6654
rect 480 6641 582 6657
rect 3382 6641 3484 6657
rect 12884 6641 12986 6657
rect 514 6607 548 6641
rect 3416 6607 3450 6641
rect 12918 6607 12952 6641
rect 13152 6634 13194 6668
rect 13228 6634 13264 6668
rect 13298 6634 13334 6668
rect 13368 6634 13404 6668
rect 13438 6634 13474 6668
rect 13508 6634 13544 6668
rect 13578 6634 13614 6668
rect 13648 6634 13684 6668
rect 13718 6634 13754 6668
rect 13788 6634 13824 6668
rect 13858 6634 13894 6668
rect 13928 6634 13964 6668
rect 13998 6634 14034 6668
rect 14068 6634 14104 6668
rect 14138 6634 14174 6668
rect 14208 6634 14244 6668
rect 14278 6634 14314 6668
rect 14348 6634 14384 6668
rect 14418 6634 14454 6668
rect 14488 6634 14524 6668
rect 14558 6634 14594 6668
rect 14628 6634 14664 6668
rect 14698 6642 16033 6668
rect 14698 6638 15733 6642
rect 15767 6638 15819 6642
rect 15853 6638 15905 6642
rect 15939 6638 15991 6642
rect 14698 6634 14774 6638
rect 344 6585 410 6598
rect 480 6591 582 6607
rect 3382 6591 3484 6607
rect 12884 6591 12986 6607
rect 13152 6604 14774 6634
rect 14808 6604 14844 6638
rect 14878 6604 14914 6638
rect 14948 6604 14984 6638
rect 15018 6604 15054 6638
rect 15088 6604 15124 6638
rect 15158 6604 15194 6638
rect 15228 6604 15264 6638
rect 15298 6604 15334 6638
rect 15368 6604 15404 6638
rect 15438 6604 15474 6638
rect 15508 6604 15544 6638
rect 15578 6604 15614 6638
rect 15648 6604 15684 6638
rect 15718 6608 15733 6638
rect 15788 6608 15819 6638
rect 15718 6604 15754 6608
rect 15788 6604 15824 6608
rect 15858 6604 15894 6638
rect 15939 6608 15964 6638
rect 16025 6608 16033 6642
rect 15928 6604 15964 6608
rect 15998 6604 16033 6608
rect 13152 6598 16033 6604
rect 344 6526 360 6585
rect 394 6526 410 6585
rect 344 6516 410 6526
rect 344 6454 360 6516
rect 394 6454 410 6516
rect 13152 6564 13194 6598
rect 13228 6564 13264 6598
rect 13298 6564 13334 6598
rect 13368 6564 13404 6598
rect 13438 6564 13474 6598
rect 13508 6564 13544 6598
rect 13578 6564 13614 6598
rect 13648 6564 13684 6598
rect 13718 6564 13754 6598
rect 13788 6564 13824 6598
rect 13858 6564 13894 6598
rect 13928 6564 13964 6598
rect 13998 6564 14034 6598
rect 14068 6564 14104 6598
rect 14138 6564 14174 6598
rect 14208 6564 14244 6598
rect 14278 6564 14314 6598
rect 14348 6564 14384 6598
rect 14418 6564 14454 6598
rect 14488 6564 14524 6598
rect 14558 6564 14594 6598
rect 14628 6564 14664 6598
rect 14698 6570 16033 6598
rect 14698 6569 15733 6570
rect 15767 6569 15819 6570
rect 15853 6569 15905 6570
rect 15939 6569 15991 6570
rect 14698 6564 14774 6569
rect 13152 6535 14774 6564
rect 14808 6535 14844 6569
rect 14878 6535 14914 6569
rect 14948 6535 14984 6569
rect 15018 6535 15054 6569
rect 15088 6535 15124 6569
rect 15158 6535 15194 6569
rect 15228 6535 15264 6569
rect 15298 6535 15334 6569
rect 15368 6535 15404 6569
rect 15438 6535 15474 6569
rect 15508 6535 15544 6569
rect 15578 6535 15614 6569
rect 15648 6535 15684 6569
rect 15718 6536 15733 6569
rect 15788 6536 15819 6569
rect 15718 6535 15754 6536
rect 15788 6535 15824 6536
rect 15858 6535 15894 6569
rect 15939 6536 15964 6569
rect 16025 6536 16033 6570
rect 15928 6535 15964 6536
rect 15998 6535 16033 6536
rect 13152 6528 16033 6535
rect 480 6487 582 6503
rect 3382 6487 3484 6503
rect 12884 6487 12986 6503
rect 13152 6494 13194 6528
rect 13228 6494 13264 6528
rect 13298 6494 13334 6528
rect 13368 6494 13404 6528
rect 13438 6494 13474 6528
rect 13508 6494 13544 6528
rect 13578 6494 13614 6528
rect 13648 6494 13684 6528
rect 13718 6494 13754 6528
rect 13788 6494 13824 6528
rect 13858 6494 13894 6528
rect 13928 6494 13964 6528
rect 13998 6494 14034 6528
rect 14068 6494 14104 6528
rect 14138 6494 14174 6528
rect 14208 6494 14244 6528
rect 14278 6494 14314 6528
rect 14348 6494 14384 6528
rect 14418 6494 14454 6528
rect 14488 6494 14524 6528
rect 14558 6494 14594 6528
rect 14628 6494 14664 6528
rect 14698 6500 16033 6528
rect 14698 6494 14774 6500
rect 344 6447 410 6454
rect 514 6453 548 6487
rect 3416 6453 3450 6487
rect 12918 6453 12952 6487
rect 13152 6466 14774 6494
rect 14808 6466 14844 6500
rect 14878 6466 14914 6500
rect 14948 6466 14984 6500
rect 15018 6466 15054 6500
rect 15088 6466 15124 6500
rect 15158 6466 15194 6500
rect 15228 6466 15264 6500
rect 15298 6466 15334 6500
rect 15368 6466 15404 6500
rect 15438 6466 15474 6500
rect 15508 6466 15544 6500
rect 15578 6466 15614 6500
rect 15648 6466 15684 6500
rect 15718 6498 15754 6500
rect 15788 6498 15824 6500
rect 15718 6466 15733 6498
rect 15788 6466 15819 6498
rect 15858 6466 15894 6500
rect 15928 6498 15964 6500
rect 15998 6498 16033 6500
rect 15939 6466 15964 6498
rect 13152 6464 15733 6466
rect 15767 6464 15819 6466
rect 15853 6464 15905 6466
rect 15939 6464 15991 6466
rect 16025 6464 16033 6498
rect 13152 6458 16033 6464
rect 344 6382 360 6447
rect 394 6382 410 6447
rect 480 6437 582 6453
rect 3382 6437 3484 6453
rect 12884 6437 12986 6453
rect 344 6378 410 6382
rect 344 6310 360 6378
rect 394 6310 410 6378
rect 13152 6424 13194 6458
rect 13228 6424 13264 6458
rect 13298 6424 13334 6458
rect 13368 6424 13404 6458
rect 13438 6424 13474 6458
rect 13508 6424 13544 6458
rect 13578 6424 13614 6458
rect 13648 6424 13684 6458
rect 13718 6424 13754 6458
rect 13788 6424 13824 6458
rect 13858 6424 13894 6458
rect 13928 6424 13964 6458
rect 13998 6424 14034 6458
rect 14068 6424 14104 6458
rect 14138 6424 14174 6458
rect 14208 6424 14244 6458
rect 14278 6424 14314 6458
rect 14348 6424 14384 6458
rect 14418 6424 14454 6458
rect 14488 6424 14524 6458
rect 14558 6424 14594 6458
rect 14628 6424 14664 6458
rect 14698 6431 16033 6458
rect 14698 6424 14774 6431
rect 13152 6397 14774 6424
rect 14808 6397 14844 6431
rect 14878 6397 14914 6431
rect 14948 6397 14984 6431
rect 15018 6397 15054 6431
rect 15088 6397 15124 6431
rect 15158 6397 15194 6431
rect 15228 6397 15264 6431
rect 15298 6397 15334 6431
rect 15368 6397 15404 6431
rect 15438 6397 15474 6431
rect 15508 6397 15544 6431
rect 15578 6397 15614 6431
rect 15648 6397 15684 6431
rect 15718 6426 15754 6431
rect 15788 6426 15824 6431
rect 15718 6397 15733 6426
rect 15788 6397 15819 6426
rect 15858 6397 15894 6431
rect 15928 6426 15964 6431
rect 15998 6426 16033 6431
rect 15939 6397 15964 6426
rect 13152 6392 15733 6397
rect 15767 6392 15819 6397
rect 15853 6392 15905 6397
rect 15939 6392 15991 6397
rect 16025 6392 16033 6426
rect 13152 6388 16033 6392
rect 13152 6354 13194 6388
rect 13228 6354 13264 6388
rect 13298 6354 13334 6388
rect 13368 6354 13404 6388
rect 13438 6354 13474 6388
rect 13508 6354 13544 6388
rect 13578 6354 13614 6388
rect 13648 6354 13684 6388
rect 13718 6354 13754 6388
rect 13788 6354 13824 6388
rect 13858 6354 13894 6388
rect 13928 6354 13964 6388
rect 13998 6354 14034 6388
rect 14068 6354 14104 6388
rect 14138 6354 14174 6388
rect 14208 6354 14244 6388
rect 14278 6354 14314 6388
rect 14348 6354 14384 6388
rect 14418 6354 14454 6388
rect 14488 6354 14524 6388
rect 14558 6354 14594 6388
rect 14628 6354 14664 6388
rect 14698 6362 16033 6388
rect 14698 6354 14774 6362
rect 480 6333 582 6349
rect 3382 6333 3484 6349
rect 12884 6333 12986 6349
rect 344 6309 410 6310
rect 344 6275 360 6309
rect 394 6275 410 6309
rect 514 6299 548 6333
rect 3416 6299 3450 6333
rect 12918 6299 12952 6333
rect 13152 6328 14774 6354
rect 14808 6328 14844 6362
rect 14878 6328 14914 6362
rect 14948 6328 14984 6362
rect 15018 6328 15054 6362
rect 15088 6328 15124 6362
rect 15158 6328 15194 6362
rect 15228 6328 15264 6362
rect 15298 6328 15334 6362
rect 15368 6328 15404 6362
rect 15438 6328 15474 6362
rect 15508 6328 15544 6362
rect 15578 6328 15614 6362
rect 15648 6328 15684 6362
rect 15718 6354 15754 6362
rect 15788 6354 15824 6362
rect 15718 6328 15733 6354
rect 15788 6328 15819 6354
rect 15858 6328 15894 6362
rect 15928 6354 15964 6362
rect 15998 6354 16033 6362
rect 15939 6328 15964 6354
rect 13152 6320 15733 6328
rect 15767 6320 15819 6328
rect 15853 6320 15905 6328
rect 15939 6320 15991 6328
rect 16025 6320 16033 6354
rect 13152 6318 16033 6320
rect 480 6283 582 6299
rect 3382 6283 3484 6299
rect 12884 6283 12986 6299
rect 13152 6284 13194 6318
rect 13228 6284 13264 6318
rect 13298 6284 13334 6318
rect 13368 6284 13404 6318
rect 13438 6284 13474 6318
rect 13508 6284 13544 6318
rect 13578 6284 13614 6318
rect 13648 6284 13684 6318
rect 13718 6284 13754 6318
rect 13788 6284 13824 6318
rect 13858 6284 13894 6318
rect 13928 6284 13964 6318
rect 13998 6284 14034 6318
rect 14068 6284 14104 6318
rect 14138 6284 14174 6318
rect 14208 6284 14244 6318
rect 14278 6284 14314 6318
rect 14348 6284 14384 6318
rect 14418 6284 14454 6318
rect 14488 6284 14524 6318
rect 14558 6284 14594 6318
rect 14628 6284 14664 6318
rect 14698 6293 16033 6318
rect 14698 6284 14774 6293
rect 344 6272 410 6275
rect 344 6206 360 6272
rect 394 6206 410 6272
rect 344 6200 410 6206
rect 344 6137 360 6200
rect 394 6137 410 6200
rect 13152 6259 14774 6284
rect 14808 6259 14844 6293
rect 14878 6259 14914 6293
rect 14948 6259 14984 6293
rect 15018 6259 15054 6293
rect 15088 6259 15124 6293
rect 15158 6259 15194 6293
rect 15228 6259 15264 6293
rect 15298 6259 15334 6293
rect 15368 6259 15404 6293
rect 15438 6259 15474 6293
rect 15508 6259 15544 6293
rect 15578 6259 15614 6293
rect 15648 6259 15684 6293
rect 15718 6282 15754 6293
rect 15788 6282 15824 6293
rect 15718 6259 15733 6282
rect 15788 6259 15819 6282
rect 15858 6259 15894 6293
rect 15928 6282 15964 6293
rect 15998 6282 16033 6293
rect 15939 6259 15964 6282
rect 13152 6248 15733 6259
rect 15767 6248 15819 6259
rect 15853 6248 15905 6259
rect 15939 6248 15991 6259
rect 16025 6248 16033 6282
rect 13152 6214 13194 6248
rect 13228 6214 13264 6248
rect 13298 6214 13334 6248
rect 13368 6214 13404 6248
rect 13438 6214 13474 6248
rect 13508 6214 13544 6248
rect 13578 6214 13614 6248
rect 13648 6214 13684 6248
rect 13718 6214 13754 6248
rect 13788 6214 13824 6248
rect 13858 6214 13894 6248
rect 13928 6214 13964 6248
rect 13998 6214 14034 6248
rect 14068 6214 14104 6248
rect 14138 6214 14174 6248
rect 14208 6214 14244 6248
rect 14278 6214 14314 6248
rect 14348 6214 14384 6248
rect 14418 6214 14454 6248
rect 14488 6214 14524 6248
rect 14558 6214 14594 6248
rect 14628 6214 14664 6248
rect 14698 6224 16033 6248
rect 14698 6214 14774 6224
rect 480 6179 582 6195
rect 3382 6179 3484 6195
rect 12884 6179 12986 6195
rect 13152 6190 14774 6214
rect 14808 6190 14844 6224
rect 14878 6190 14914 6224
rect 14948 6190 14984 6224
rect 15018 6190 15054 6224
rect 15088 6190 15124 6224
rect 15158 6190 15194 6224
rect 15228 6190 15264 6224
rect 15298 6190 15334 6224
rect 15368 6190 15404 6224
rect 15438 6190 15474 6224
rect 15508 6190 15544 6224
rect 15578 6190 15614 6224
rect 15648 6190 15684 6224
rect 15718 6210 15754 6224
rect 15788 6210 15824 6224
rect 15718 6190 15733 6210
rect 15788 6190 15819 6210
rect 15858 6190 15894 6224
rect 15928 6210 15964 6224
rect 15998 6210 16033 6224
rect 15939 6190 15964 6210
rect 514 6145 548 6179
rect 3416 6145 3450 6179
rect 12918 6145 12952 6179
rect 13152 6178 15733 6190
rect 344 6128 410 6137
rect 480 6129 582 6145
rect 3382 6129 3484 6145
rect 12884 6129 12986 6145
rect 13152 6144 13194 6178
rect 13228 6144 13264 6178
rect 13298 6144 13334 6178
rect 13368 6144 13404 6178
rect 13438 6144 13474 6178
rect 13508 6144 13544 6178
rect 13578 6144 13614 6178
rect 13648 6144 13684 6178
rect 13718 6144 13754 6178
rect 13788 6144 13824 6178
rect 13858 6144 13894 6178
rect 13928 6144 13964 6178
rect 13998 6144 14034 6178
rect 14068 6144 14104 6178
rect 14138 6144 14174 6178
rect 14208 6144 14244 6178
rect 14278 6144 14314 6178
rect 14348 6144 14384 6178
rect 14418 6144 14454 6178
rect 14488 6144 14524 6178
rect 14558 6144 14594 6178
rect 14628 6144 14664 6178
rect 14698 6176 15733 6178
rect 15767 6176 15819 6190
rect 15853 6176 15905 6190
rect 15939 6176 15991 6190
rect 16025 6176 16033 6210
rect 14698 6155 16033 6176
rect 14698 6144 14774 6155
rect 344 6068 360 6128
rect 394 6068 410 6128
rect 344 6049 410 6068
rect 13152 6121 14774 6144
rect 14808 6121 14844 6155
rect 14878 6121 14914 6155
rect 14948 6121 14984 6155
rect 15018 6121 15054 6155
rect 15088 6121 15124 6155
rect 15158 6121 15194 6155
rect 15228 6121 15264 6155
rect 15298 6121 15334 6155
rect 15368 6121 15404 6155
rect 15438 6121 15474 6155
rect 15508 6121 15544 6155
rect 15578 6121 15614 6155
rect 15648 6121 15684 6155
rect 15718 6138 15754 6155
rect 15788 6138 15824 6155
rect 15718 6121 15733 6138
rect 15788 6121 15819 6138
rect 15858 6121 15894 6155
rect 15928 6138 15964 6155
rect 15998 6138 16033 6155
rect 15939 6121 15964 6138
rect 13152 6108 15733 6121
rect 13152 6074 13194 6108
rect 13228 6074 13264 6108
rect 13298 6074 13334 6108
rect 13368 6074 13404 6108
rect 13438 6074 13474 6108
rect 13508 6074 13544 6108
rect 13578 6074 13614 6108
rect 13648 6074 13684 6108
rect 13718 6074 13754 6108
rect 13788 6074 13824 6108
rect 13858 6074 13894 6108
rect 13928 6074 13964 6108
rect 13998 6074 14034 6108
rect 14068 6074 14104 6108
rect 14138 6074 14174 6108
rect 14208 6074 14244 6108
rect 14278 6074 14314 6108
rect 14348 6074 14384 6108
rect 14418 6074 14454 6108
rect 14488 6074 14524 6108
rect 14558 6074 14594 6108
rect 14628 6074 14664 6108
rect 14698 6104 15733 6108
rect 15767 6104 15819 6121
rect 15853 6104 15905 6121
rect 15939 6104 15991 6121
rect 16025 6104 16033 6138
rect 14698 6086 16033 6104
rect 14698 6074 14774 6086
rect 13152 6052 14774 6074
rect 14808 6052 14844 6086
rect 14878 6052 14914 6086
rect 14948 6052 14984 6086
rect 15018 6052 15054 6086
rect 15088 6052 15124 6086
rect 15158 6052 15194 6086
rect 15228 6052 15264 6086
rect 15298 6052 15334 6086
rect 15368 6052 15404 6086
rect 15438 6052 15474 6086
rect 15508 6052 15544 6086
rect 15578 6052 15614 6086
rect 15648 6052 15684 6086
rect 15718 6066 15754 6086
rect 15788 6066 15824 6086
rect 15718 6052 15733 6066
rect 15788 6052 15819 6066
rect 15858 6052 15894 6086
rect 15928 6066 15964 6086
rect 15998 6066 16033 6086
rect 15939 6052 15964 6066
rect 13152 6049 15733 6052
rect 344 6033 14647 6049
rect 344 5999 360 6033
rect 423 5999 429 6033
rect 495 5999 498 6033
rect 532 5999 533 6033
rect 601 5999 605 6033
rect 670 5999 677 6033
rect 739 6032 774 6033
rect 808 6032 843 6033
rect 739 5999 765 6032
rect 808 5999 837 6032
rect 877 5999 912 6033
rect 948 5999 981 6033
rect 1020 5999 1050 6033
rect 1092 5999 1119 6033
rect 1164 5999 1188 6033
rect 1236 5999 1257 6033
rect 1308 5999 1326 6033
rect 1380 5999 1395 6033
rect 1452 5999 1464 6033
rect 1524 5999 1533 6033
rect 1596 5999 1602 6033
rect 1668 5999 1671 6033
rect 1705 5999 1706 6033
rect 1774 5999 1778 6033
rect 1843 5999 1850 6033
rect 1912 5999 1922 6033
rect 1981 5999 1994 6033
rect 2050 5999 2066 6033
rect 2119 5999 2138 6033
rect 2188 5999 2210 6033
rect 2257 5999 2282 6033
rect 2326 5999 2354 6033
rect 2395 5999 2426 6033
rect 2464 5999 2498 6033
rect 2533 5999 2568 6033
rect 2604 5999 2637 6033
rect 2676 5999 2706 6033
rect 2748 5999 2775 6033
rect 2820 5999 2844 6033
rect 2892 5999 2913 6033
rect 2964 5999 2982 6033
rect 3036 5999 3051 6033
rect 3108 5999 3120 6033
rect 3180 5999 3189 6033
rect 3252 5999 3257 6033
rect 3324 5999 3325 6033
rect 3359 5999 3362 6033
rect 3427 5999 3434 6033
rect 3495 5999 3506 6033
rect 3563 5999 3578 6033
rect 3631 5999 3650 6033
rect 3699 5999 3722 6033
rect 3767 5999 3794 6033
rect 3835 5999 3866 6033
rect 3903 5999 3937 6033
rect 3972 5999 4005 6033
rect 4044 5999 4073 6033
rect 4116 5999 4141 6033
rect 4188 5999 4209 6033
rect 4260 5999 4277 6033
rect 4332 5999 4345 6033
rect 4404 5999 4413 6033
rect 4476 5999 4481 6033
rect 4548 5999 4549 6033
rect 4583 5999 4617 6033
rect 4651 6032 4685 6033
rect 4719 6032 4753 6033
rect 4652 5999 4685 6032
rect 4724 5999 4753 6032
rect 4807 5999 4821 6033
rect 4879 5999 4889 6033
rect 4951 5999 4957 6033
rect 5023 5999 5025 6033
rect 5059 5999 5061 6033
rect 5127 5999 5133 6033
rect 5195 5999 5205 6033
rect 5263 5999 5277 6033
rect 5331 5999 5349 6033
rect 5399 5999 5421 6033
rect 5467 5999 5493 6033
rect 5535 5999 5565 6033
rect 5603 5999 5637 6033
rect 5671 5999 5705 6033
rect 5743 5999 5773 6033
rect 5815 5999 5841 6033
rect 5887 5999 5909 6033
rect 5943 5999 5977 6033
rect 6011 5999 6045 6033
rect 6079 5999 6113 6033
rect 6147 5999 6181 6033
rect 6229 5999 6249 6033
rect 6303 5999 6317 6033
rect 6376 5999 6385 6033
rect 6449 5999 6453 6033
rect 6487 5999 6488 6033
rect 6555 5999 6561 6033
rect 6623 5999 6634 6033
rect 6691 5999 6707 6033
rect 6759 5999 6780 6033
rect 6827 5999 6861 6033
rect 6895 5999 6929 6033
rect 6963 5999 6997 6033
rect 7031 5999 7065 6033
rect 7103 5999 7133 6033
rect 7175 5999 7201 6033
rect 7247 5999 7269 6033
rect 7319 5999 7337 6033
rect 7391 5999 7405 6033
rect 7463 5999 7473 6033
rect 7535 5999 7541 6033
rect 7607 5999 7609 6033
rect 7643 5999 7677 6033
rect 7711 5999 7745 6033
rect 7779 5999 7813 6033
rect 7847 5999 7881 6033
rect 7915 5999 7932 6033
rect 7983 5999 8004 6033
rect 8051 5999 8076 6033
rect 8119 5999 8148 6033
rect 8187 5999 8220 6033
rect 8255 5999 8289 6033
rect 8326 5999 8357 6033
rect 8398 5999 8425 6033
rect 8470 5999 8493 6033
rect 8527 5999 8561 6033
rect 8595 5999 8629 6033
rect 8663 5999 8697 6033
rect 8731 5999 8765 6033
rect 8824 5999 8833 6033
rect 8896 5999 8901 6033
rect 8968 5999 8969 6033
rect 9003 5999 9006 6033
rect 9071 5999 9078 6033
rect 9139 5999 9150 6033
rect 9207 5999 9222 6033
rect 9275 5999 9294 6033
rect 9343 5999 9377 6033
rect 9411 5999 9445 6033
rect 9479 5999 9513 6033
rect 9547 5999 9581 6033
rect 9615 5999 9628 6033
rect 9683 5999 9700 6033
rect 9751 5999 9772 6033
rect 9819 5999 9844 6033
rect 9887 5999 9916 6033
rect 9955 5999 9988 6033
rect 10023 5999 10057 6033
rect 10094 5999 10125 6033
rect 10166 5999 10193 6033
rect 10227 5999 10261 6033
rect 10295 5999 10329 6033
rect 10363 5999 10397 6033
rect 10431 5999 10465 6033
rect 10499 5999 10533 6033
rect 10572 5999 10601 6033
rect 10644 5999 10669 6033
rect 10716 5999 10737 6033
rect 10788 5999 10805 6033
rect 10860 5999 10873 6033
rect 10932 5999 10941 6033
rect 11004 5999 11009 6033
rect 11076 5999 11077 6033
rect 11111 5999 11114 6033
rect 11179 5999 11186 6033
rect 11247 5999 11258 6033
rect 11315 5999 11330 6033
rect 11383 5999 11402 6033
rect 11451 5999 11474 6033
rect 11519 5999 11546 6033
rect 11587 5999 11618 6033
rect 11655 5999 11689 6033
rect 11724 5999 11757 6033
rect 11796 5999 11825 6033
rect 11868 5999 11893 6033
rect 11940 5999 11961 6033
rect 12012 5999 12029 6033
rect 12084 5999 12097 6033
rect 12156 5999 12165 6033
rect 12228 5999 12233 6033
rect 12300 5999 12301 6033
rect 12335 5999 12338 6033
rect 12403 5999 12410 6033
rect 12471 5999 12482 6033
rect 12539 5999 12554 6033
rect 12607 5999 12626 6033
rect 12675 5999 12698 6033
rect 12743 5999 12770 6033
rect 12811 5999 12842 6033
rect 12879 5999 12913 6033
rect 12948 5999 12981 6033
rect 13020 5999 13049 6033
rect 13092 5999 13117 6033
rect 13151 5999 13165 6033
rect 13219 5999 13240 6033
rect 13287 5999 13315 6033
rect 13355 5999 13389 6033
rect 13424 5999 13457 6033
rect 13499 5999 13525 6033
rect 13574 5999 13593 6033
rect 13649 5999 13661 6033
rect 13724 5999 13729 6033
rect 13763 5999 13765 6033
rect 13831 5999 13840 6033
rect 13899 5999 13915 6033
rect 13967 5999 13990 6033
rect 14035 5999 14065 6033
rect 14103 5999 14137 6033
rect 14174 5999 14205 6033
rect 14249 5999 14273 6033
rect 14324 5999 14341 6033
rect 14399 5999 14409 6033
rect 14474 5999 14477 6033
rect 14511 5999 14515 6033
rect 14579 5999 14613 6033
rect 344 5998 765 5999
rect 799 5998 837 5999
rect 871 5998 4618 5999
rect 4652 5998 4690 5999
rect 4724 5998 14647 5999
rect 344 5983 14647 5998
rect 14740 6032 15733 6049
rect 15767 6032 15819 6052
rect 15853 6032 15905 6052
rect 15939 6032 15991 6052
rect 16025 6032 16033 6066
rect 14740 6017 16033 6032
rect 14740 5983 14774 6017
rect 14808 5983 14844 6017
rect 14878 5983 14914 6017
rect 14948 5983 14984 6017
rect 15018 5983 15054 6017
rect 15088 5983 15124 6017
rect 15158 5983 15194 6017
rect 15228 5983 15264 6017
rect 15298 5983 15334 6017
rect 15368 5983 15404 6017
rect 15438 5983 15474 6017
rect 15508 5983 15544 6017
rect 15578 5983 15614 6017
rect 15648 5983 15684 6017
rect 15718 5994 15754 6017
rect 15788 5994 15824 6017
rect 15718 5983 15733 5994
rect 15788 5983 15819 5994
rect 15858 5983 15894 6017
rect 15928 5994 15964 6017
rect 15998 5994 16033 6017
rect 15939 5983 15964 5994
rect 11482 5951 11564 5975
rect 11482 5917 11506 5951
rect 11540 5917 11564 5951
rect 11482 5882 11564 5917
rect 14740 5960 15733 5983
rect 15767 5960 15819 5983
rect 15853 5960 15905 5983
rect 15939 5960 15991 5983
rect 16025 5960 16033 5994
rect 14740 5948 16033 5960
rect 14740 5914 14774 5948
rect 14808 5914 14844 5948
rect 14878 5914 14914 5948
rect 14948 5914 14984 5948
rect 15018 5914 15054 5948
rect 15088 5914 15124 5948
rect 15158 5914 15194 5948
rect 15228 5914 15264 5948
rect 15298 5914 15334 5948
rect 15368 5914 15404 5948
rect 15438 5914 15474 5948
rect 15508 5914 15544 5948
rect 15578 5914 15614 5948
rect 15648 5914 15684 5948
rect 15718 5922 15754 5948
rect 15788 5922 15824 5948
rect 15718 5914 15733 5922
rect 15788 5914 15819 5922
rect 15858 5914 15894 5948
rect 15928 5922 15964 5948
rect 15998 5922 16033 5948
rect 15939 5914 15964 5922
rect 11482 5848 11506 5882
rect 11540 5848 11564 5882
rect 11626 5888 11728 5904
rect 14528 5888 14630 5904
rect 14740 5888 15733 5914
rect 15767 5888 15819 5914
rect 15853 5888 15905 5914
rect 15939 5888 15991 5914
rect 16025 5888 16033 5922
rect 344 5799 10922 5815
rect 344 5731 360 5799
rect 394 5765 428 5799
rect 468 5765 496 5799
rect 540 5765 564 5799
rect 612 5765 632 5799
rect 684 5765 700 5799
rect 756 5765 768 5799
rect 828 5765 836 5799
rect 900 5765 904 5799
rect 1006 5765 1010 5799
rect 1074 5765 1082 5799
rect 1142 5765 1154 5799
rect 1210 5765 1226 5799
rect 1278 5765 1298 5799
rect 1346 5765 1370 5799
rect 1414 5765 1442 5799
rect 1482 5765 1514 5799
rect 1550 5765 1584 5799
rect 1620 5765 1652 5799
rect 1692 5765 1720 5799
rect 1764 5765 1788 5799
rect 1836 5765 1856 5799
rect 1908 5765 1924 5799
rect 1980 5765 1992 5799
rect 2052 5765 2060 5799
rect 2124 5765 2128 5799
rect 2230 5765 2234 5799
rect 2298 5765 2306 5799
rect 2366 5765 2378 5799
rect 2434 5765 2450 5799
rect 2502 5765 2522 5799
rect 2570 5765 2594 5799
rect 2638 5765 2666 5799
rect 2706 5765 2738 5799
rect 2774 5765 2808 5799
rect 2844 5765 2876 5799
rect 2916 5765 2944 5799
rect 2988 5765 3012 5799
rect 3060 5765 3080 5799
rect 3132 5765 3148 5799
rect 3204 5765 3216 5799
rect 3276 5765 3284 5799
rect 3348 5765 3352 5799
rect 3454 5765 3458 5799
rect 3522 5765 3530 5799
rect 3590 5765 3602 5799
rect 3658 5765 3674 5799
rect 3726 5765 3746 5799
rect 3794 5765 3818 5799
rect 3862 5765 3890 5799
rect 3930 5765 3962 5799
rect 3998 5765 4032 5799
rect 4068 5765 4100 5799
rect 4140 5765 4168 5799
rect 4212 5765 4236 5799
rect 4284 5765 4304 5799
rect 4356 5765 4372 5799
rect 4428 5765 4440 5799
rect 4500 5765 4508 5799
rect 4572 5765 4576 5799
rect 4678 5765 4682 5799
rect 4746 5765 4754 5799
rect 4814 5765 4826 5799
rect 4882 5765 4898 5799
rect 4950 5765 4970 5799
rect 5018 5765 5042 5799
rect 5086 5765 5114 5799
rect 5154 5765 5186 5799
rect 5222 5765 5256 5799
rect 5292 5765 5324 5799
rect 5364 5765 5392 5799
rect 5436 5765 5460 5799
rect 5508 5765 5528 5799
rect 5580 5765 5596 5799
rect 5652 5765 5664 5799
rect 5724 5765 5732 5799
rect 5797 5765 5800 5799
rect 5834 5765 5836 5799
rect 5902 5765 5909 5799
rect 5970 5765 6004 5799
rect 6038 5765 6072 5799
rect 6106 5765 6140 5799
rect 6174 5765 6195 5799
rect 6242 5765 6269 5799
rect 6310 5765 6342 5799
rect 6378 5765 6412 5799
rect 6449 5765 6480 5799
rect 6522 5765 6548 5799
rect 6595 5765 6616 5799
rect 6668 5765 6684 5799
rect 6741 5765 6752 5799
rect 6814 5765 6820 5799
rect 6854 5765 6888 5799
rect 6922 5765 6956 5799
rect 6990 5765 7024 5799
rect 7058 5765 7069 5799
rect 7126 5765 7141 5799
rect 7194 5765 7213 5799
rect 7262 5765 7285 5799
rect 7330 5765 7357 5799
rect 7398 5765 7429 5799
rect 7466 5765 7500 5799
rect 7535 5765 7568 5799
rect 7607 5765 7636 5799
rect 7670 5765 7704 5799
rect 7738 5765 7772 5799
rect 7806 5765 7840 5799
rect 7874 5765 7908 5799
rect 7966 5765 7976 5799
rect 8038 5765 8044 5799
rect 8110 5765 8112 5799
rect 8146 5765 8148 5799
rect 8215 5765 8220 5799
rect 8284 5765 8292 5799
rect 8353 5765 8364 5799
rect 8422 5765 8436 5799
rect 8491 5765 8526 5799
rect 8560 5765 8595 5799
rect 8629 5765 8664 5799
rect 8698 5765 8733 5799
rect 8767 5765 8790 5799
rect 8836 5765 8862 5799
rect 8905 5765 8934 5799
rect 8974 5765 9006 5799
rect 9043 5765 9078 5799
rect 9112 5765 9147 5799
rect 9184 5765 9216 5799
rect 9256 5765 9285 5799
rect 9328 5765 9354 5799
rect 9388 5765 9423 5799
rect 9457 5765 9492 5799
rect 9526 5765 9561 5799
rect 9595 5765 9628 5799
rect 9664 5765 9699 5799
rect 9734 5765 9768 5799
rect 9806 5765 9837 5799
rect 9878 5765 9906 5799
rect 9950 5765 9975 5799
rect 10022 5765 10044 5799
rect 10094 5765 10113 5799
rect 10166 5765 10182 5799
rect 10216 5765 10251 5799
rect 10285 5765 10320 5799
rect 10354 5765 10389 5799
rect 10423 5765 10458 5799
rect 10521 5765 10527 5799
rect 10593 5765 10596 5799
rect 10630 5765 10631 5799
rect 10699 5765 10703 5799
rect 10768 5765 10775 5799
rect 10837 5765 10847 5799
rect 10906 5765 10922 5799
rect 394 5749 10922 5765
rect 394 5731 410 5749
rect 344 5724 410 5731
rect 344 5659 360 5724
rect 394 5659 410 5724
rect 344 5649 410 5659
rect 344 5587 360 5649
rect 394 5587 410 5649
rect 10856 5730 10922 5749
rect 10856 5676 10872 5730
rect 10906 5676 10922 5730
rect 10856 5661 10922 5676
rect 344 5575 410 5587
rect 344 5515 360 5575
rect 394 5515 410 5575
rect 344 5501 410 5515
rect 344 5443 360 5501
rect 394 5443 410 5501
rect 344 5427 410 5443
rect 344 5371 360 5427
rect 394 5371 410 5427
rect 344 5333 410 5371
rect 344 5287 360 5333
rect 394 5287 410 5333
rect 344 5261 410 5287
rect 344 5217 360 5261
rect 394 5217 410 5261
rect 344 5189 410 5217
rect 344 5147 360 5189
rect 394 5147 410 5189
rect 344 5117 410 5147
rect 344 5077 360 5117
rect 394 5077 410 5117
rect 344 5045 410 5077
rect 344 5007 360 5045
rect 394 5007 410 5045
rect 344 4973 410 5007
rect 344 4937 360 4973
rect 394 4937 410 4973
rect 344 4902 410 4937
rect 344 4867 360 4902
rect 394 4867 410 4902
rect 344 4833 410 4867
rect 344 4795 360 4833
rect 394 4795 410 4833
rect 344 4764 410 4795
rect 344 4723 360 4764
rect 394 4723 410 4764
rect 344 4695 410 4723
rect 344 4651 360 4695
rect 394 4651 410 4695
rect 344 4626 410 4651
rect 344 4579 360 4626
rect 394 4579 410 4626
rect 344 4557 410 4579
rect 344 4507 360 4557
rect 394 4507 410 4557
rect 344 4488 410 4507
rect 344 4435 360 4488
rect 394 4435 410 4488
rect 344 4419 410 4435
rect 344 4363 360 4419
rect 394 4363 410 4419
rect 344 4350 410 4363
rect 344 4291 360 4350
rect 394 4291 410 4350
rect 344 4281 410 4291
rect 480 5625 514 5641
rect 480 5557 514 5591
rect 480 5489 514 5523
rect 480 5421 514 5455
rect 480 5353 514 5377
rect 480 5285 514 5305
rect 480 5217 514 5233
rect 480 5149 514 5161
rect 480 5081 514 5089
rect 480 5013 514 5017
rect 480 4907 514 4911
rect 480 4835 514 4843
rect 480 4763 514 4775
rect 480 4691 514 4707
rect 480 4619 514 4639
rect 480 4547 514 4571
rect 480 4469 514 4503
rect 480 4401 514 4435
rect 480 4333 514 4367
rect 480 4283 514 4299
rect 1336 5625 1370 5641
rect 1336 5557 1370 5591
rect 1336 5489 1370 5523
rect 1336 5421 1370 5455
rect 1336 5353 1370 5377
rect 1336 5285 1370 5305
rect 1336 5217 1370 5233
rect 1336 5149 1370 5161
rect 1336 5081 1370 5089
rect 1336 5013 1370 5017
rect 1336 4907 1370 4911
rect 1336 4835 1370 4843
rect 1336 4763 1370 4775
rect 1336 4691 1370 4707
rect 1336 4619 1370 4639
rect 1336 4547 1370 4571
rect 1336 4469 1370 4503
rect 1336 4401 1370 4435
rect 1336 4333 1370 4367
rect 1336 4283 1370 4299
rect 2192 5625 2226 5641
rect 2192 5557 2226 5591
rect 2192 5489 2226 5523
rect 2192 5421 2226 5455
rect 2192 5353 2226 5377
rect 2192 5285 2226 5305
rect 2192 5217 2226 5233
rect 2192 5149 2226 5161
rect 2192 5081 2226 5089
rect 2192 5013 2226 5017
rect 2192 4907 2226 4911
rect 2192 4835 2226 4843
rect 2192 4763 2226 4775
rect 2192 4691 2226 4707
rect 2192 4619 2226 4639
rect 2192 4547 2226 4571
rect 2192 4469 2226 4503
rect 2192 4401 2226 4435
rect 2192 4333 2226 4367
rect 2192 4283 2226 4299
rect 3048 5625 3082 5641
rect 3048 5557 3082 5591
rect 3048 5489 3082 5523
rect 3048 5421 3082 5455
rect 3048 5353 3082 5377
rect 3048 5285 3082 5305
rect 3048 5217 3082 5233
rect 3048 5149 3082 5161
rect 3048 5081 3082 5089
rect 3048 5013 3082 5017
rect 3048 4907 3082 4911
rect 3048 4835 3082 4843
rect 3048 4763 3082 4775
rect 3048 4691 3082 4707
rect 3048 4619 3082 4639
rect 3048 4547 3082 4571
rect 3048 4469 3082 4503
rect 3048 4401 3082 4435
rect 3048 4333 3082 4367
rect 3048 4283 3082 4299
rect 3904 5625 3938 5641
rect 3904 5557 3938 5591
rect 3904 5489 3938 5523
rect 3904 5421 3938 5455
rect 3904 5353 3938 5377
rect 3904 5285 3938 5305
rect 3904 5217 3938 5233
rect 3904 5149 3938 5161
rect 3904 5081 3938 5089
rect 3904 5013 3938 5017
rect 3904 4907 3938 4911
rect 3904 4835 3938 4843
rect 3904 4763 3938 4775
rect 3904 4691 3938 4707
rect 3904 4619 3938 4639
rect 3904 4547 3938 4571
rect 3904 4469 3938 4503
rect 3904 4401 3938 4435
rect 3904 4333 3938 4367
rect 3904 4283 3938 4299
rect 4760 5625 4794 5641
rect 4760 5557 4794 5591
rect 4760 5489 4794 5523
rect 4760 5421 4794 5455
rect 4760 5353 4794 5377
rect 4760 5285 4794 5305
rect 4760 5217 4794 5233
rect 4760 5149 4794 5161
rect 4760 5081 4794 5089
rect 4760 5013 4794 5017
rect 4760 4907 4794 4911
rect 4760 4835 4794 4843
rect 4760 4763 4794 4775
rect 4760 4691 4794 4707
rect 4760 4619 4794 4639
rect 4760 4547 4794 4571
rect 4760 4469 4794 4503
rect 4760 4401 4794 4435
rect 4760 4333 4794 4367
rect 4760 4283 4794 4299
rect 5616 5625 5650 5641
rect 5616 5557 5650 5591
rect 5616 5489 5650 5523
rect 5616 5421 5650 5455
rect 5616 5353 5650 5377
rect 5616 5285 5650 5305
rect 5616 5217 5650 5233
rect 5616 5149 5650 5161
rect 5616 5081 5650 5089
rect 5616 5013 5650 5017
rect 5616 4907 5650 4911
rect 5616 4835 5650 4843
rect 5616 4763 5650 4775
rect 5616 4691 5650 4707
rect 5616 4619 5650 4639
rect 5616 4547 5650 4571
rect 5616 4469 5650 4503
rect 5616 4401 5650 4435
rect 5616 4333 5650 4367
rect 5616 4283 5650 4299
rect 6472 5625 6506 5641
rect 6472 5557 6506 5591
rect 6472 5489 6506 5523
rect 6472 5421 6506 5455
rect 6472 5353 6506 5377
rect 6472 5285 6506 5305
rect 6472 5217 6506 5233
rect 6472 5149 6506 5161
rect 6472 5081 6506 5089
rect 6472 5013 6506 5017
rect 6472 4907 6506 4911
rect 6472 4835 6506 4843
rect 6472 4763 6506 4775
rect 6472 4691 6506 4707
rect 6472 4619 6506 4639
rect 6472 4547 6506 4571
rect 6472 4469 6506 4503
rect 6472 4401 6506 4435
rect 6472 4333 6506 4367
rect 6472 4283 6506 4299
rect 7328 5625 7362 5641
rect 7328 5557 7362 5591
rect 7328 5489 7362 5523
rect 7328 5421 7362 5455
rect 7328 5353 7362 5377
rect 7328 5285 7362 5305
rect 7328 5217 7362 5233
rect 7328 5149 7362 5161
rect 7328 5081 7362 5089
rect 7328 5013 7362 5017
rect 7328 4907 7362 4911
rect 7328 4835 7362 4843
rect 7328 4763 7362 4775
rect 7328 4691 7362 4707
rect 7328 4619 7362 4639
rect 7328 4547 7362 4571
rect 7328 4469 7362 4503
rect 7328 4401 7362 4435
rect 7328 4333 7362 4367
rect 7328 4283 7362 4299
rect 8184 5625 8218 5641
rect 8184 5557 8218 5591
rect 8184 5489 8218 5523
rect 8184 5421 8218 5455
rect 8184 5353 8218 5377
rect 8184 5285 8218 5305
rect 8184 5217 8218 5233
rect 8184 5149 8218 5161
rect 8184 5081 8218 5089
rect 8184 5013 8218 5017
rect 8184 4907 8218 4911
rect 8184 4835 8218 4843
rect 8184 4763 8218 4775
rect 8184 4691 8218 4707
rect 8184 4619 8218 4639
rect 8184 4547 8218 4571
rect 8184 4469 8218 4503
rect 8184 4401 8218 4435
rect 8184 4333 8218 4367
rect 8184 4283 8218 4299
rect 9040 5625 9074 5641
rect 9040 5557 9074 5591
rect 9040 5489 9074 5523
rect 9040 5421 9074 5455
rect 9040 5353 9074 5377
rect 9040 5285 9074 5305
rect 9040 5217 9074 5233
rect 9040 5149 9074 5161
rect 9040 5081 9074 5089
rect 9040 5013 9074 5017
rect 9040 4907 9074 4911
rect 9040 4835 9074 4843
rect 9040 4763 9074 4775
rect 9040 4691 9074 4707
rect 9040 4619 9074 4639
rect 9040 4547 9074 4571
rect 9040 4469 9074 4503
rect 9040 4401 9074 4435
rect 9040 4333 9074 4367
rect 9040 4283 9074 4299
rect 9896 5625 9930 5641
rect 9896 5557 9930 5591
rect 9896 5489 9930 5523
rect 9896 5421 9930 5455
rect 9896 5353 9930 5377
rect 9896 5285 9930 5305
rect 9896 5217 9930 5233
rect 9896 5149 9930 5161
rect 9896 5081 9930 5089
rect 9896 5013 9930 5017
rect 9896 4907 9930 4911
rect 9896 4835 9930 4843
rect 9896 4763 9930 4775
rect 9896 4691 9930 4707
rect 9896 4619 9930 4639
rect 9896 4547 9930 4571
rect 9896 4469 9930 4503
rect 9896 4401 9930 4435
rect 9896 4333 9930 4367
rect 9896 4283 9930 4299
rect 10752 5625 10786 5641
rect 10752 5557 10786 5591
rect 10752 5489 10786 5523
rect 10752 5421 10786 5455
rect 10752 5353 10786 5377
rect 10752 5285 10786 5305
rect 10752 5217 10786 5233
rect 10752 5149 10786 5161
rect 10752 5081 10786 5089
rect 10752 5013 10786 5017
rect 10752 4907 10786 4911
rect 10752 4835 10786 4843
rect 10752 4763 10786 4775
rect 10752 4691 10786 4707
rect 10752 4619 10786 4639
rect 10752 4547 10786 4571
rect 10752 4469 10786 4503
rect 10752 4401 10786 4435
rect 10752 4333 10786 4367
rect 10752 4283 10786 4299
rect 10856 5604 10872 5661
rect 10906 5604 10922 5661
rect 10856 5592 10922 5604
rect 10856 5532 10872 5592
rect 10906 5532 10922 5592
rect 10856 5523 10922 5532
rect 10856 5460 10872 5523
rect 10906 5460 10922 5523
rect 10856 5454 10922 5460
rect 10856 5388 10872 5454
rect 10906 5388 10922 5454
rect 10856 5385 10922 5388
rect 10856 5351 10872 5385
rect 10906 5351 10922 5385
rect 10856 5350 10922 5351
rect 10856 5282 10872 5350
rect 10906 5282 10922 5350
rect 10856 5278 10922 5282
rect 10856 5213 10872 5278
rect 10906 5213 10922 5278
rect 10856 5206 10922 5213
rect 10856 5144 10872 5206
rect 10906 5144 10922 5206
rect 10856 5134 10922 5144
rect 10856 5075 10872 5134
rect 10906 5075 10922 5134
rect 10856 5062 10922 5075
rect 10856 5006 10872 5062
rect 10906 5006 10922 5062
rect 10856 4990 10922 5006
rect 10856 4937 10872 4990
rect 10906 4937 10922 4990
rect 10856 4918 10922 4937
rect 10856 4868 10872 4918
rect 10906 4868 10922 4918
rect 10856 4846 10922 4868
rect 10856 4799 10872 4846
rect 10906 4799 10922 4846
rect 10856 4774 10922 4799
rect 10856 4730 10872 4774
rect 10906 4730 10922 4774
rect 10856 4702 10922 4730
rect 10856 4661 10872 4702
rect 10906 4661 10922 4702
rect 10856 4630 10922 4661
rect 10856 4592 10872 4630
rect 10906 4592 10922 4630
rect 10856 4558 10922 4592
rect 10856 4523 10872 4558
rect 10906 4523 10922 4558
rect 10856 4488 10922 4523
rect 10856 4452 10872 4488
rect 10906 4452 10922 4488
rect 10856 4419 10922 4452
rect 10856 4380 10872 4419
rect 10906 4380 10922 4419
rect 10856 4350 10922 4380
rect 10856 4308 10872 4350
rect 10906 4308 10922 4350
rect 344 4219 360 4281
rect 394 4219 410 4281
rect 10856 4281 10922 4308
rect 344 4212 410 4219
rect 344 4178 360 4212
rect 394 4178 410 4212
rect 602 4205 632 4239
rect 670 4205 704 4239
rect 745 4205 772 4239
rect 824 4205 840 4239
rect 903 4205 908 4239
rect 942 4205 948 4239
rect 1010 4205 1027 4239
rect 1078 4205 1106 4239
rect 1146 4205 1180 4239
rect 1219 4205 1248 4239
rect 1458 4205 1488 4239
rect 1526 4205 1560 4239
rect 1601 4205 1628 4239
rect 1680 4205 1696 4239
rect 1759 4205 1764 4239
rect 1798 4205 1804 4239
rect 1866 4205 1883 4239
rect 1934 4205 1962 4239
rect 2002 4205 2036 4239
rect 2075 4205 2104 4239
rect 2314 4205 2344 4239
rect 2382 4205 2416 4239
rect 2457 4205 2484 4239
rect 2536 4205 2552 4239
rect 2615 4205 2620 4239
rect 2654 4205 2660 4239
rect 2722 4205 2739 4239
rect 2790 4205 2818 4239
rect 2858 4205 2892 4239
rect 2931 4205 2960 4239
rect 3170 4205 3200 4239
rect 3238 4205 3272 4239
rect 3313 4205 3340 4239
rect 3392 4205 3408 4239
rect 3471 4205 3476 4239
rect 3510 4205 3516 4239
rect 3578 4205 3595 4239
rect 3646 4205 3674 4239
rect 3714 4205 3748 4239
rect 3787 4205 3816 4239
rect 4026 4205 4056 4239
rect 4094 4205 4128 4239
rect 4169 4205 4196 4239
rect 4248 4205 4264 4239
rect 4327 4205 4332 4239
rect 4366 4205 4372 4239
rect 4434 4205 4451 4239
rect 4502 4205 4530 4239
rect 4570 4205 4604 4239
rect 4643 4205 4672 4239
rect 4882 4205 4912 4239
rect 4950 4205 4984 4239
rect 5025 4205 5052 4239
rect 5104 4205 5120 4239
rect 5183 4205 5188 4239
rect 5222 4205 5228 4239
rect 5290 4205 5307 4239
rect 5358 4205 5386 4239
rect 5426 4205 5460 4239
rect 5499 4205 5528 4239
rect 5738 4205 5768 4239
rect 5806 4205 5840 4239
rect 5881 4205 5908 4239
rect 5960 4205 5976 4239
rect 6039 4205 6044 4239
rect 6078 4205 6084 4239
rect 6146 4205 6163 4239
rect 6214 4205 6242 4239
rect 6282 4205 6316 4239
rect 6355 4205 6384 4239
rect 6594 4205 6624 4239
rect 6662 4205 6696 4239
rect 6737 4205 6764 4239
rect 6816 4205 6832 4239
rect 6895 4205 6900 4239
rect 6934 4205 6940 4239
rect 7002 4205 7019 4239
rect 7070 4205 7098 4239
rect 7138 4205 7172 4239
rect 7211 4205 7240 4239
rect 7450 4205 7480 4239
rect 7518 4205 7552 4239
rect 7593 4205 7620 4239
rect 7672 4205 7688 4239
rect 7751 4205 7756 4239
rect 7790 4205 7796 4239
rect 7858 4205 7875 4239
rect 7926 4205 7954 4239
rect 7994 4205 8028 4239
rect 8067 4205 8096 4239
rect 8306 4205 8336 4239
rect 8374 4205 8408 4239
rect 8449 4205 8476 4239
rect 8528 4205 8544 4239
rect 8607 4205 8612 4239
rect 8646 4205 8652 4239
rect 8714 4205 8731 4239
rect 8782 4205 8810 4239
rect 8850 4205 8884 4239
rect 8923 4205 8952 4239
rect 9162 4205 9192 4239
rect 9230 4205 9264 4239
rect 9305 4205 9332 4239
rect 9384 4205 9400 4239
rect 9463 4205 9468 4239
rect 9502 4205 9508 4239
rect 9570 4205 9587 4239
rect 9638 4205 9666 4239
rect 9706 4205 9740 4239
rect 9779 4205 9808 4239
rect 10018 4205 10048 4239
rect 10086 4205 10120 4239
rect 10161 4205 10188 4239
rect 10240 4205 10256 4239
rect 10319 4205 10324 4239
rect 10358 4205 10364 4239
rect 10426 4205 10443 4239
rect 10494 4205 10522 4239
rect 10562 4205 10596 4239
rect 10635 4205 10664 4239
rect 10856 4236 10872 4281
rect 10906 4236 10922 4281
rect 10856 4212 10922 4236
rect 344 4159 410 4178
rect 10856 4178 10872 4212
rect 10906 4178 10922 4212
rect 10856 4159 10922 4178
rect 344 4143 10922 4159
rect 344 4109 360 4143
rect 394 4139 429 4143
rect 463 4139 498 4143
rect 532 4139 567 4143
rect 601 4139 636 4143
rect 413 4109 429 4139
rect 486 4109 498 4139
rect 559 4109 567 4139
rect 632 4109 636 4139
rect 670 4139 705 4143
rect 670 4109 671 4139
rect 344 4105 379 4109
rect 413 4105 452 4109
rect 486 4105 525 4109
rect 559 4105 598 4109
rect 632 4105 671 4109
rect 739 4139 774 4143
rect 808 4139 843 4143
rect 877 4139 912 4143
rect 946 4139 981 4143
rect 1015 4139 1050 4143
rect 1084 4139 1119 4143
rect 1153 4139 1188 4143
rect 1222 4139 1257 4143
rect 739 4109 744 4139
rect 808 4109 817 4139
rect 877 4109 890 4139
rect 946 4109 963 4139
rect 1015 4109 1036 4139
rect 1084 4109 1109 4139
rect 1153 4109 1182 4139
rect 1222 4109 1255 4139
rect 1291 4109 1326 4143
rect 1360 4139 1395 4143
rect 1429 4139 1464 4143
rect 1498 4139 1533 4143
rect 1567 4139 1602 4143
rect 1636 4139 1671 4143
rect 1705 4139 1740 4143
rect 1774 4139 1809 4143
rect 1843 4139 1878 4143
rect 1362 4109 1395 4139
rect 1435 4109 1464 4139
rect 1508 4109 1533 4139
rect 1581 4109 1602 4139
rect 1654 4109 1671 4139
rect 1727 4109 1740 4139
rect 1800 4109 1809 4139
rect 1873 4109 1878 4139
rect 1912 4139 1947 4143
rect 705 4105 744 4109
rect 778 4105 817 4109
rect 851 4105 890 4109
rect 924 4105 963 4109
rect 997 4105 1036 4109
rect 1070 4105 1109 4109
rect 1143 4105 1182 4109
rect 1216 4105 1255 4109
rect 1289 4105 1328 4109
rect 1362 4105 1401 4109
rect 1435 4105 1474 4109
rect 1508 4105 1547 4109
rect 1581 4105 1620 4109
rect 1654 4105 1693 4109
rect 1727 4105 1766 4109
rect 1800 4105 1839 4109
rect 1873 4105 1912 4109
rect 1946 4109 1947 4139
rect 1981 4139 2016 4143
rect 2050 4139 2085 4143
rect 2119 4139 2154 4143
rect 2188 4139 2223 4143
rect 2257 4139 2292 4143
rect 2326 4139 2361 4143
rect 2395 4139 2430 4143
rect 2464 4139 2499 4143
rect 1981 4109 1985 4139
rect 2050 4109 2058 4139
rect 2119 4109 2131 4139
rect 2188 4109 2204 4139
rect 2257 4109 2277 4139
rect 2326 4109 2350 4139
rect 2395 4109 2423 4139
rect 2464 4109 2496 4139
rect 2533 4109 2568 4143
rect 2602 4139 2637 4143
rect 2671 4139 2706 4143
rect 2740 4139 2775 4143
rect 2809 4139 2844 4143
rect 2878 4139 2913 4143
rect 2947 4139 2982 4143
rect 3016 4139 3051 4143
rect 3085 4139 3120 4143
rect 3154 4139 3188 4143
rect 2603 4109 2637 4139
rect 2676 4109 2706 4139
rect 2749 4109 2775 4139
rect 2822 4109 2844 4139
rect 2895 4109 2913 4139
rect 2968 4109 2982 4139
rect 3041 4109 3051 4139
rect 3114 4109 3120 4139
rect 3187 4109 3188 4139
rect 3222 4139 3256 4143
rect 3290 4139 3324 4143
rect 3358 4139 3392 4143
rect 3426 4139 3460 4143
rect 3494 4139 3528 4143
rect 3562 4139 3596 4143
rect 3630 4139 3664 4143
rect 3222 4109 3226 4139
rect 3290 4109 3299 4139
rect 3358 4109 3372 4139
rect 3426 4109 3444 4139
rect 3494 4109 3516 4139
rect 3562 4109 3588 4139
rect 3630 4109 3660 4139
rect 3698 4109 3732 4143
rect 3766 4109 3800 4143
rect 3834 4139 3868 4143
rect 3902 4139 3936 4143
rect 3970 4139 4004 4143
rect 4038 4139 4072 4143
rect 4106 4139 4140 4143
rect 4174 4139 4208 4143
rect 4242 4139 4276 4143
rect 4310 4139 4344 4143
rect 3838 4109 3868 4139
rect 3910 4109 3936 4139
rect 3982 4109 4004 4139
rect 4054 4109 4072 4139
rect 4126 4109 4140 4139
rect 4198 4109 4208 4139
rect 4270 4109 4276 4139
rect 4342 4109 4344 4139
rect 4378 4139 4412 4143
rect 4446 4139 4480 4143
rect 4514 4139 4548 4143
rect 4582 4139 4616 4143
rect 4650 4139 4684 4143
rect 4718 4139 4752 4143
rect 4786 4139 4820 4143
rect 4854 4139 4888 4143
rect 4378 4109 4380 4139
rect 4446 4109 4452 4139
rect 4514 4109 4524 4139
rect 4582 4109 4596 4139
rect 4650 4109 4668 4139
rect 4718 4109 4740 4139
rect 4786 4109 4812 4139
rect 4854 4109 4884 4139
rect 4922 4109 4956 4143
rect 4990 4109 5024 4143
rect 5058 4139 5092 4143
rect 5126 4139 5160 4143
rect 5194 4139 5228 4143
rect 5262 4139 5296 4143
rect 5330 4139 5364 4143
rect 5398 4139 5432 4143
rect 5466 4139 5500 4143
rect 5534 4139 5568 4143
rect 5062 4109 5092 4139
rect 5134 4109 5160 4139
rect 5206 4109 5228 4139
rect 5278 4109 5296 4139
rect 5350 4109 5364 4139
rect 5422 4109 5432 4139
rect 5494 4109 5500 4139
rect 5566 4109 5568 4139
rect 5602 4139 5636 4143
rect 5670 4139 5704 4143
rect 5738 4139 5772 4143
rect 5806 4139 5840 4143
rect 5874 4139 5908 4143
rect 5942 4139 5976 4143
rect 6010 4139 6044 4143
rect 6078 4139 6112 4143
rect 5602 4109 5604 4139
rect 5670 4109 5676 4139
rect 5738 4109 5748 4139
rect 5806 4109 5820 4139
rect 5874 4109 5892 4139
rect 5942 4109 5964 4139
rect 6010 4109 6036 4139
rect 6078 4109 6108 4139
rect 6146 4109 6180 4143
rect 6214 4109 6248 4143
rect 6282 4139 6316 4143
rect 6350 4139 6384 4143
rect 6418 4139 6452 4143
rect 6486 4139 6520 4143
rect 6554 4139 6588 4143
rect 6622 4139 6656 4143
rect 6690 4139 6724 4143
rect 6758 4139 6792 4143
rect 6286 4109 6316 4139
rect 6358 4109 6384 4139
rect 6430 4109 6452 4139
rect 6502 4109 6520 4139
rect 6574 4109 6588 4139
rect 6646 4109 6656 4139
rect 6718 4109 6724 4139
rect 6790 4109 6792 4139
rect 6826 4139 6860 4143
rect 6894 4139 6928 4143
rect 6962 4139 6996 4143
rect 7030 4139 7064 4143
rect 7098 4139 7132 4143
rect 7166 4139 7200 4143
rect 7234 4139 7268 4143
rect 7302 4139 7336 4143
rect 6826 4109 6828 4139
rect 6894 4109 6900 4139
rect 6962 4109 6972 4139
rect 7030 4109 7044 4139
rect 7098 4109 7116 4139
rect 7166 4109 7188 4139
rect 7234 4109 7260 4139
rect 7302 4109 7332 4139
rect 7370 4109 7404 4143
rect 7438 4109 7472 4143
rect 7506 4139 7540 4143
rect 7574 4139 7608 4143
rect 7642 4139 7676 4143
rect 7710 4139 7744 4143
rect 7778 4139 7812 4143
rect 7846 4139 7880 4143
rect 7914 4139 7948 4143
rect 7982 4139 8016 4143
rect 7510 4109 7540 4139
rect 7582 4109 7608 4139
rect 7654 4109 7676 4139
rect 7726 4109 7744 4139
rect 7798 4109 7812 4139
rect 7870 4109 7880 4139
rect 7942 4109 7948 4139
rect 8014 4109 8016 4139
rect 8050 4139 8084 4143
rect 8118 4139 8152 4143
rect 8186 4139 8220 4143
rect 8254 4139 8288 4143
rect 8322 4139 8356 4143
rect 8390 4139 8424 4143
rect 8458 4139 8492 4143
rect 8526 4139 8560 4143
rect 8050 4109 8052 4139
rect 8118 4109 8124 4139
rect 8186 4109 8196 4139
rect 8254 4109 8268 4139
rect 8322 4109 8340 4139
rect 8390 4109 8412 4139
rect 8458 4109 8484 4139
rect 8526 4109 8556 4139
rect 8594 4109 8628 4143
rect 8662 4109 8696 4143
rect 8730 4139 8764 4143
rect 8798 4139 8832 4143
rect 8866 4139 8900 4143
rect 8934 4139 8968 4143
rect 9002 4139 9036 4143
rect 9070 4139 9104 4143
rect 9138 4139 9172 4143
rect 9206 4139 9240 4143
rect 8734 4109 8764 4139
rect 8806 4109 8832 4139
rect 8878 4109 8900 4139
rect 8950 4109 8968 4139
rect 9022 4109 9036 4139
rect 9094 4109 9104 4139
rect 9166 4109 9172 4139
rect 9238 4109 9240 4139
rect 9274 4139 9308 4143
rect 9342 4139 9376 4143
rect 9410 4139 9444 4143
rect 9478 4139 9512 4143
rect 9546 4139 9580 4143
rect 9614 4139 9648 4143
rect 9682 4139 9716 4143
rect 9750 4139 9784 4143
rect 9274 4109 9276 4139
rect 9342 4109 9348 4139
rect 9410 4109 9420 4139
rect 9478 4109 9492 4139
rect 9546 4109 9564 4139
rect 9614 4109 9636 4139
rect 9682 4109 9708 4139
rect 9750 4109 9780 4139
rect 9818 4109 9852 4143
rect 9886 4109 9920 4143
rect 9954 4139 9988 4143
rect 10022 4139 10056 4143
rect 10090 4139 10124 4143
rect 10158 4139 10192 4143
rect 10226 4139 10260 4143
rect 10294 4139 10328 4143
rect 10362 4139 10396 4143
rect 10430 4139 10464 4143
rect 9958 4109 9988 4139
rect 10030 4109 10056 4139
rect 10102 4109 10124 4139
rect 10174 4109 10192 4139
rect 10246 4109 10260 4139
rect 10318 4109 10328 4139
rect 10390 4109 10396 4139
rect 10462 4109 10464 4139
rect 10498 4139 10532 4143
rect 10566 4139 10600 4143
rect 10634 4139 10668 4143
rect 10702 4139 10736 4143
rect 10770 4139 10804 4143
rect 10838 4139 10872 4143
rect 10498 4109 10500 4139
rect 10566 4109 10572 4139
rect 10634 4109 10644 4139
rect 10702 4109 10716 4139
rect 10770 4109 10788 4139
rect 10838 4109 10860 4139
rect 10906 4109 10922 4143
rect 1946 4105 1985 4109
rect 2019 4105 2058 4109
rect 2092 4105 2131 4109
rect 2165 4105 2204 4109
rect 2238 4105 2277 4109
rect 2311 4105 2350 4109
rect 2384 4105 2423 4109
rect 2457 4105 2496 4109
rect 2530 4105 2569 4109
rect 2603 4105 2642 4109
rect 2676 4105 2715 4109
rect 2749 4105 2788 4109
rect 2822 4105 2861 4109
rect 2895 4105 2934 4109
rect 2968 4105 3007 4109
rect 3041 4105 3080 4109
rect 3114 4105 3153 4109
rect 3187 4105 3226 4109
rect 3260 4105 3299 4109
rect 3333 4105 3372 4109
rect 3406 4105 3444 4109
rect 3478 4105 3516 4109
rect 3550 4105 3588 4109
rect 3622 4105 3660 4109
rect 3694 4105 3732 4109
rect 3766 4105 3804 4109
rect 3838 4105 3876 4109
rect 3910 4105 3948 4109
rect 3982 4105 4020 4109
rect 4054 4105 4092 4109
rect 4126 4105 4164 4109
rect 4198 4105 4236 4109
rect 4270 4105 4308 4109
rect 4342 4105 4380 4109
rect 4414 4105 4452 4109
rect 4486 4105 4524 4109
rect 4558 4105 4596 4109
rect 4630 4105 4668 4109
rect 4702 4105 4740 4109
rect 4774 4105 4812 4109
rect 4846 4105 4884 4109
rect 4918 4105 4956 4109
rect 4990 4105 5028 4109
rect 5062 4105 5100 4109
rect 5134 4105 5172 4109
rect 5206 4105 5244 4109
rect 5278 4105 5316 4109
rect 5350 4105 5388 4109
rect 5422 4105 5460 4109
rect 5494 4105 5532 4109
rect 5566 4105 5604 4109
rect 5638 4105 5676 4109
rect 5710 4105 5748 4109
rect 5782 4105 5820 4109
rect 5854 4105 5892 4109
rect 5926 4105 5964 4109
rect 5998 4105 6036 4109
rect 6070 4105 6108 4109
rect 6142 4105 6180 4109
rect 6214 4105 6252 4109
rect 6286 4105 6324 4109
rect 6358 4105 6396 4109
rect 6430 4105 6468 4109
rect 6502 4105 6540 4109
rect 6574 4105 6612 4109
rect 6646 4105 6684 4109
rect 6718 4105 6756 4109
rect 6790 4105 6828 4109
rect 6862 4105 6900 4109
rect 6934 4105 6972 4109
rect 7006 4105 7044 4109
rect 7078 4105 7116 4109
rect 7150 4105 7188 4109
rect 7222 4105 7260 4109
rect 7294 4105 7332 4109
rect 7366 4105 7404 4109
rect 7438 4105 7476 4109
rect 7510 4105 7548 4109
rect 7582 4105 7620 4109
rect 7654 4105 7692 4109
rect 7726 4105 7764 4109
rect 7798 4105 7836 4109
rect 7870 4105 7908 4109
rect 7942 4105 7980 4109
rect 8014 4105 8052 4109
rect 8086 4105 8124 4109
rect 8158 4105 8196 4109
rect 8230 4105 8268 4109
rect 8302 4105 8340 4109
rect 8374 4105 8412 4109
rect 8446 4105 8484 4109
rect 8518 4105 8556 4109
rect 8590 4105 8628 4109
rect 8662 4105 8700 4109
rect 8734 4105 8772 4109
rect 8806 4105 8844 4109
rect 8878 4105 8916 4109
rect 8950 4105 8988 4109
rect 9022 4105 9060 4109
rect 9094 4105 9132 4109
rect 9166 4105 9204 4109
rect 9238 4105 9276 4109
rect 9310 4105 9348 4109
rect 9382 4105 9420 4109
rect 9454 4105 9492 4109
rect 9526 4105 9564 4109
rect 9598 4105 9636 4109
rect 9670 4105 9708 4109
rect 9742 4105 9780 4109
rect 9814 4105 9852 4109
rect 9886 4105 9924 4109
rect 9958 4105 9996 4109
rect 10030 4105 10068 4109
rect 10102 4105 10140 4109
rect 10174 4105 10212 4109
rect 10246 4105 10284 4109
rect 10318 4105 10356 4109
rect 10390 4105 10428 4109
rect 10462 4105 10500 4109
rect 10534 4105 10572 4109
rect 10606 4105 10644 4109
rect 10678 4105 10716 4109
rect 10750 4105 10788 4109
rect 10822 4105 10860 4109
rect 10894 4105 10922 4109
rect 344 4093 10922 4105
rect 11482 5813 11564 5848
rect 11660 5854 11694 5888
rect 14562 5854 14596 5888
rect 14740 5879 16033 5888
rect 11658 5838 11696 5854
rect 14528 5838 14630 5854
rect 14740 5845 14774 5879
rect 14808 5845 14844 5879
rect 14878 5845 14914 5879
rect 14948 5845 14984 5879
rect 15018 5845 15054 5879
rect 15088 5845 15124 5879
rect 15158 5845 15194 5879
rect 15228 5845 15264 5879
rect 15298 5845 15334 5879
rect 15368 5845 15404 5879
rect 15438 5845 15474 5879
rect 15508 5845 15544 5879
rect 15578 5845 15614 5879
rect 15648 5845 15684 5879
rect 15718 5850 15754 5879
rect 15788 5850 15824 5879
rect 15718 5845 15733 5850
rect 15788 5845 15819 5850
rect 15858 5845 15894 5879
rect 15928 5850 15964 5879
rect 15998 5850 16033 5879
rect 15939 5845 15964 5850
rect 11482 5779 11506 5813
rect 11540 5779 11564 5813
rect 11482 5744 11564 5779
rect 14740 5816 15733 5845
rect 15767 5816 15819 5845
rect 15853 5816 15905 5845
rect 15939 5816 15991 5845
rect 16025 5816 16033 5850
rect 14740 5810 16033 5816
rect 14740 5776 14774 5810
rect 14808 5776 14844 5810
rect 14878 5776 14914 5810
rect 14948 5776 14984 5810
rect 15018 5776 15054 5810
rect 15088 5776 15124 5810
rect 15158 5776 15194 5810
rect 15228 5776 15264 5810
rect 15298 5776 15334 5810
rect 15368 5776 15404 5810
rect 15438 5776 15474 5810
rect 15508 5776 15544 5810
rect 15578 5776 15614 5810
rect 15648 5776 15684 5810
rect 15718 5778 15754 5810
rect 15788 5778 15824 5810
rect 15718 5776 15733 5778
rect 15788 5776 15819 5778
rect 15858 5776 15894 5810
rect 15928 5778 15964 5810
rect 15998 5778 16033 5810
rect 15939 5776 15964 5778
rect 11482 5710 11506 5744
rect 11540 5710 11564 5744
rect 11626 5734 11728 5750
rect 14528 5734 14630 5750
rect 14740 5744 15733 5776
rect 15767 5744 15819 5776
rect 15853 5744 15905 5776
rect 15939 5744 15991 5776
rect 16025 5744 16033 5778
rect 14740 5741 16033 5744
rect 11482 5675 11564 5710
rect 11660 5700 11694 5734
rect 14562 5700 14596 5734
rect 14740 5707 14774 5741
rect 14808 5707 14844 5741
rect 14878 5707 14914 5741
rect 14948 5707 14984 5741
rect 15018 5707 15054 5741
rect 15088 5707 15124 5741
rect 15158 5707 15194 5741
rect 15228 5707 15264 5741
rect 15298 5707 15334 5741
rect 15368 5707 15404 5741
rect 15438 5707 15474 5741
rect 15508 5707 15544 5741
rect 15578 5707 15614 5741
rect 15648 5707 15684 5741
rect 15718 5707 15754 5741
rect 15788 5707 15824 5741
rect 15858 5707 15894 5741
rect 15928 5707 15964 5741
rect 15998 5707 16033 5741
rect 14740 5706 16033 5707
rect 11626 5684 11728 5700
rect 14528 5684 14630 5700
rect 11482 5641 11506 5675
rect 11540 5641 11564 5675
rect 11482 5606 11564 5641
rect 11482 5599 11506 5606
rect 11482 5565 11500 5599
rect 11540 5572 11564 5606
rect 14740 5672 15733 5706
rect 15767 5672 15819 5706
rect 15853 5672 15905 5706
rect 15939 5672 15991 5706
rect 16025 5672 16033 5706
rect 14740 5638 14774 5672
rect 14808 5638 14844 5672
rect 14878 5638 14914 5672
rect 14948 5638 14984 5672
rect 15018 5638 15054 5672
rect 15088 5638 15124 5672
rect 15158 5638 15194 5672
rect 15228 5638 15264 5672
rect 15298 5638 15334 5672
rect 15368 5638 15404 5672
rect 15438 5638 15474 5672
rect 15508 5638 15544 5672
rect 15578 5638 15614 5672
rect 15648 5638 15684 5672
rect 15718 5638 15754 5672
rect 15788 5638 15824 5672
rect 15858 5638 15894 5672
rect 15928 5638 15964 5672
rect 15998 5638 16033 5672
rect 14740 5634 16033 5638
rect 14740 5603 15733 5634
rect 15767 5603 15819 5634
rect 15853 5603 15905 5634
rect 15939 5603 15991 5634
rect 11626 5580 11728 5596
rect 14528 5580 14630 5596
rect 11534 5565 11564 5572
rect 11482 5537 11564 5565
rect 11660 5546 11694 5580
rect 14562 5546 14596 5580
rect 14740 5569 14774 5603
rect 14808 5569 14844 5603
rect 14878 5569 14914 5603
rect 14948 5569 14984 5603
rect 15018 5569 15054 5603
rect 15088 5569 15124 5603
rect 15158 5569 15194 5603
rect 15228 5569 15264 5603
rect 15298 5569 15334 5603
rect 15368 5569 15404 5603
rect 15438 5569 15474 5603
rect 15508 5569 15544 5603
rect 15578 5569 15614 5603
rect 15648 5569 15684 5603
rect 15718 5600 15733 5603
rect 15788 5600 15819 5603
rect 15718 5569 15754 5600
rect 15788 5569 15824 5600
rect 15858 5569 15894 5603
rect 15939 5600 15964 5603
rect 16025 5600 16033 5634
rect 15928 5569 15964 5600
rect 15998 5569 16033 5600
rect 14740 5562 16033 5569
rect 11482 5525 11506 5537
rect 11482 5491 11500 5525
rect 11540 5503 11564 5537
rect 11626 5530 11728 5546
rect 14528 5530 14630 5546
rect 14740 5534 15733 5562
rect 15767 5534 15819 5562
rect 15853 5534 15905 5562
rect 15939 5534 15991 5562
rect 11534 5491 11564 5503
rect 11482 5468 11564 5491
rect 11482 5451 11506 5468
rect 11482 5417 11500 5451
rect 11540 5434 11564 5468
rect 14740 5500 14774 5534
rect 14808 5500 14844 5534
rect 14878 5500 14914 5534
rect 14948 5500 14984 5534
rect 15018 5500 15054 5534
rect 15088 5500 15124 5534
rect 15158 5500 15194 5534
rect 15228 5500 15264 5534
rect 15298 5500 15334 5534
rect 15368 5500 15404 5534
rect 15438 5500 15474 5534
rect 15508 5500 15544 5534
rect 15578 5500 15614 5534
rect 15648 5500 15684 5534
rect 15718 5528 15733 5534
rect 15788 5528 15819 5534
rect 15718 5500 15754 5528
rect 15788 5500 15824 5528
rect 15858 5500 15894 5534
rect 15939 5528 15964 5534
rect 16025 5528 16033 5562
rect 15928 5500 15964 5528
rect 15998 5500 16033 5528
rect 14740 5490 16033 5500
rect 14740 5465 15733 5490
rect 15767 5465 15819 5490
rect 15853 5465 15905 5490
rect 15939 5465 15991 5490
rect 11534 5417 11564 5434
rect 11626 5426 11728 5442
rect 14528 5426 14630 5442
rect 14740 5431 14774 5465
rect 14808 5431 14844 5465
rect 14878 5431 14914 5465
rect 14948 5431 14984 5465
rect 15018 5431 15054 5465
rect 15088 5431 15124 5465
rect 15158 5431 15194 5465
rect 15228 5431 15264 5465
rect 15298 5431 15334 5465
rect 15368 5431 15404 5465
rect 15438 5431 15474 5465
rect 15508 5431 15544 5465
rect 15578 5431 15614 5465
rect 15648 5431 15684 5465
rect 15718 5456 15733 5465
rect 15788 5456 15819 5465
rect 15718 5431 15754 5456
rect 15788 5431 15824 5456
rect 15858 5431 15894 5465
rect 15939 5456 15964 5465
rect 16025 5456 16033 5490
rect 15928 5431 15964 5456
rect 15998 5431 16033 5456
rect 11482 5399 11564 5417
rect 11482 5377 11506 5399
rect 11482 5343 11500 5377
rect 11540 5365 11564 5399
rect 11660 5392 11694 5426
rect 14562 5392 14596 5426
rect 14740 5418 16033 5431
rect 14740 5396 15733 5418
rect 15767 5396 15819 5418
rect 15853 5396 15905 5418
rect 15939 5396 15991 5418
rect 11626 5376 11728 5392
rect 14528 5376 14630 5392
rect 11534 5343 11564 5365
rect 11482 5330 11564 5343
rect 11482 5303 11506 5330
rect 11482 5269 11500 5303
rect 11540 5296 11564 5330
rect 11534 5269 11564 5296
rect 14740 5362 14774 5396
rect 14808 5362 14844 5396
rect 14878 5362 14914 5396
rect 14948 5362 14984 5396
rect 15018 5362 15054 5396
rect 15088 5362 15124 5396
rect 15158 5362 15194 5396
rect 15228 5362 15264 5396
rect 15298 5362 15334 5396
rect 15368 5362 15404 5396
rect 15438 5362 15474 5396
rect 15508 5362 15544 5396
rect 15578 5362 15614 5396
rect 15648 5362 15684 5396
rect 15718 5384 15733 5396
rect 15788 5384 15819 5396
rect 15718 5362 15754 5384
rect 15788 5362 15824 5384
rect 15858 5362 15894 5396
rect 15939 5384 15964 5396
rect 16025 5384 16033 5418
rect 15928 5362 15964 5384
rect 15998 5362 16033 5384
rect 14740 5346 16033 5362
rect 14740 5327 15733 5346
rect 15767 5327 15819 5346
rect 15853 5327 15905 5346
rect 15939 5327 15991 5346
rect 14740 5293 14774 5327
rect 14808 5293 14844 5327
rect 14878 5293 14914 5327
rect 14948 5293 14984 5327
rect 15018 5293 15054 5327
rect 15088 5293 15124 5327
rect 15158 5293 15194 5327
rect 15228 5293 15264 5327
rect 15298 5293 15334 5327
rect 15368 5293 15404 5327
rect 15438 5293 15474 5327
rect 15508 5293 15544 5327
rect 15578 5293 15614 5327
rect 15648 5293 15684 5327
rect 15718 5312 15733 5327
rect 15788 5312 15819 5327
rect 15718 5293 15754 5312
rect 15788 5293 15824 5312
rect 15858 5293 15894 5327
rect 15939 5312 15964 5327
rect 16025 5312 16033 5346
rect 15928 5293 15964 5312
rect 15998 5293 16033 5312
rect 11626 5272 11728 5288
rect 14528 5272 14630 5288
rect 14740 5274 16033 5293
rect 11482 5261 11564 5269
rect 11482 5229 11506 5261
rect 11482 5195 11500 5229
rect 11540 5227 11564 5261
rect 11660 5238 11694 5272
rect 14562 5238 14596 5272
rect 14740 5258 15733 5274
rect 15767 5258 15819 5274
rect 15853 5258 15905 5274
rect 15939 5258 15991 5274
rect 11534 5195 11564 5227
rect 11626 5222 11728 5238
rect 14528 5222 14630 5238
rect 14740 5224 14774 5258
rect 14808 5224 14844 5258
rect 14878 5224 14914 5258
rect 14948 5224 14984 5258
rect 15018 5224 15054 5258
rect 15088 5224 15124 5258
rect 15158 5224 15194 5258
rect 15228 5224 15264 5258
rect 15298 5224 15334 5258
rect 15368 5224 15404 5258
rect 15438 5224 15474 5258
rect 15508 5224 15544 5258
rect 15578 5224 15614 5258
rect 15648 5224 15684 5258
rect 15718 5240 15733 5258
rect 15788 5240 15819 5258
rect 15718 5224 15754 5240
rect 15788 5224 15824 5240
rect 15858 5224 15894 5258
rect 15939 5240 15964 5258
rect 16025 5240 16033 5274
rect 15928 5224 15964 5240
rect 15998 5224 16033 5240
rect 11482 5192 11564 5195
rect 11482 5158 11506 5192
rect 11540 5158 11564 5192
rect 11482 5155 11564 5158
rect 11482 5121 11500 5155
rect 11534 5123 11564 5155
rect 14740 5202 16033 5224
rect 14740 5190 15733 5202
rect 15767 5190 15819 5202
rect 15853 5190 15905 5202
rect 15939 5190 15991 5202
rect 14740 5156 14774 5190
rect 14808 5156 14844 5190
rect 14878 5156 14914 5190
rect 14948 5156 14984 5190
rect 15018 5156 15054 5190
rect 15088 5156 15124 5190
rect 15158 5156 15194 5190
rect 15228 5156 15264 5190
rect 15298 5156 15334 5190
rect 15368 5156 15404 5190
rect 15438 5156 15474 5190
rect 15508 5156 15544 5190
rect 15578 5156 15614 5190
rect 15648 5156 15684 5190
rect 15718 5168 15733 5190
rect 15788 5168 15819 5190
rect 15718 5156 15754 5168
rect 15788 5156 15824 5168
rect 15858 5156 15894 5190
rect 15939 5168 15964 5190
rect 16025 5168 16033 5202
rect 15928 5156 15964 5168
rect 15998 5156 16033 5168
rect 11482 5089 11506 5121
rect 11540 5089 11564 5123
rect 11626 5118 11728 5134
rect 14528 5118 14630 5134
rect 14740 5130 16033 5156
rect 14740 5122 15733 5130
rect 15767 5122 15819 5130
rect 15853 5122 15905 5130
rect 15939 5122 15991 5130
rect 11482 5081 11564 5089
rect 11660 5084 11694 5118
rect 14562 5084 14596 5118
rect 14740 5088 14774 5122
rect 14808 5088 14844 5122
rect 14878 5088 14914 5122
rect 14948 5088 14984 5122
rect 15018 5088 15054 5122
rect 15088 5088 15124 5122
rect 15158 5088 15194 5122
rect 15228 5088 15264 5122
rect 15298 5088 15334 5122
rect 15368 5088 15404 5122
rect 15438 5088 15474 5122
rect 15508 5088 15544 5122
rect 15578 5088 15614 5122
rect 15648 5088 15684 5122
rect 15718 5096 15733 5122
rect 15788 5096 15819 5122
rect 15718 5088 15754 5096
rect 15788 5088 15824 5096
rect 15858 5088 15894 5122
rect 15939 5096 15964 5122
rect 16025 5096 16033 5130
rect 15928 5088 15964 5096
rect 15998 5088 16033 5096
rect 11482 5047 11500 5081
rect 11534 5054 11564 5081
rect 11626 5068 11728 5084
rect 14528 5068 14630 5084
rect 11482 5020 11506 5047
rect 11540 5020 11564 5054
rect 11482 5007 11564 5020
rect 11482 4973 11500 5007
rect 11534 4985 11564 5007
rect 11482 4951 11506 4973
rect 11540 4951 11564 4985
rect 14740 5058 16033 5088
rect 14740 5054 15733 5058
rect 15767 5054 15819 5058
rect 15853 5054 15905 5058
rect 15939 5054 15991 5058
rect 14740 5020 14774 5054
rect 14808 5020 14844 5054
rect 14878 5020 14914 5054
rect 14948 5020 14984 5054
rect 15018 5020 15054 5054
rect 15088 5020 15124 5054
rect 15158 5020 15194 5054
rect 15228 5020 15264 5054
rect 15298 5020 15334 5054
rect 15368 5020 15404 5054
rect 15438 5020 15474 5054
rect 15508 5020 15544 5054
rect 15578 5020 15614 5054
rect 15648 5020 15684 5054
rect 15718 5024 15733 5054
rect 15788 5024 15819 5054
rect 15718 5020 15754 5024
rect 15788 5020 15824 5024
rect 15858 5020 15894 5054
rect 15939 5024 15964 5054
rect 16025 5024 16033 5058
rect 15928 5020 15964 5024
rect 15998 5020 16033 5024
rect 14740 4986 16033 5020
rect 11626 4964 11728 4980
rect 14528 4964 14630 4980
rect 11482 4933 11564 4951
rect 11482 4899 11500 4933
rect 11534 4916 11564 4933
rect 11660 4930 11694 4964
rect 14562 4930 14596 4964
rect 14740 4952 14774 4986
rect 14808 4952 14844 4986
rect 14878 4952 14914 4986
rect 14948 4952 14984 4986
rect 15018 4952 15054 4986
rect 15088 4952 15124 4986
rect 15158 4952 15194 4986
rect 15228 4952 15264 4986
rect 15298 4952 15334 4986
rect 15368 4952 15404 4986
rect 15438 4952 15474 4986
rect 15508 4952 15544 4986
rect 15578 4952 15614 4986
rect 15648 4952 15684 4986
rect 15718 4952 15733 4986
rect 15788 4952 15819 4986
rect 15858 4952 15894 4986
rect 15939 4952 15964 4986
rect 16025 4952 16033 4986
rect 11482 4882 11506 4899
rect 11540 4882 11564 4916
rect 11626 4914 11728 4930
rect 14528 4914 14630 4930
rect 14740 4918 16033 4952
rect 11482 4859 11564 4882
rect 11482 4825 11500 4859
rect 11534 4847 11564 4859
rect 11482 4813 11506 4825
rect 11540 4813 11564 4847
rect 14740 4884 14774 4918
rect 14808 4884 14844 4918
rect 14878 4884 14914 4918
rect 14948 4884 14984 4918
rect 15018 4884 15054 4918
rect 15088 4884 15124 4918
rect 15158 4884 15194 4918
rect 15228 4884 15264 4918
rect 15298 4884 15334 4918
rect 15368 4884 15404 4918
rect 15438 4884 15474 4918
rect 15508 4884 15544 4918
rect 15578 4884 15614 4918
rect 15648 4884 15684 4918
rect 15718 4914 15754 4918
rect 15788 4914 15824 4918
rect 15718 4884 15733 4914
rect 15788 4884 15819 4914
rect 15858 4884 15894 4918
rect 15928 4914 15964 4918
rect 15998 4914 16033 4918
rect 15939 4884 15964 4914
rect 14740 4880 15733 4884
rect 15767 4880 15819 4884
rect 15853 4880 15905 4884
rect 15939 4880 15991 4884
rect 16025 4880 16033 4914
rect 14740 4850 16033 4880
rect 11482 4786 11564 4813
rect 11626 4810 11728 4826
rect 14528 4810 14630 4826
rect 14740 4816 14774 4850
rect 14808 4816 14844 4850
rect 14878 4816 14914 4850
rect 14948 4816 14984 4850
rect 15018 4816 15054 4850
rect 15088 4816 15124 4850
rect 15158 4816 15194 4850
rect 15228 4816 15264 4850
rect 15298 4816 15334 4850
rect 15368 4816 15404 4850
rect 15438 4816 15474 4850
rect 15508 4816 15544 4850
rect 15578 4816 15614 4850
rect 15648 4816 15684 4850
rect 15718 4842 15754 4850
rect 15788 4842 15824 4850
rect 15718 4816 15733 4842
rect 15788 4816 15819 4842
rect 15858 4816 15894 4850
rect 15928 4842 15964 4850
rect 15998 4842 16033 4850
rect 15939 4816 15964 4842
rect 11482 4752 11500 4786
rect 11534 4778 11564 4786
rect 11482 4744 11506 4752
rect 11540 4744 11564 4778
rect 11660 4776 11694 4810
rect 14562 4776 14596 4810
rect 14740 4808 15733 4816
rect 15767 4808 15819 4816
rect 15853 4808 15905 4816
rect 15939 4808 15991 4816
rect 16025 4808 16033 4842
rect 14740 4782 16033 4808
rect 11626 4760 11728 4776
rect 14528 4760 14630 4776
rect 11482 4713 11564 4744
rect 11482 4679 11500 4713
rect 11534 4709 11564 4713
rect 11482 4675 11506 4679
rect 11540 4675 11564 4709
rect 11482 4640 11564 4675
rect 14740 4748 14774 4782
rect 14808 4748 14844 4782
rect 14878 4748 14914 4782
rect 14948 4748 14984 4782
rect 15018 4748 15054 4782
rect 15088 4748 15124 4782
rect 15158 4748 15194 4782
rect 15228 4748 15264 4782
rect 15298 4748 15334 4782
rect 15368 4748 15404 4782
rect 15438 4748 15474 4782
rect 15508 4748 15544 4782
rect 15578 4748 15614 4782
rect 15648 4748 15684 4782
rect 15718 4770 15754 4782
rect 15788 4770 15824 4782
rect 15718 4748 15733 4770
rect 15788 4748 15819 4770
rect 15858 4748 15894 4782
rect 15928 4770 15964 4782
rect 15998 4770 16033 4782
rect 15939 4748 15964 4770
rect 14740 4736 15733 4748
rect 15767 4736 15819 4748
rect 15853 4736 15905 4748
rect 15939 4736 15991 4748
rect 16025 4736 16033 4770
rect 14740 4714 16033 4736
rect 14740 4680 14774 4714
rect 14808 4680 14844 4714
rect 14878 4680 14914 4714
rect 14948 4680 14984 4714
rect 15018 4680 15054 4714
rect 15088 4680 15124 4714
rect 15158 4680 15194 4714
rect 15228 4680 15264 4714
rect 15298 4680 15334 4714
rect 15368 4680 15404 4714
rect 15438 4680 15474 4714
rect 15508 4680 15544 4714
rect 15578 4680 15614 4714
rect 15648 4680 15684 4714
rect 15718 4698 15754 4714
rect 15788 4698 15824 4714
rect 15718 4680 15733 4698
rect 15788 4680 15819 4698
rect 15858 4680 15894 4714
rect 15928 4698 15964 4714
rect 15998 4698 16033 4714
rect 15939 4680 15964 4698
rect 11626 4656 11728 4672
rect 14528 4656 14630 4672
rect 14740 4664 15733 4680
rect 15767 4664 15819 4680
rect 15853 4664 15905 4680
rect 15939 4664 15991 4680
rect 16025 4664 16033 4698
rect 11482 4606 11500 4640
rect 11540 4606 11564 4640
rect 11660 4622 11694 4656
rect 14562 4622 14596 4656
rect 14740 4646 16033 4664
rect 11626 4606 11728 4622
rect 14528 4606 14630 4622
rect 14740 4612 14774 4646
rect 14808 4612 14844 4646
rect 14878 4612 14914 4646
rect 14948 4612 14984 4646
rect 15018 4612 15054 4646
rect 15088 4612 15124 4646
rect 15158 4612 15194 4646
rect 15228 4612 15264 4646
rect 15298 4612 15334 4646
rect 15368 4612 15404 4646
rect 15438 4612 15474 4646
rect 15508 4612 15544 4646
rect 15578 4612 15614 4646
rect 15648 4612 15684 4646
rect 15718 4626 15754 4646
rect 15788 4626 15824 4646
rect 15718 4612 15733 4626
rect 15788 4612 15819 4626
rect 15858 4612 15894 4646
rect 15928 4626 15964 4646
rect 15998 4626 16033 4646
rect 15939 4612 15964 4626
rect 11482 4571 11564 4606
rect 11482 4567 11506 4571
rect 11482 4533 11500 4567
rect 11540 4537 11564 4571
rect 11534 4533 11564 4537
rect 11482 4502 11564 4533
rect 14740 4592 15733 4612
rect 15767 4592 15819 4612
rect 15853 4592 15905 4612
rect 15939 4592 15991 4612
rect 16025 4592 16033 4626
rect 14740 4578 16033 4592
rect 14740 4544 14774 4578
rect 14808 4544 14844 4578
rect 14878 4544 14914 4578
rect 14948 4544 14984 4578
rect 15018 4544 15054 4578
rect 15088 4544 15124 4578
rect 15158 4544 15194 4578
rect 15228 4544 15264 4578
rect 15298 4544 15334 4578
rect 15368 4544 15404 4578
rect 15438 4544 15474 4578
rect 15508 4544 15544 4578
rect 15578 4544 15614 4578
rect 15648 4544 15684 4578
rect 15718 4554 15754 4578
rect 15788 4554 15824 4578
rect 15718 4544 15733 4554
rect 15788 4544 15819 4554
rect 15858 4544 15894 4578
rect 15928 4554 15964 4578
rect 15998 4554 16033 4578
rect 15939 4544 15964 4554
rect 14740 4520 15733 4544
rect 15767 4520 15819 4544
rect 15853 4520 15905 4544
rect 15939 4520 15991 4544
rect 16025 4520 16033 4554
rect 11626 4502 11728 4518
rect 14528 4502 14630 4518
rect 14740 4510 16033 4520
rect 11482 4494 11506 4502
rect 11482 4460 11500 4494
rect 11540 4468 11564 4502
rect 11660 4468 11694 4502
rect 14562 4468 14596 4502
rect 14740 4476 14774 4510
rect 14808 4476 14844 4510
rect 14878 4476 14914 4510
rect 14948 4476 14984 4510
rect 15018 4476 15054 4510
rect 15088 4476 15124 4510
rect 15158 4476 15194 4510
rect 15228 4476 15264 4510
rect 15298 4476 15334 4510
rect 15368 4476 15404 4510
rect 15438 4476 15474 4510
rect 15508 4476 15544 4510
rect 15578 4476 15614 4510
rect 15648 4476 15684 4510
rect 15718 4482 15754 4510
rect 15788 4482 15824 4510
rect 15718 4476 15733 4482
rect 15788 4476 15819 4482
rect 15858 4476 15894 4510
rect 15928 4482 15964 4510
rect 15998 4482 16033 4510
rect 15939 4476 15964 4482
rect 11534 4460 11564 4468
rect 11482 4433 11564 4460
rect 11626 4452 11728 4468
rect 14528 4452 14630 4468
rect 11482 4421 11506 4433
rect 11482 4387 11500 4421
rect 11540 4399 11564 4433
rect 11534 4387 11564 4399
rect 11482 4364 11564 4387
rect 14740 4448 15733 4476
rect 15767 4448 15819 4476
rect 15853 4448 15905 4476
rect 15939 4448 15991 4476
rect 16025 4448 16033 4482
rect 14740 4442 16033 4448
rect 14740 4408 14774 4442
rect 14808 4408 14844 4442
rect 14878 4408 14914 4442
rect 14948 4408 14984 4442
rect 15018 4408 15054 4442
rect 15088 4408 15124 4442
rect 15158 4408 15194 4442
rect 15228 4408 15264 4442
rect 15298 4408 15334 4442
rect 15368 4408 15404 4442
rect 15438 4408 15474 4442
rect 15508 4408 15544 4442
rect 15578 4408 15614 4442
rect 15648 4408 15684 4442
rect 15718 4410 15754 4442
rect 15788 4410 15824 4442
rect 15718 4408 15733 4410
rect 15788 4408 15819 4410
rect 15858 4408 15894 4442
rect 15928 4410 15964 4442
rect 15998 4410 16033 4442
rect 15939 4408 15964 4410
rect 14740 4376 15733 4408
rect 15767 4376 15819 4408
rect 15853 4376 15905 4408
rect 15939 4376 15991 4408
rect 16025 4376 16033 4410
rect 14740 4374 16033 4376
rect 11482 4348 11506 4364
rect 11482 4314 11500 4348
rect 11540 4330 11564 4364
rect 11626 4348 11728 4364
rect 14528 4348 14630 4364
rect 11534 4314 11564 4330
rect 11660 4314 11694 4348
rect 14562 4314 14596 4348
rect 14740 4340 14774 4374
rect 14808 4340 14844 4374
rect 14878 4340 14914 4374
rect 14948 4340 14984 4374
rect 15018 4340 15054 4374
rect 15088 4340 15124 4374
rect 15158 4340 15194 4374
rect 15228 4340 15264 4374
rect 15298 4340 15334 4374
rect 15368 4340 15404 4374
rect 15438 4340 15474 4374
rect 15508 4340 15544 4374
rect 15578 4340 15614 4374
rect 15648 4340 15684 4374
rect 15718 4340 15754 4374
rect 15788 4340 15824 4374
rect 15858 4340 15894 4374
rect 15928 4340 15964 4374
rect 15998 4340 16033 4374
rect 14740 4338 16033 4340
rect 11482 4295 11564 4314
rect 11626 4298 11728 4314
rect 14528 4298 14630 4314
rect 14740 4306 15733 4338
rect 15767 4306 15819 4338
rect 15853 4306 15905 4338
rect 15939 4306 15991 4338
rect 11482 4275 11506 4295
rect 11482 4241 11500 4275
rect 11540 4261 11564 4295
rect 11534 4241 11564 4261
rect 11482 4226 11564 4241
rect 11482 4202 11506 4226
rect 11482 4168 11500 4202
rect 11540 4192 11564 4226
rect 14740 4272 14774 4306
rect 14808 4272 14844 4306
rect 14878 4272 14914 4306
rect 14948 4272 14984 4306
rect 15018 4272 15054 4306
rect 15088 4272 15124 4306
rect 15158 4272 15194 4306
rect 15228 4272 15264 4306
rect 15298 4272 15334 4306
rect 15368 4272 15404 4306
rect 15438 4272 15474 4306
rect 15508 4272 15544 4306
rect 15578 4272 15614 4306
rect 15648 4272 15684 4306
rect 15718 4304 15733 4306
rect 15788 4304 15819 4306
rect 15718 4272 15754 4304
rect 15788 4272 15824 4304
rect 15858 4272 15894 4306
rect 15939 4304 15964 4306
rect 16025 4304 16033 4338
rect 15928 4272 15964 4304
rect 15998 4272 16033 4304
rect 14740 4266 16033 4272
rect 14740 4246 15733 4266
rect 14740 4238 15554 4246
rect 15588 4238 15626 4246
rect 15660 4238 15733 4246
rect 15767 4238 15819 4266
rect 15853 4238 15905 4266
rect 15939 4238 15991 4266
rect 11626 4194 11728 4210
rect 14528 4194 14630 4210
rect 14740 4204 14774 4238
rect 14808 4204 14844 4238
rect 14878 4204 14914 4238
rect 14948 4204 14984 4238
rect 15018 4204 15054 4238
rect 15088 4204 15124 4238
rect 15158 4204 15194 4238
rect 15228 4204 15264 4238
rect 15298 4204 15334 4238
rect 15368 4204 15404 4238
rect 15438 4204 15474 4238
rect 15508 4204 15544 4238
rect 15588 4212 15614 4238
rect 15660 4212 15684 4238
rect 15578 4204 15614 4212
rect 15648 4204 15684 4212
rect 15718 4232 15733 4238
rect 15788 4232 15819 4238
rect 15718 4204 15754 4232
rect 15788 4204 15824 4232
rect 15858 4204 15894 4238
rect 15939 4232 15964 4238
rect 16025 4232 16033 4266
rect 15928 4204 15964 4232
rect 15998 4204 16033 4232
rect 14740 4194 16033 4204
rect 11534 4168 11564 4192
rect 11482 4157 11564 4168
rect 11660 4160 11694 4194
rect 14562 4160 14596 4194
rect 14740 4173 15733 4194
rect 14740 4170 15484 4173
rect 15518 4170 15560 4173
rect 15594 4170 15636 4173
rect 15670 4170 15733 4173
rect 15767 4170 15819 4194
rect 15853 4170 15905 4194
rect 15939 4170 15991 4194
rect 11482 4129 11506 4157
rect 11482 4095 11500 4129
rect 11540 4123 11564 4157
rect 11626 4144 11728 4160
rect 14528 4144 14630 4160
rect 11534 4095 11564 4123
rect 11482 4088 11564 4095
rect 11482 4056 11506 4088
rect 11482 4022 11500 4056
rect 11540 4054 11564 4088
rect 11534 4051 11564 4054
rect 14740 4136 14774 4170
rect 14808 4136 14844 4170
rect 14878 4136 14914 4170
rect 14948 4136 14984 4170
rect 15018 4136 15054 4170
rect 15088 4136 15124 4170
rect 15158 4136 15194 4170
rect 15228 4136 15264 4170
rect 15298 4136 15334 4170
rect 15368 4136 15404 4170
rect 15438 4136 15474 4170
rect 15518 4139 15544 4170
rect 15594 4139 15614 4170
rect 15670 4139 15684 4170
rect 15508 4136 15544 4139
rect 15578 4136 15614 4139
rect 15648 4136 15684 4139
rect 15718 4160 15733 4170
rect 15788 4160 15819 4170
rect 15718 4136 15754 4160
rect 15788 4136 15824 4160
rect 15858 4136 15894 4170
rect 15939 4160 15964 4170
rect 16025 4160 16033 4194
rect 15928 4136 15964 4160
rect 15998 4136 16033 4160
rect 14740 4122 16033 4136
rect 14740 4102 15733 4122
rect 15767 4102 15819 4122
rect 15853 4102 15905 4122
rect 15939 4102 15991 4122
rect 14740 4068 14774 4102
rect 14808 4068 14844 4102
rect 14878 4068 14914 4102
rect 14948 4068 14984 4102
rect 15018 4068 15054 4102
rect 15088 4068 15124 4102
rect 15158 4068 15194 4102
rect 15228 4068 15264 4102
rect 15298 4068 15334 4102
rect 15368 4068 15404 4102
rect 15438 4088 15474 4102
rect 15508 4092 15544 4102
rect 15578 4092 15614 4102
rect 15648 4092 15684 4102
rect 15439 4068 15474 4088
rect 15518 4068 15544 4092
rect 15594 4068 15614 4092
rect 15670 4068 15684 4092
rect 15718 4088 15733 4102
rect 15788 4088 15819 4102
rect 15718 4068 15754 4088
rect 15788 4068 15824 4088
rect 15858 4068 15894 4102
rect 15939 4088 15964 4102
rect 16025 4088 16033 4122
rect 15928 4068 15964 4088
rect 15998 4068 16033 4088
rect 14740 4054 15405 4068
rect 15439 4058 15484 4068
rect 15518 4058 15560 4068
rect 15594 4058 15636 4068
rect 15670 4058 16033 4068
rect 15439 4054 16033 4058
rect 14740 4051 16033 4054
rect 11534 4022 11583 4051
rect 11482 4019 11583 4022
rect 11482 3985 11506 4019
rect 11540 4017 11583 4019
rect 11622 4017 11656 4051
rect 11691 4017 11726 4051
rect 11763 4017 11795 4051
rect 11835 4017 11864 4051
rect 11907 4017 11933 4051
rect 11979 4017 12002 4051
rect 12051 4017 12071 4051
rect 12123 4017 12140 4051
rect 12195 4017 12209 4051
rect 12267 4017 12278 4051
rect 12339 4017 12347 4051
rect 12411 4017 12416 4051
rect 12483 4017 12485 4051
rect 12519 4017 12521 4051
rect 12588 4017 12593 4051
rect 12657 4017 12665 4051
rect 12726 4017 12737 4051
rect 12795 4017 12809 4051
rect 12864 4017 12881 4051
rect 12933 4017 12953 4051
rect 13002 4017 13025 4051
rect 13071 4017 13097 4051
rect 13140 4017 13169 4051
rect 13209 4017 13241 4051
rect 13278 4017 13313 4051
rect 13347 4017 13382 4051
rect 13419 4017 13451 4051
rect 13491 4017 13520 4051
rect 13563 4017 13589 4051
rect 13635 4017 13658 4051
rect 13707 4017 13727 4051
rect 13779 4017 13796 4051
rect 13851 4017 13865 4051
rect 13923 4017 13934 4051
rect 13995 4017 14002 4051
rect 14067 4017 14070 4051
rect 14104 4017 14105 4051
rect 14172 4017 14177 4051
rect 14240 4017 14249 4051
rect 14308 4017 14321 4051
rect 14376 4017 14393 4051
rect 14444 4017 14465 4051
rect 14512 4017 14537 4051
rect 14580 4017 14609 4051
rect 14648 4017 14681 4051
rect 14716 4017 14753 4051
rect 14787 4034 14825 4051
rect 14859 4034 14897 4051
rect 14931 4034 14969 4051
rect 15003 4034 15041 4051
rect 15075 4034 15113 4051
rect 15147 4034 15185 4051
rect 15219 4034 15257 4051
rect 15291 4034 15329 4051
rect 15363 4050 16033 4051
rect 15363 4034 15733 4050
rect 15767 4034 15819 4050
rect 15853 4034 15905 4050
rect 15939 4034 15991 4050
rect 14808 4017 14825 4034
rect 14878 4017 14897 4034
rect 14948 4017 14969 4034
rect 15018 4017 15041 4034
rect 15088 4017 15113 4034
rect 15158 4017 15185 4034
rect 15228 4017 15257 4034
rect 15298 4017 15329 4034
rect 11540 3985 11564 4017
rect 11482 3950 11564 3985
rect 344 3909 10962 3925
rect 344 3907 470 3909
rect 504 3907 538 3909
rect 572 3907 606 3909
rect 640 3907 674 3909
rect 344 3906 379 3907
rect 344 3872 360 3906
rect 413 3873 452 3907
rect 504 3875 525 3907
rect 572 3875 598 3907
rect 640 3875 671 3907
rect 708 3875 742 3909
rect 776 3907 810 3909
rect 844 3907 878 3909
rect 912 3907 946 3909
rect 980 3907 1014 3909
rect 1048 3907 1082 3909
rect 1116 3907 1150 3909
rect 1184 3907 1218 3909
rect 778 3875 810 3907
rect 851 3875 878 3907
rect 924 3875 946 3907
rect 997 3875 1014 3907
rect 1070 3875 1082 3907
rect 1143 3875 1150 3907
rect 1216 3875 1218 3907
rect 1252 3907 1286 3909
rect 1320 3907 1354 3909
rect 1388 3907 1422 3909
rect 1456 3907 1490 3909
rect 1524 3907 1558 3909
rect 1592 3907 1626 3909
rect 1660 3907 1694 3909
rect 1252 3875 1255 3907
rect 1320 3875 1328 3907
rect 1388 3875 1401 3907
rect 1456 3875 1474 3907
rect 1524 3875 1547 3907
rect 1592 3875 1620 3907
rect 1660 3875 1693 3907
rect 1728 3875 1762 3909
rect 1796 3907 1830 3909
rect 1864 3907 1898 3909
rect 1932 3907 1966 3909
rect 2000 3907 2034 3909
rect 2068 3907 2102 3909
rect 2136 3907 2170 3909
rect 1800 3875 1830 3907
rect 1873 3875 1898 3907
rect 1946 3875 1966 3907
rect 2019 3875 2034 3907
rect 2092 3875 2102 3907
rect 2165 3875 2170 3907
rect 2204 3907 2238 3909
rect 486 3873 525 3875
rect 559 3873 598 3875
rect 632 3873 671 3875
rect 705 3873 744 3875
rect 778 3873 817 3875
rect 851 3873 890 3875
rect 924 3873 963 3875
rect 997 3873 1036 3875
rect 1070 3873 1109 3875
rect 1143 3873 1182 3875
rect 1216 3873 1255 3875
rect 1289 3873 1328 3875
rect 1362 3873 1401 3875
rect 1435 3873 1474 3875
rect 1508 3873 1547 3875
rect 1581 3873 1620 3875
rect 1654 3873 1693 3875
rect 1727 3873 1766 3875
rect 1800 3873 1839 3875
rect 1873 3873 1912 3875
rect 1946 3873 1985 3875
rect 2019 3873 2058 3875
rect 2092 3873 2131 3875
rect 2165 3873 2204 3875
rect 2272 3907 2306 3909
rect 2340 3907 2374 3909
rect 2408 3907 2442 3909
rect 2476 3907 2510 3909
rect 2544 3907 2578 3909
rect 2612 3907 2646 3909
rect 2272 3875 2277 3907
rect 2340 3875 2350 3907
rect 2408 3875 2423 3907
rect 2476 3875 2496 3907
rect 2544 3875 2569 3907
rect 2612 3875 2642 3907
rect 2680 3875 2714 3909
rect 2748 3907 2782 3909
rect 2816 3907 2850 3909
rect 2884 3907 2918 3909
rect 2952 3907 2986 3909
rect 3020 3907 3054 3909
rect 3088 3907 3122 3909
rect 3156 3907 3190 3909
rect 2749 3875 2782 3907
rect 2822 3875 2850 3907
rect 2895 3875 2918 3907
rect 2968 3875 2986 3907
rect 3041 3875 3054 3907
rect 3114 3875 3122 3907
rect 3187 3875 3190 3907
rect 3224 3907 3258 3909
rect 3292 3907 3326 3909
rect 3360 3907 3394 3909
rect 3428 3907 3462 3909
rect 3496 3907 3530 3909
rect 3564 3907 3598 3909
rect 3632 3907 3666 3909
rect 3700 3907 3734 3909
rect 3224 3875 3226 3907
rect 3292 3875 3299 3907
rect 3360 3875 3372 3907
rect 3428 3875 3444 3907
rect 3496 3875 3516 3907
rect 3564 3875 3588 3907
rect 3632 3875 3660 3907
rect 3700 3875 3732 3907
rect 3768 3875 3802 3909
rect 3836 3907 3870 3909
rect 3904 3907 3938 3909
rect 3972 3907 4006 3909
rect 4040 3907 4074 3909
rect 4108 3907 4142 3909
rect 4176 3907 4210 3909
rect 4244 3907 4278 3909
rect 4312 3907 4346 3909
rect 3838 3875 3870 3907
rect 3910 3875 3938 3907
rect 3982 3875 4006 3907
rect 4054 3875 4074 3907
rect 4126 3875 4142 3907
rect 4198 3875 4210 3907
rect 4270 3875 4278 3907
rect 4342 3875 4346 3907
rect 4380 3907 4414 3909
rect 2238 3873 2277 3875
rect 2311 3873 2350 3875
rect 2384 3873 2423 3875
rect 2457 3873 2496 3875
rect 2530 3873 2569 3875
rect 2603 3873 2642 3875
rect 2676 3873 2715 3875
rect 2749 3873 2788 3875
rect 2822 3873 2861 3875
rect 2895 3873 2934 3875
rect 2968 3873 3007 3875
rect 3041 3873 3080 3875
rect 3114 3873 3153 3875
rect 3187 3873 3226 3875
rect 3260 3873 3299 3875
rect 3333 3873 3372 3875
rect 3406 3873 3444 3875
rect 3478 3873 3516 3875
rect 3550 3873 3588 3875
rect 3622 3873 3660 3875
rect 3694 3873 3732 3875
rect 3766 3873 3804 3875
rect 3838 3873 3876 3875
rect 3910 3873 3948 3875
rect 3982 3873 4020 3875
rect 4054 3873 4092 3875
rect 4126 3873 4164 3875
rect 4198 3873 4236 3875
rect 4270 3873 4308 3875
rect 4342 3873 4380 3875
rect 4448 3907 4482 3909
rect 4516 3907 4550 3909
rect 4584 3907 4618 3909
rect 4652 3907 4686 3909
rect 4720 3907 4754 3909
rect 4788 3907 4822 3909
rect 4856 3907 4890 3909
rect 4924 3907 4958 3909
rect 4448 3875 4452 3907
rect 4516 3875 4524 3907
rect 4584 3875 4596 3907
rect 4652 3875 4668 3907
rect 4720 3875 4740 3907
rect 4788 3875 4812 3907
rect 4856 3875 4884 3907
rect 4924 3875 4956 3907
rect 4992 3875 5026 3909
rect 5060 3907 5094 3909
rect 5128 3907 5162 3909
rect 5196 3907 5230 3909
rect 5264 3907 5298 3909
rect 5332 3907 5366 3909
rect 5400 3907 5434 3909
rect 5468 3907 5502 3909
rect 5536 3907 5570 3909
rect 5062 3875 5094 3907
rect 5134 3875 5162 3907
rect 5206 3875 5230 3907
rect 5278 3875 5298 3907
rect 5350 3875 5366 3907
rect 5422 3875 5434 3907
rect 5494 3875 5502 3907
rect 5566 3875 5570 3907
rect 5604 3907 5638 3909
rect 4414 3873 4452 3875
rect 4486 3873 4524 3875
rect 4558 3873 4596 3875
rect 4630 3873 4668 3875
rect 4702 3873 4740 3875
rect 4774 3873 4812 3875
rect 4846 3873 4884 3875
rect 4918 3873 4956 3875
rect 4990 3873 5028 3875
rect 5062 3873 5100 3875
rect 5134 3873 5172 3875
rect 5206 3873 5244 3875
rect 5278 3873 5316 3875
rect 5350 3873 5388 3875
rect 5422 3873 5460 3875
rect 5494 3873 5532 3875
rect 5566 3873 5604 3875
rect 5672 3907 5706 3909
rect 5740 3907 5774 3909
rect 5808 3907 5842 3909
rect 5876 3907 5910 3909
rect 5944 3907 5978 3909
rect 6012 3907 6046 3909
rect 6080 3907 6114 3909
rect 6148 3907 6182 3909
rect 5672 3875 5676 3907
rect 5740 3875 5748 3907
rect 5808 3875 5820 3907
rect 5876 3875 5892 3907
rect 5944 3875 5964 3907
rect 6012 3875 6036 3907
rect 6080 3875 6108 3907
rect 6148 3875 6180 3907
rect 6216 3875 6250 3909
rect 6284 3907 6318 3909
rect 6352 3907 6386 3909
rect 6420 3907 6454 3909
rect 6488 3907 6522 3909
rect 6556 3907 6590 3909
rect 6624 3907 6658 3909
rect 6692 3907 6726 3909
rect 6760 3907 6794 3909
rect 6286 3875 6318 3907
rect 6358 3875 6386 3907
rect 6430 3875 6454 3907
rect 6502 3875 6522 3907
rect 6574 3875 6590 3907
rect 6646 3875 6658 3907
rect 6718 3875 6726 3907
rect 6790 3875 6794 3907
rect 6828 3907 6862 3909
rect 5638 3873 5676 3875
rect 5710 3873 5748 3875
rect 5782 3873 5820 3875
rect 5854 3873 5892 3875
rect 5926 3873 5964 3875
rect 5998 3873 6036 3875
rect 6070 3873 6108 3875
rect 6142 3873 6180 3875
rect 6214 3873 6252 3875
rect 6286 3873 6324 3875
rect 6358 3873 6396 3875
rect 6430 3873 6468 3875
rect 6502 3873 6540 3875
rect 6574 3873 6612 3875
rect 6646 3873 6684 3875
rect 6718 3873 6756 3875
rect 6790 3873 6828 3875
rect 6896 3907 6930 3909
rect 6964 3907 6998 3909
rect 7032 3907 7066 3909
rect 7100 3907 7134 3909
rect 7168 3907 7202 3909
rect 7236 3907 7270 3909
rect 7304 3907 7338 3909
rect 7372 3907 7406 3909
rect 6896 3875 6900 3907
rect 6964 3875 6972 3907
rect 7032 3875 7044 3907
rect 7100 3875 7116 3907
rect 7168 3875 7188 3907
rect 7236 3875 7260 3907
rect 7304 3875 7332 3907
rect 7372 3875 7404 3907
rect 7440 3875 7474 3909
rect 7508 3907 7542 3909
rect 7576 3907 7610 3909
rect 7644 3907 7678 3909
rect 7712 3907 7746 3909
rect 7780 3907 7814 3909
rect 7848 3907 7882 3909
rect 7916 3907 7950 3909
rect 7984 3907 8018 3909
rect 7510 3875 7542 3907
rect 7582 3875 7610 3907
rect 7654 3875 7678 3907
rect 7726 3875 7746 3907
rect 7798 3875 7814 3907
rect 7870 3875 7882 3907
rect 7942 3875 7950 3907
rect 8014 3875 8018 3907
rect 8052 3907 8086 3909
rect 6862 3873 6900 3875
rect 6934 3873 6972 3875
rect 7006 3873 7044 3875
rect 7078 3873 7116 3875
rect 7150 3873 7188 3875
rect 7222 3873 7260 3875
rect 7294 3873 7332 3875
rect 7366 3873 7404 3875
rect 7438 3873 7476 3875
rect 7510 3873 7548 3875
rect 7582 3873 7620 3875
rect 7654 3873 7692 3875
rect 7726 3873 7764 3875
rect 7798 3873 7836 3875
rect 7870 3873 7908 3875
rect 7942 3873 7980 3875
rect 8014 3873 8052 3875
rect 8120 3907 8154 3909
rect 8188 3907 8222 3909
rect 8256 3907 8290 3909
rect 8324 3907 8359 3909
rect 8393 3907 8428 3909
rect 8462 3907 8497 3909
rect 8531 3907 8566 3909
rect 8600 3907 8635 3909
rect 8669 3907 8704 3909
rect 8738 3907 8773 3909
rect 8120 3875 8124 3907
rect 8188 3875 8196 3907
rect 8256 3875 8268 3907
rect 8324 3875 8340 3907
rect 8393 3875 8412 3907
rect 8462 3875 8484 3907
rect 8531 3875 8556 3907
rect 8600 3875 8628 3907
rect 8669 3875 8700 3907
rect 8738 3875 8772 3907
rect 8807 3875 8842 3909
rect 8876 3907 8911 3909
rect 8945 3907 8980 3909
rect 9014 3907 9049 3909
rect 9083 3907 9118 3909
rect 9152 3907 9187 3909
rect 9221 3907 9256 3909
rect 9290 3907 9325 3909
rect 9359 3907 9394 3909
rect 9428 3907 9463 3909
rect 9497 3907 9532 3909
rect 9566 3907 9601 3909
rect 8878 3875 8911 3907
rect 8950 3875 8980 3907
rect 9022 3875 9049 3907
rect 9094 3875 9118 3907
rect 9166 3875 9187 3907
rect 9238 3875 9256 3907
rect 9310 3875 9325 3907
rect 9382 3875 9394 3907
rect 9454 3875 9463 3907
rect 9526 3875 9532 3907
rect 9598 3875 9601 3907
rect 9635 3907 9670 3909
rect 9635 3875 9636 3907
rect 8086 3873 8124 3875
rect 8158 3873 8196 3875
rect 8230 3873 8268 3875
rect 8302 3873 8340 3875
rect 8374 3873 8412 3875
rect 8446 3873 8484 3875
rect 8518 3873 8556 3875
rect 8590 3873 8628 3875
rect 8662 3873 8700 3875
rect 8734 3873 8772 3875
rect 8806 3873 8844 3875
rect 8878 3873 8916 3875
rect 8950 3873 8988 3875
rect 9022 3873 9060 3875
rect 9094 3873 9132 3875
rect 9166 3873 9204 3875
rect 9238 3873 9276 3875
rect 9310 3873 9348 3875
rect 9382 3873 9420 3875
rect 9454 3873 9492 3875
rect 9526 3873 9564 3875
rect 9598 3873 9636 3875
rect 9704 3907 9739 3909
rect 9773 3907 9808 3909
rect 9842 3907 9877 3909
rect 9911 3907 9946 3909
rect 9980 3907 10015 3909
rect 10049 3907 10084 3909
rect 10118 3907 10153 3909
rect 10187 3907 10222 3909
rect 10256 3907 10291 3909
rect 10325 3907 10360 3909
rect 10394 3907 10429 3909
rect 9704 3875 9708 3907
rect 9773 3875 9780 3907
rect 9842 3875 9852 3907
rect 9911 3875 9924 3907
rect 9980 3875 9996 3907
rect 10049 3875 10068 3907
rect 10118 3875 10140 3907
rect 10187 3875 10212 3907
rect 10256 3875 10284 3907
rect 10325 3875 10356 3907
rect 10394 3875 10428 3907
rect 10463 3875 10498 3909
rect 10532 3907 10567 3909
rect 10601 3907 10636 3909
rect 10670 3907 10705 3909
rect 10739 3907 10774 3909
rect 10808 3907 10843 3909
rect 10877 3907 10912 3909
rect 10534 3875 10567 3907
rect 10606 3875 10636 3907
rect 10678 3875 10705 3907
rect 10750 3875 10774 3907
rect 10822 3875 10843 3907
rect 10894 3875 10912 3907
rect 10946 3875 10962 3909
rect 9670 3873 9708 3875
rect 9742 3873 9780 3875
rect 9814 3873 9852 3875
rect 9886 3873 9924 3875
rect 9958 3873 9996 3875
rect 10030 3873 10068 3875
rect 10102 3873 10140 3875
rect 10174 3873 10212 3875
rect 10246 3873 10284 3875
rect 10318 3873 10356 3875
rect 10390 3873 10428 3875
rect 10462 3873 10500 3875
rect 10534 3873 10572 3875
rect 10606 3873 10644 3875
rect 10678 3873 10716 3875
rect 10750 3873 10788 3875
rect 10822 3873 10860 3875
rect 10894 3873 10962 3875
rect 394 3872 10962 3873
rect 344 3859 10962 3872
rect 344 3835 410 3859
rect 344 3801 360 3835
rect 394 3801 410 3835
rect 10896 3839 10962 3859
rect 10896 3805 10912 3839
rect 10946 3805 10962 3839
rect 344 3790 410 3801
rect 344 3730 360 3790
rect 394 3730 410 3790
rect 586 3769 588 3803
rect 622 3769 632 3803
rect 690 3769 711 3803
rect 758 3769 790 3803
rect 826 3769 860 3803
rect 903 3769 928 3803
rect 982 3769 996 3803
rect 1061 3769 1064 3803
rect 1098 3769 1106 3803
rect 1166 3769 1185 3803
rect 1234 3769 1264 3803
rect 1302 3769 1318 3803
rect 1442 3769 1444 3803
rect 1478 3769 1488 3803
rect 1546 3769 1567 3803
rect 1614 3769 1646 3803
rect 1682 3769 1716 3803
rect 1759 3769 1784 3803
rect 1838 3769 1852 3803
rect 1917 3769 1920 3803
rect 1954 3769 1962 3803
rect 2022 3769 2041 3803
rect 2090 3769 2120 3803
rect 2158 3769 2174 3803
rect 2298 3769 2300 3803
rect 2334 3769 2344 3803
rect 2402 3769 2423 3803
rect 2470 3769 2502 3803
rect 2538 3769 2572 3803
rect 2615 3769 2640 3803
rect 2694 3769 2708 3803
rect 2773 3769 2776 3803
rect 2810 3769 2818 3803
rect 2878 3769 2897 3803
rect 2946 3769 2976 3803
rect 3014 3769 3030 3803
rect 3154 3769 3156 3803
rect 3190 3769 3200 3803
rect 3258 3769 3279 3803
rect 3326 3769 3358 3803
rect 3394 3769 3428 3803
rect 3471 3769 3496 3803
rect 3550 3769 3564 3803
rect 3629 3769 3632 3803
rect 3666 3769 3674 3803
rect 3734 3769 3753 3803
rect 3802 3769 3832 3803
rect 3870 3769 3886 3803
rect 4010 3769 4012 3803
rect 4046 3769 4056 3803
rect 4114 3769 4135 3803
rect 4182 3769 4214 3803
rect 4250 3769 4284 3803
rect 4327 3769 4352 3803
rect 4406 3769 4420 3803
rect 4485 3769 4488 3803
rect 4522 3769 4530 3803
rect 4590 3769 4609 3803
rect 4658 3769 4688 3803
rect 4726 3769 4742 3803
rect 4866 3769 4868 3803
rect 4902 3769 4912 3803
rect 4970 3769 4991 3803
rect 5038 3769 5070 3803
rect 5106 3769 5140 3803
rect 5183 3769 5208 3803
rect 5262 3769 5276 3803
rect 5341 3769 5344 3803
rect 5378 3769 5386 3803
rect 5446 3769 5465 3803
rect 5514 3769 5544 3803
rect 5582 3769 5598 3803
rect 5722 3769 5724 3803
rect 5758 3769 5768 3803
rect 5826 3769 5847 3803
rect 5894 3769 5926 3803
rect 5962 3769 5996 3803
rect 6039 3769 6064 3803
rect 6118 3769 6132 3803
rect 6197 3769 6200 3803
rect 6234 3769 6242 3803
rect 6302 3769 6321 3803
rect 6370 3769 6400 3803
rect 6438 3769 6454 3803
rect 6578 3769 6580 3803
rect 6614 3769 6624 3803
rect 6682 3769 6703 3803
rect 6750 3769 6782 3803
rect 6818 3769 6852 3803
rect 6895 3769 6920 3803
rect 6974 3769 6988 3803
rect 7053 3769 7056 3803
rect 7090 3769 7098 3803
rect 7158 3769 7177 3803
rect 7226 3769 7256 3803
rect 7294 3769 7310 3803
rect 7434 3769 7436 3803
rect 7470 3769 7480 3803
rect 7538 3769 7559 3803
rect 7606 3769 7638 3803
rect 7674 3769 7708 3803
rect 7751 3769 7776 3803
rect 7830 3769 7844 3803
rect 7909 3769 7912 3803
rect 7946 3769 7954 3803
rect 8014 3769 8033 3803
rect 8082 3769 8112 3803
rect 8150 3769 8166 3803
rect 8290 3769 8292 3803
rect 8326 3769 8336 3803
rect 8394 3769 8415 3803
rect 8462 3769 8494 3803
rect 8530 3769 8564 3803
rect 8607 3769 8632 3803
rect 8686 3769 8700 3803
rect 8765 3769 8768 3803
rect 8802 3769 8810 3803
rect 8870 3769 8889 3803
rect 8938 3769 8968 3803
rect 9006 3769 9022 3803
rect 9146 3769 9148 3803
rect 9182 3769 9192 3803
rect 9250 3769 9271 3803
rect 9318 3769 9350 3803
rect 9386 3769 9420 3803
rect 9463 3769 9488 3803
rect 9542 3769 9556 3803
rect 9621 3769 9624 3803
rect 9658 3769 9666 3803
rect 9726 3769 9745 3803
rect 9794 3769 9824 3803
rect 9862 3769 9878 3803
rect 10002 3769 10004 3803
rect 10038 3769 10048 3803
rect 10106 3769 10127 3803
rect 10174 3769 10206 3803
rect 10242 3769 10276 3803
rect 10319 3769 10344 3803
rect 10398 3769 10412 3803
rect 10477 3769 10480 3803
rect 10514 3769 10522 3803
rect 10582 3769 10601 3803
rect 10650 3769 10680 3803
rect 10718 3769 10734 3803
rect 10896 3790 10962 3805
rect 344 3718 410 3730
rect 344 3659 360 3718
rect 394 3659 410 3718
rect 10896 3735 10912 3790
rect 10946 3735 10962 3790
rect 10896 3718 10962 3735
rect 344 3646 410 3659
rect 344 3589 360 3646
rect 394 3589 410 3646
rect 344 3574 410 3589
rect 344 3519 360 3574
rect 394 3519 410 3574
rect 344 3502 410 3519
rect 344 3449 360 3502
rect 394 3449 410 3502
rect 344 3430 410 3449
rect 344 3379 360 3430
rect 394 3379 410 3430
rect 344 3358 410 3379
rect 344 3309 360 3358
rect 394 3309 410 3358
rect 344 3286 410 3309
rect 344 3239 360 3286
rect 394 3239 410 3286
rect 344 3214 410 3239
rect 344 3169 360 3214
rect 394 3169 410 3214
rect 344 3142 410 3169
rect 344 3099 360 3142
rect 394 3099 410 3142
rect 344 3070 410 3099
rect 344 3029 360 3070
rect 394 3029 410 3070
rect 344 2998 410 3029
rect 344 2959 360 2998
rect 394 2959 410 2998
rect 344 2926 410 2959
rect 344 2889 360 2926
rect 394 2889 410 2926
rect 344 2854 410 2889
rect 344 2819 360 2854
rect 394 2819 410 2854
rect 344 2783 410 2819
rect 344 2748 360 2783
rect 394 2748 410 2783
rect 344 2713 410 2748
rect 344 2676 360 2713
rect 394 2676 410 2713
rect 344 2643 410 2676
rect 344 2604 360 2643
rect 394 2604 410 2643
rect 344 2573 410 2604
rect 344 2532 360 2573
rect 394 2532 410 2573
rect 344 2503 410 2532
rect 344 2460 360 2503
rect 394 2460 410 2503
rect 344 2433 410 2460
rect 344 2388 360 2433
rect 394 2388 410 2433
rect 344 2363 410 2388
rect 344 2316 360 2363
rect 394 2316 410 2363
rect 500 3659 534 3675
rect 500 3591 534 3612
rect 500 3523 534 3540
rect 500 3455 534 3468
rect 500 3387 534 3396
rect 500 3319 534 3324
rect 500 3251 534 3252
rect 500 3214 534 3217
rect 500 3142 534 3149
rect 500 3070 534 3081
rect 500 2998 534 3013
rect 500 2926 534 2945
rect 500 2854 534 2877
rect 500 2782 534 2809
rect 500 2707 534 2741
rect 500 2639 534 2673
rect 500 2571 534 2605
rect 500 2503 534 2537
rect 500 2435 534 2469
rect 500 2367 534 2401
rect 500 2317 534 2333
rect 1356 3664 1390 3675
rect 1356 3592 1390 3625
rect 1356 3523 1390 3557
rect 1356 3455 1390 3486
rect 1356 3387 1390 3414
rect 1356 3319 1390 3342
rect 1356 3251 1390 3270
rect 1356 3183 1390 3198
rect 1356 3115 1390 3126
rect 1356 3047 1390 3054
rect 1356 2979 1390 2982
rect 1356 2944 1390 2945
rect 1356 2872 1390 2877
rect 1356 2800 1390 2809
rect 1356 2728 1390 2741
rect 1356 2656 1390 2673
rect 1356 2584 1390 2605
rect 1356 2512 1390 2537
rect 1356 2440 1390 2469
rect 1356 2368 1390 2401
rect 1356 2317 1390 2333
rect 2212 3664 2246 3675
rect 2212 3592 2246 3625
rect 2212 3523 2246 3557
rect 2212 3455 2246 3486
rect 2212 3387 2246 3414
rect 2212 3319 2246 3342
rect 2212 3251 2246 3270
rect 2212 3183 2246 3198
rect 2212 3115 2246 3126
rect 2212 3047 2246 3054
rect 2212 2979 2246 2982
rect 2212 2944 2246 2945
rect 2212 2872 2246 2877
rect 2212 2800 2246 2809
rect 2212 2728 2246 2741
rect 2212 2656 2246 2673
rect 2212 2584 2246 2605
rect 2212 2512 2246 2537
rect 2212 2440 2246 2469
rect 2212 2368 2246 2401
rect 2212 2317 2246 2333
rect 3068 3664 3102 3675
rect 3068 3592 3102 3625
rect 3068 3523 3102 3557
rect 3068 3455 3102 3486
rect 3068 3387 3102 3414
rect 3068 3319 3102 3342
rect 3068 3251 3102 3270
rect 3068 3183 3102 3198
rect 3068 3115 3102 3126
rect 3068 3047 3102 3054
rect 3068 2979 3102 2982
rect 3068 2944 3102 2945
rect 3068 2872 3102 2877
rect 3068 2800 3102 2809
rect 3068 2728 3102 2741
rect 3068 2656 3102 2673
rect 3068 2584 3102 2605
rect 3068 2512 3102 2537
rect 3068 2440 3102 2469
rect 3068 2368 3102 2401
rect 3068 2317 3102 2333
rect 3924 3664 3958 3675
rect 3924 3592 3958 3625
rect 3924 3523 3958 3557
rect 3924 3455 3958 3486
rect 3924 3387 3958 3414
rect 3924 3319 3958 3342
rect 3924 3251 3958 3270
rect 3924 3183 3958 3198
rect 3924 3115 3958 3126
rect 3924 3047 3958 3054
rect 3924 2979 3958 2982
rect 3924 2944 3958 2945
rect 3924 2872 3958 2877
rect 3924 2800 3958 2809
rect 3924 2728 3958 2741
rect 3924 2656 3958 2673
rect 3924 2584 3958 2605
rect 3924 2512 3958 2537
rect 3924 2440 3958 2469
rect 3924 2368 3958 2401
rect 3924 2317 3958 2333
rect 4780 3664 4814 3675
rect 4780 3592 4814 3625
rect 4780 3523 4814 3557
rect 4780 3455 4814 3486
rect 4780 3387 4814 3414
rect 4780 3319 4814 3342
rect 4780 3251 4814 3270
rect 4780 3183 4814 3198
rect 4780 3115 4814 3126
rect 4780 3047 4814 3054
rect 4780 2979 4814 2982
rect 4780 2944 4814 2945
rect 4780 2872 4814 2877
rect 4780 2800 4814 2809
rect 4780 2728 4814 2741
rect 4780 2656 4814 2673
rect 4780 2584 4814 2605
rect 4780 2512 4814 2537
rect 4780 2440 4814 2469
rect 4780 2368 4814 2401
rect 4780 2317 4814 2333
rect 5636 3664 5670 3675
rect 5636 3592 5670 3625
rect 5636 3523 5670 3557
rect 5636 3455 5670 3486
rect 5636 3387 5670 3414
rect 5636 3319 5670 3342
rect 5636 3251 5670 3270
rect 5636 3183 5670 3198
rect 5636 3115 5670 3126
rect 5636 3047 5670 3054
rect 5636 2979 5670 2982
rect 5636 2944 5670 2945
rect 5636 2872 5670 2877
rect 5636 2800 5670 2809
rect 5636 2728 5670 2741
rect 5636 2656 5670 2673
rect 5636 2584 5670 2605
rect 5636 2512 5670 2537
rect 5636 2440 5670 2469
rect 5636 2368 5670 2401
rect 5636 2317 5670 2333
rect 6492 3664 6526 3675
rect 6492 3592 6526 3625
rect 6492 3523 6526 3557
rect 6492 3455 6526 3486
rect 6492 3387 6526 3414
rect 6492 3319 6526 3342
rect 6492 3251 6526 3270
rect 6492 3183 6526 3198
rect 6492 3115 6526 3126
rect 6492 3047 6526 3054
rect 6492 2979 6526 2982
rect 6492 2944 6526 2945
rect 6492 2872 6526 2877
rect 6492 2800 6526 2809
rect 6492 2728 6526 2741
rect 6492 2656 6526 2673
rect 6492 2584 6526 2605
rect 6492 2512 6526 2537
rect 6492 2440 6526 2469
rect 6492 2368 6526 2401
rect 6492 2317 6526 2333
rect 7348 3664 7382 3675
rect 7348 3592 7382 3625
rect 7348 3523 7382 3557
rect 7348 3455 7382 3486
rect 7348 3387 7382 3414
rect 7348 3319 7382 3342
rect 7348 3251 7382 3270
rect 7348 3183 7382 3198
rect 7348 3115 7382 3126
rect 7348 3047 7382 3054
rect 7348 2979 7382 2982
rect 7348 2944 7382 2945
rect 7348 2872 7382 2877
rect 7348 2800 7382 2809
rect 7348 2728 7382 2741
rect 7348 2656 7382 2673
rect 7348 2584 7382 2605
rect 7348 2512 7382 2537
rect 7348 2440 7382 2469
rect 7348 2368 7382 2401
rect 7348 2317 7382 2333
rect 8204 3664 8238 3675
rect 8204 3592 8238 3625
rect 8204 3523 8238 3557
rect 8204 3455 8238 3486
rect 8204 3387 8238 3414
rect 8204 3319 8238 3342
rect 8204 3251 8238 3270
rect 8204 3183 8238 3198
rect 8204 3115 8238 3126
rect 8204 3047 8238 3054
rect 8204 2979 8238 2982
rect 8204 2944 8238 2945
rect 8204 2872 8238 2877
rect 8204 2800 8238 2809
rect 8204 2728 8238 2741
rect 8204 2656 8238 2673
rect 8204 2584 8238 2605
rect 8204 2512 8238 2537
rect 8204 2440 8238 2469
rect 8204 2368 8238 2401
rect 8204 2317 8238 2333
rect 9060 3664 9094 3675
rect 9060 3592 9094 3625
rect 9060 3523 9094 3557
rect 9060 3455 9094 3486
rect 9060 3387 9094 3414
rect 9060 3319 9094 3342
rect 9060 3251 9094 3270
rect 9060 3183 9094 3198
rect 9060 3115 9094 3126
rect 9060 3047 9094 3054
rect 9060 2979 9094 2982
rect 9060 2944 9094 2945
rect 9060 2872 9094 2877
rect 9060 2800 9094 2809
rect 9060 2728 9094 2741
rect 9060 2656 9094 2673
rect 9060 2584 9094 2605
rect 9060 2512 9094 2537
rect 9060 2440 9094 2469
rect 9060 2368 9094 2401
rect 9060 2317 9094 2333
rect 9916 3664 9950 3675
rect 9916 3592 9950 3625
rect 9916 3523 9950 3557
rect 9916 3455 9950 3486
rect 9916 3387 9950 3414
rect 9916 3319 9950 3342
rect 9916 3251 9950 3270
rect 9916 3183 9950 3198
rect 9916 3115 9950 3126
rect 9916 3047 9950 3054
rect 9916 2979 9950 2982
rect 9916 2944 9950 2945
rect 9916 2872 9950 2877
rect 9916 2800 9950 2809
rect 9916 2728 9950 2741
rect 9916 2656 9950 2673
rect 9916 2584 9950 2605
rect 9916 2512 9950 2537
rect 9916 2440 9950 2469
rect 9916 2368 9950 2401
rect 9916 2317 9950 2333
rect 10772 3664 10806 3675
rect 10772 3592 10806 3625
rect 10772 3523 10806 3557
rect 10772 3455 10806 3486
rect 10772 3387 10806 3414
rect 10772 3319 10806 3342
rect 10772 3251 10806 3270
rect 10772 3183 10806 3198
rect 10772 3115 10806 3126
rect 10772 3047 10806 3054
rect 10772 2979 10806 2982
rect 10772 2944 10806 2945
rect 10772 2872 10806 2877
rect 10772 2800 10806 2809
rect 10772 2728 10806 2741
rect 10772 2656 10806 2673
rect 10772 2584 10806 2605
rect 10772 2512 10806 2537
rect 10772 2440 10806 2469
rect 10772 2368 10806 2401
rect 10772 2317 10806 2333
rect 10896 3665 10912 3718
rect 10946 3665 10962 3718
rect 10896 3646 10962 3665
rect 10896 3595 10912 3646
rect 10946 3595 10962 3646
rect 10896 3574 10962 3595
rect 10896 3525 10912 3574
rect 10946 3525 10962 3574
rect 10896 3502 10962 3525
rect 10896 3455 10912 3502
rect 10946 3455 10962 3502
rect 10896 3430 10962 3455
rect 10896 3385 10912 3430
rect 10946 3385 10962 3430
rect 10896 3358 10962 3385
rect 10896 3315 10912 3358
rect 10946 3315 10962 3358
rect 10896 3286 10962 3315
rect 10896 3245 10912 3286
rect 10946 3245 10962 3286
rect 10896 3214 10962 3245
rect 10896 3175 10912 3214
rect 10946 3175 10962 3214
rect 10896 3142 10962 3175
rect 10896 3105 10912 3142
rect 10946 3105 10962 3142
rect 10896 3070 10962 3105
rect 10896 3035 10912 3070
rect 10946 3035 10962 3070
rect 10896 2999 10962 3035
rect 10896 2964 10912 2999
rect 10946 2964 10962 2999
rect 10896 2929 10962 2964
rect 10896 2892 10912 2929
rect 10946 2892 10962 2929
rect 10896 2859 10962 2892
rect 10896 2820 10912 2859
rect 10946 2820 10962 2859
rect 10896 2789 10962 2820
rect 10896 2748 10912 2789
rect 10946 2748 10962 2789
rect 10896 2719 10962 2748
rect 10896 2676 10912 2719
rect 10946 2676 10962 2719
rect 10896 2649 10962 2676
rect 10896 2604 10912 2649
rect 10946 2604 10962 2649
rect 10896 2578 10962 2604
rect 10896 2532 10912 2578
rect 10946 2532 10962 2578
rect 10896 2507 10962 2532
rect 10896 2460 10912 2507
rect 10946 2460 10962 2507
rect 10896 2436 10962 2460
rect 10896 2388 10912 2436
rect 10946 2388 10962 2436
rect 10896 2365 10962 2388
rect 344 2293 410 2316
rect 344 2244 360 2293
rect 394 2244 410 2293
rect 344 2239 410 2244
rect 10896 2316 10912 2365
rect 10946 2316 10962 2365
rect 10896 2294 10962 2316
rect 10896 2260 10912 2294
rect 10946 2260 10962 2294
rect 10896 2239 10962 2260
rect 344 2223 10962 2239
rect 344 2189 360 2223
rect 394 2189 429 2223
rect 490 2189 498 2223
rect 562 2189 567 2223
rect 634 2189 636 2223
rect 670 2189 705 2223
rect 739 2189 774 2223
rect 808 2189 843 2223
rect 877 2189 912 2223
rect 946 2189 981 2223
rect 1015 2189 1050 2223
rect 1103 2189 1119 2223
rect 1175 2189 1188 2223
rect 1247 2189 1256 2223
rect 1290 2189 1324 2223
rect 1358 2189 1392 2223
rect 1426 2189 1458 2223
rect 1494 2189 1528 2223
rect 1564 2189 1596 2223
rect 1636 2189 1664 2223
rect 1698 2189 1732 2223
rect 1766 2189 1800 2223
rect 1834 2189 1868 2223
rect 1902 2189 1912 2223
rect 1970 2189 1984 2223
rect 2038 2189 2056 2223
rect 2106 2189 2140 2223
rect 2174 2189 2208 2223
rect 2242 2189 2276 2223
rect 2310 2189 2317 2223
rect 2378 2189 2389 2223
rect 2446 2189 2461 2223
rect 2514 2189 2548 2223
rect 2582 2189 2616 2223
rect 2650 2189 2684 2223
rect 2718 2189 2752 2223
rect 2815 2189 2820 2223
rect 2887 2189 2888 2223
rect 2922 2189 2925 2223
rect 2990 2189 3024 2223
rect 3058 2189 3092 2223
rect 3126 2189 3160 2223
rect 3194 2189 3219 2223
rect 3262 2189 3291 2223
rect 3330 2189 3363 2223
rect 3398 2189 3432 2223
rect 3469 2189 3500 2223
rect 3541 2189 3568 2223
rect 3613 2189 3636 2223
rect 3670 2189 3704 2223
rect 3738 2189 3772 2223
rect 3806 2189 3840 2223
rect 3874 2189 3908 2223
rect 3942 2189 3976 2223
rect 4027 2189 4044 2223
rect 4099 2189 4112 2223
rect 4171 2189 4180 2223
rect 4214 2189 4248 2223
rect 4282 2189 4316 2223
rect 4350 2189 4384 2223
rect 4418 2189 4452 2223
rect 4486 2189 4488 2223
rect 4554 2189 4560 2223
rect 4622 2189 4632 2223
rect 4690 2189 4724 2223
rect 4758 2189 4792 2223
rect 4826 2189 4860 2223
rect 4916 2189 4928 2223
rect 4988 2189 4996 2223
rect 5060 2189 5064 2223
rect 5098 2189 5132 2223
rect 5166 2189 5200 2223
rect 5234 2189 5268 2223
rect 5302 2189 5336 2223
rect 5381 2189 5404 2223
rect 5453 2189 5472 2223
rect 5525 2189 5540 2223
rect 5574 2189 5608 2223
rect 5642 2189 5676 2223
rect 5710 2189 5741 2223
rect 5778 2189 5812 2223
rect 5847 2189 5880 2223
rect 5919 2189 5948 2223
rect 5982 2189 6016 2223
rect 6050 2189 6084 2223
rect 6118 2189 6152 2223
rect 6186 2189 6211 2223
rect 6254 2189 6283 2223
rect 6322 2189 6355 2223
rect 6390 2189 6424 2223
rect 6458 2189 6492 2223
rect 6526 2189 6560 2223
rect 6594 2189 6628 2223
rect 6663 2189 6696 2223
rect 6735 2189 6764 2223
rect 6807 2189 6832 2223
rect 6879 2189 6900 2223
rect 6951 2189 6968 2223
rect 7023 2189 7036 2223
rect 7095 2189 7104 2223
rect 7167 2189 7172 2223
rect 7239 2189 7240 2223
rect 7274 2189 7277 2223
rect 7342 2189 7349 2223
rect 7410 2189 7421 2223
rect 7478 2189 7493 2223
rect 7546 2189 7565 2223
rect 7614 2189 7637 2223
rect 7682 2189 7709 2223
rect 7750 2189 7781 2223
rect 7818 2189 7852 2223
rect 7887 2189 7920 2223
rect 7959 2189 7988 2223
rect 8031 2189 8056 2223
rect 8103 2189 8124 2223
rect 8175 2189 8192 2223
rect 8247 2189 8260 2223
rect 8319 2189 8328 2223
rect 8391 2189 8396 2223
rect 8463 2189 8464 2223
rect 8498 2189 8501 2223
rect 8566 2189 8573 2223
rect 8634 2189 8645 2223
rect 8702 2189 8717 2223
rect 8770 2189 8789 2223
rect 8838 2189 8861 2223
rect 8906 2189 8933 2223
rect 8974 2189 9005 2223
rect 9042 2189 9076 2223
rect 9111 2189 9144 2223
rect 9183 2189 9212 2223
rect 9255 2189 9280 2223
rect 9327 2189 9348 2223
rect 9399 2189 9416 2223
rect 9471 2189 9484 2223
rect 9543 2189 9552 2223
rect 9615 2189 9620 2223
rect 9687 2189 9688 2223
rect 9722 2189 9725 2223
rect 9790 2189 9797 2223
rect 9858 2189 9869 2223
rect 9926 2189 9941 2223
rect 9994 2189 10013 2223
rect 10062 2189 10085 2223
rect 10130 2189 10157 2223
rect 10198 2189 10229 2223
rect 10266 2189 10300 2223
rect 10335 2189 10368 2223
rect 10407 2189 10436 2223
rect 10479 2189 10504 2223
rect 10551 2189 10572 2223
rect 10623 2189 10640 2223
rect 10695 2189 10708 2223
rect 10767 2189 10776 2223
rect 10839 2189 10844 2223
rect 10911 2189 10912 2223
rect 10946 2189 10962 2223
rect 344 2173 10962 2189
rect 11482 3916 11506 3950
rect 11540 3916 11564 3950
rect 14740 4000 14774 4017
rect 14808 4000 14844 4017
rect 14878 4000 14914 4017
rect 14948 4000 14984 4017
rect 15018 4000 15054 4017
rect 15088 4000 15124 4017
rect 15158 4000 15194 4017
rect 15228 4000 15264 4017
rect 15298 4000 15334 4017
rect 15368 4000 15404 4034
rect 15438 4016 15474 4034
rect 15439 4000 15474 4016
rect 15508 4012 15544 4034
rect 15578 4012 15614 4034
rect 15648 4012 15684 4034
rect 15518 4000 15544 4012
rect 15594 4000 15614 4012
rect 15670 4000 15684 4012
rect 15718 4016 15733 4034
rect 15788 4016 15819 4034
rect 15718 4000 15754 4016
rect 15788 4000 15824 4016
rect 15858 4000 15894 4034
rect 15939 4016 15964 4034
rect 16025 4016 16033 4050
rect 15928 4000 15964 4016
rect 15998 4000 16033 4016
rect 14740 3982 15405 4000
rect 15439 3982 15484 4000
rect 14740 3978 15484 3982
rect 15518 3978 15560 4000
rect 15594 3978 15636 4000
rect 15670 3978 16033 4000
rect 14740 3966 15733 3978
rect 15767 3966 15819 3978
rect 15853 3966 15905 3978
rect 15939 3966 15991 3978
rect 14740 3932 14774 3966
rect 14808 3932 14844 3966
rect 14878 3932 14914 3966
rect 14948 3932 14984 3966
rect 15018 3932 15054 3966
rect 15088 3932 15124 3966
rect 15158 3932 15194 3966
rect 15228 3932 15264 3966
rect 15298 3932 15334 3966
rect 15368 3932 15404 3966
rect 15438 3932 15474 3966
rect 15508 3932 15544 3966
rect 15578 3932 15614 3966
rect 15648 3932 15684 3966
rect 15718 3944 15733 3966
rect 15788 3944 15819 3966
rect 15718 3932 15754 3944
rect 15788 3932 15824 3944
rect 15858 3932 15894 3966
rect 15939 3944 15964 3966
rect 16025 3944 16033 3978
rect 15928 3932 15964 3944
rect 15998 3932 16033 3944
rect 11482 3881 11564 3916
rect 11626 3908 11728 3924
rect 14528 3908 14630 3924
rect 11482 3844 11506 3881
rect 11540 3844 11564 3881
rect 11660 3874 11694 3908
rect 14562 3874 14596 3908
rect 14740 3898 15484 3932
rect 15518 3898 15560 3932
rect 15594 3898 15636 3932
rect 15670 3906 16033 3932
rect 15670 3898 15733 3906
rect 15767 3898 15819 3906
rect 15853 3898 15905 3906
rect 15939 3898 15991 3906
rect 11626 3858 11728 3874
rect 14528 3858 14630 3874
rect 14740 3864 14774 3898
rect 14808 3864 14844 3898
rect 14878 3864 14914 3898
rect 14948 3864 14984 3898
rect 15018 3864 15054 3898
rect 15088 3864 15124 3898
rect 15158 3864 15194 3898
rect 15228 3864 15264 3898
rect 15298 3864 15334 3898
rect 15368 3864 15404 3898
rect 15438 3864 15474 3898
rect 15508 3864 15544 3898
rect 15578 3864 15614 3898
rect 15648 3864 15684 3898
rect 15718 3872 15733 3898
rect 15788 3872 15819 3898
rect 15718 3864 15754 3872
rect 15788 3864 15824 3872
rect 15858 3864 15894 3898
rect 15939 3872 15964 3898
rect 16025 3872 16033 3906
rect 15928 3864 15964 3872
rect 15998 3864 16033 3872
rect 14740 3859 16033 3864
rect 11482 3812 11564 3844
rect 11482 3772 11506 3812
rect 11540 3772 11564 3812
rect 11482 3743 11564 3772
rect 14740 3830 15554 3859
rect 15588 3830 15626 3859
rect 15660 3834 16033 3859
rect 15660 3830 15733 3834
rect 15767 3830 15819 3834
rect 15853 3830 15905 3834
rect 15939 3830 15991 3834
rect 14740 3796 14774 3830
rect 14808 3796 14844 3830
rect 14878 3796 14914 3830
rect 14948 3796 14984 3830
rect 15018 3796 15054 3830
rect 15088 3796 15124 3830
rect 15158 3796 15194 3830
rect 15228 3796 15264 3830
rect 15298 3796 15334 3830
rect 15368 3796 15404 3830
rect 15438 3796 15474 3830
rect 15508 3796 15544 3830
rect 15588 3825 15614 3830
rect 15660 3825 15684 3830
rect 15578 3796 15614 3825
rect 15648 3796 15684 3825
rect 15718 3800 15733 3830
rect 15788 3800 15819 3830
rect 15718 3796 15754 3800
rect 15788 3796 15824 3800
rect 15858 3796 15894 3830
rect 15939 3800 15964 3830
rect 16025 3800 16033 3834
rect 15928 3796 15964 3800
rect 15998 3796 16033 3800
rect 11626 3754 11728 3770
rect 14528 3754 14630 3770
rect 14740 3762 16033 3796
rect 11482 3700 11506 3743
rect 11540 3700 11564 3743
rect 11660 3720 11694 3754
rect 14562 3720 14596 3754
rect 14740 3728 14774 3762
rect 14808 3728 14844 3762
rect 14878 3728 14914 3762
rect 14948 3728 14984 3762
rect 15018 3728 15054 3762
rect 15088 3728 15124 3762
rect 15158 3728 15194 3762
rect 15228 3728 15264 3762
rect 15298 3728 15334 3762
rect 15368 3728 15404 3762
rect 15438 3728 15474 3762
rect 15508 3728 15544 3762
rect 15578 3728 15614 3762
rect 15648 3728 15684 3762
rect 15718 3728 15733 3762
rect 15788 3728 15819 3762
rect 15858 3728 15894 3762
rect 15939 3728 15964 3762
rect 16025 3728 16033 3762
rect 11626 3704 11728 3720
rect 14528 3704 14630 3720
rect 11482 3674 11564 3700
rect 11482 3628 11506 3674
rect 11540 3628 11564 3674
rect 11482 3605 11564 3628
rect 14740 3694 16033 3728
rect 14740 3660 14774 3694
rect 14808 3660 14844 3694
rect 14878 3660 14914 3694
rect 14948 3660 14984 3694
rect 15018 3660 15054 3694
rect 15088 3660 15124 3694
rect 15158 3660 15194 3694
rect 15228 3660 15264 3694
rect 15298 3660 15334 3694
rect 15368 3660 15404 3694
rect 15438 3660 15474 3694
rect 15508 3660 15544 3694
rect 15578 3660 15614 3694
rect 15648 3660 15684 3694
rect 15718 3690 15754 3694
rect 15788 3690 15824 3694
rect 15718 3660 15733 3690
rect 15788 3660 15819 3690
rect 15858 3660 15894 3694
rect 15928 3690 15964 3694
rect 15998 3690 16033 3694
rect 15939 3660 15964 3690
rect 14740 3656 15733 3660
rect 15767 3656 15819 3660
rect 15853 3656 15905 3660
rect 15939 3656 15991 3660
rect 16025 3656 16033 3690
rect 14740 3626 16033 3656
rect 11482 3556 11506 3605
rect 11540 3556 11564 3605
rect 11626 3600 11728 3616
rect 14528 3600 14630 3616
rect 11660 3566 11694 3600
rect 14562 3566 14596 3600
rect 14740 3592 14774 3626
rect 14808 3592 14844 3626
rect 14878 3592 14914 3626
rect 14948 3592 14984 3626
rect 15018 3592 15054 3626
rect 15088 3592 15124 3626
rect 15158 3592 15194 3626
rect 15228 3592 15264 3626
rect 15298 3592 15334 3626
rect 15368 3592 15404 3626
rect 15438 3592 15474 3626
rect 15508 3592 15544 3626
rect 15578 3592 15614 3626
rect 15648 3592 15684 3626
rect 15718 3618 15754 3626
rect 15788 3618 15824 3626
rect 15718 3592 15733 3618
rect 15788 3592 15819 3618
rect 15858 3592 15894 3626
rect 15928 3618 15964 3626
rect 15998 3618 16033 3626
rect 15939 3592 15964 3618
rect 14740 3584 15733 3592
rect 15767 3584 15819 3592
rect 15853 3584 15905 3592
rect 15939 3584 15991 3592
rect 16025 3584 16033 3618
rect 11482 3536 11564 3556
rect 11626 3550 11728 3566
rect 14528 3550 14630 3566
rect 14740 3558 16033 3584
rect 11482 3484 11506 3536
rect 11540 3484 11564 3536
rect 11482 3467 11564 3484
rect 11482 3412 11506 3467
rect 11540 3412 11564 3467
rect 14740 3524 14774 3558
rect 14808 3524 14844 3558
rect 14878 3524 14914 3558
rect 14948 3524 14984 3558
rect 15018 3524 15054 3558
rect 15088 3524 15124 3558
rect 15158 3524 15194 3558
rect 15228 3524 15264 3558
rect 15298 3524 15334 3558
rect 15368 3524 15404 3558
rect 15438 3524 15474 3558
rect 15508 3524 15544 3558
rect 15578 3524 15614 3558
rect 15648 3524 15684 3558
rect 15718 3546 15754 3558
rect 15788 3546 15824 3558
rect 15718 3524 15733 3546
rect 15788 3524 15819 3546
rect 15858 3524 15894 3558
rect 15928 3546 15964 3558
rect 15998 3546 16033 3558
rect 15939 3524 15964 3546
rect 14740 3512 15733 3524
rect 15767 3512 15819 3524
rect 15853 3512 15905 3524
rect 15939 3512 15991 3524
rect 16025 3512 16033 3546
rect 14740 3490 16033 3512
rect 11626 3446 11728 3462
rect 14528 3446 14630 3462
rect 14740 3456 14774 3490
rect 14808 3456 14844 3490
rect 14878 3456 14914 3490
rect 14948 3456 14984 3490
rect 15018 3456 15054 3490
rect 15088 3456 15124 3490
rect 15158 3456 15194 3490
rect 15228 3456 15264 3490
rect 15298 3456 15334 3490
rect 15368 3456 15404 3490
rect 15438 3456 15474 3490
rect 15508 3456 15544 3490
rect 15578 3456 15614 3490
rect 15648 3456 15684 3490
rect 15718 3474 15754 3490
rect 15788 3474 15824 3490
rect 15718 3456 15733 3474
rect 15788 3456 15819 3474
rect 15858 3456 15894 3490
rect 15928 3474 15964 3490
rect 15998 3474 16033 3490
rect 15939 3456 15964 3474
rect 11660 3412 11694 3446
rect 14562 3412 14596 3446
rect 14740 3440 15733 3456
rect 15767 3440 15819 3456
rect 15853 3440 15905 3456
rect 15939 3440 15991 3456
rect 16025 3440 16033 3474
rect 14740 3422 16033 3440
rect 11482 3398 11564 3412
rect 11482 3340 11506 3398
rect 11540 3340 11564 3398
rect 11626 3396 11728 3412
rect 14528 3396 14630 3412
rect 11482 3329 11564 3340
rect 11482 3268 11506 3329
rect 11540 3268 11564 3329
rect 14740 3388 14774 3422
rect 14808 3388 14844 3422
rect 14878 3388 14914 3422
rect 14948 3388 14984 3422
rect 15018 3388 15054 3422
rect 15088 3388 15124 3422
rect 15158 3388 15194 3422
rect 15228 3388 15264 3422
rect 15298 3388 15334 3422
rect 15368 3388 15404 3422
rect 15438 3388 15474 3422
rect 15508 3388 15544 3422
rect 15578 3388 15614 3422
rect 15648 3388 15684 3422
rect 15718 3402 15754 3422
rect 15788 3402 15824 3422
rect 15718 3388 15733 3402
rect 15788 3388 15819 3402
rect 15858 3388 15894 3422
rect 15928 3402 15964 3422
rect 15998 3402 16033 3422
rect 15939 3388 15964 3402
rect 14740 3368 15733 3388
rect 15767 3368 15819 3388
rect 15853 3368 15905 3388
rect 15939 3368 15991 3388
rect 16025 3368 16033 3402
rect 14740 3354 16033 3368
rect 14740 3320 14774 3354
rect 14808 3320 14844 3354
rect 14878 3320 14914 3354
rect 14948 3320 14984 3354
rect 15018 3320 15054 3354
rect 15088 3320 15124 3354
rect 15158 3320 15194 3354
rect 15228 3320 15264 3354
rect 15298 3320 15334 3354
rect 15368 3320 15404 3354
rect 15438 3320 15474 3354
rect 15508 3320 15544 3354
rect 15578 3320 15614 3354
rect 15648 3320 15684 3354
rect 15718 3330 15754 3354
rect 15788 3330 15824 3354
rect 15718 3320 15733 3330
rect 15788 3320 15819 3330
rect 15858 3320 15894 3354
rect 15928 3330 15964 3354
rect 15998 3330 16033 3354
rect 15939 3320 15964 3330
rect 11626 3292 11728 3308
rect 14528 3292 14630 3308
rect 14740 3296 15733 3320
rect 15767 3296 15819 3320
rect 15853 3296 15905 3320
rect 15939 3296 15991 3320
rect 16025 3296 16033 3330
rect 11482 3260 11564 3268
rect 11482 3196 11506 3260
rect 11540 3196 11564 3260
rect 11660 3258 11694 3292
rect 14562 3258 14596 3292
rect 14740 3286 16033 3296
rect 11626 3242 11728 3258
rect 14528 3242 14630 3258
rect 14740 3252 14774 3286
rect 14808 3252 14844 3286
rect 14878 3252 14914 3286
rect 14948 3252 14984 3286
rect 15018 3252 15054 3286
rect 15088 3252 15124 3286
rect 15158 3252 15194 3286
rect 15228 3252 15264 3286
rect 15298 3252 15334 3286
rect 15368 3252 15404 3286
rect 15438 3252 15474 3286
rect 15508 3252 15544 3286
rect 15578 3252 15614 3286
rect 15648 3252 15684 3286
rect 15718 3258 15754 3286
rect 15788 3258 15824 3286
rect 15718 3252 15733 3258
rect 15788 3252 15819 3258
rect 15858 3252 15894 3286
rect 15928 3258 15964 3286
rect 15998 3258 16033 3286
rect 15939 3252 15964 3258
rect 11482 3191 11564 3196
rect 11482 3124 11506 3191
rect 11540 3124 11564 3191
rect 14740 3224 15733 3252
rect 15767 3224 15819 3252
rect 15853 3224 15905 3252
rect 15939 3224 15991 3252
rect 16025 3224 16033 3258
rect 14740 3218 16033 3224
rect 14740 3184 14774 3218
rect 14808 3184 14844 3218
rect 14878 3184 14914 3218
rect 14948 3184 14984 3218
rect 15018 3184 15054 3218
rect 15088 3184 15124 3218
rect 15158 3184 15194 3218
rect 15228 3184 15264 3218
rect 15298 3184 15334 3218
rect 15368 3184 15404 3218
rect 15438 3184 15474 3218
rect 15508 3184 15544 3218
rect 15578 3184 15614 3218
rect 15648 3184 15684 3218
rect 15718 3186 15754 3218
rect 15788 3186 15824 3218
rect 15718 3184 15733 3186
rect 15788 3184 15819 3186
rect 15858 3184 15894 3218
rect 15928 3186 15964 3218
rect 15998 3186 16033 3218
rect 15939 3184 15964 3186
rect 11626 3138 11728 3154
rect 14528 3138 14630 3154
rect 14740 3152 15733 3184
rect 15767 3152 15819 3184
rect 15853 3152 15905 3184
rect 15939 3152 15991 3184
rect 16025 3152 16033 3186
rect 14740 3150 16033 3152
rect 11482 3122 11564 3124
rect 11482 3088 11506 3122
rect 11540 3088 11564 3122
rect 11660 3104 11694 3138
rect 14562 3104 14596 3138
rect 14740 3116 14774 3150
rect 14808 3116 14844 3150
rect 14878 3116 14914 3150
rect 14948 3116 14984 3150
rect 15018 3116 15054 3150
rect 15088 3116 15124 3150
rect 15158 3116 15194 3150
rect 15228 3116 15264 3150
rect 15298 3116 15334 3150
rect 15368 3116 15404 3150
rect 15438 3116 15474 3150
rect 15508 3116 15544 3150
rect 15578 3116 15614 3150
rect 15648 3116 15684 3150
rect 15718 3116 15754 3150
rect 15788 3116 15824 3150
rect 15858 3116 15894 3150
rect 15928 3116 15964 3150
rect 15998 3116 16033 3150
rect 14740 3114 16033 3116
rect 11626 3088 11728 3104
rect 14528 3088 14630 3104
rect 11482 3086 11564 3088
rect 11482 3019 11506 3086
rect 11540 3019 11564 3086
rect 11482 3014 11564 3019
rect 11482 2950 11506 3014
rect 11540 2950 11564 3014
rect 14740 3082 15733 3114
rect 15767 3082 15819 3114
rect 15853 3082 15905 3114
rect 15939 3082 15991 3114
rect 14740 3048 14774 3082
rect 14808 3048 14844 3082
rect 14878 3048 14914 3082
rect 14948 3048 14984 3082
rect 15018 3048 15054 3082
rect 15088 3048 15124 3082
rect 15158 3048 15194 3082
rect 15228 3048 15264 3082
rect 15298 3048 15334 3082
rect 15368 3048 15404 3082
rect 15438 3048 15474 3082
rect 15508 3048 15544 3082
rect 15578 3048 15614 3082
rect 15648 3048 15684 3082
rect 15718 3080 15733 3082
rect 15788 3080 15819 3082
rect 15718 3048 15754 3080
rect 15788 3048 15824 3080
rect 15858 3048 15894 3082
rect 15939 3080 15964 3082
rect 16025 3080 16033 3114
rect 15928 3048 15964 3080
rect 15998 3048 16033 3080
rect 14740 3042 16033 3048
rect 14740 3014 15733 3042
rect 15767 3014 15819 3042
rect 15853 3014 15905 3042
rect 15939 3014 15991 3042
rect 11626 2984 11728 3000
rect 14528 2984 14630 3000
rect 11660 2950 11694 2984
rect 14562 2950 14596 2984
rect 14740 2980 14774 3014
rect 14808 2980 14844 3014
rect 14878 2980 14914 3014
rect 14948 2980 14984 3014
rect 15018 2980 15054 3014
rect 15088 2980 15124 3014
rect 15158 2980 15194 3014
rect 15228 2980 15264 3014
rect 15298 2980 15334 3014
rect 15368 2980 15404 3014
rect 15438 2980 15474 3014
rect 15508 2980 15544 3014
rect 15578 2980 15614 3014
rect 15648 2980 15684 3014
rect 15718 3008 15733 3014
rect 15788 3008 15819 3014
rect 15718 2980 15754 3008
rect 15788 2980 15824 3008
rect 15858 2980 15894 3014
rect 15939 3008 15964 3014
rect 16025 3008 16033 3042
rect 15928 2980 15964 3008
rect 15998 2980 16033 3008
rect 14740 2970 16033 2980
rect 11482 2942 11564 2950
rect 11482 2881 11506 2942
rect 11540 2881 11564 2942
rect 11626 2934 11728 2950
rect 14528 2934 14630 2950
rect 14740 2946 15733 2970
rect 15767 2946 15819 2970
rect 15853 2946 15905 2970
rect 15939 2946 15991 2970
rect 11482 2870 11564 2881
rect 11482 2812 11506 2870
rect 11540 2812 11564 2870
rect 14740 2912 14774 2946
rect 14808 2912 14844 2946
rect 14878 2912 14914 2946
rect 14948 2912 14984 2946
rect 15018 2912 15054 2946
rect 15088 2912 15124 2946
rect 15158 2912 15194 2946
rect 15228 2912 15264 2946
rect 15298 2912 15334 2946
rect 15368 2912 15404 2946
rect 15438 2912 15474 2946
rect 15508 2912 15544 2946
rect 15578 2912 15614 2946
rect 15648 2912 15684 2946
rect 15718 2936 15733 2946
rect 15788 2936 15819 2946
rect 15718 2912 15754 2936
rect 15788 2912 15824 2936
rect 15858 2912 15894 2946
rect 15939 2936 15964 2946
rect 16025 2936 16033 2970
rect 15928 2912 15964 2936
rect 15998 2912 16033 2936
rect 14740 2898 16033 2912
rect 14740 2878 15733 2898
rect 15767 2878 15819 2898
rect 15853 2878 15905 2898
rect 15939 2878 15991 2898
rect 11626 2830 11728 2846
rect 14528 2830 14630 2846
rect 14740 2844 14774 2878
rect 14808 2844 14844 2878
rect 14878 2844 14914 2878
rect 14948 2844 14984 2878
rect 15018 2844 15054 2878
rect 15088 2844 15124 2878
rect 15158 2844 15194 2878
rect 15228 2844 15264 2878
rect 15298 2844 15334 2878
rect 15368 2844 15404 2878
rect 15438 2844 15474 2878
rect 15508 2844 15544 2878
rect 15578 2844 15614 2878
rect 15648 2844 15684 2878
rect 15718 2864 15733 2878
rect 15788 2864 15819 2878
rect 15718 2844 15754 2864
rect 15788 2844 15824 2864
rect 15858 2844 15894 2878
rect 15939 2864 15964 2878
rect 16025 2864 16033 2898
rect 15928 2844 15964 2864
rect 15998 2844 16033 2864
rect 11482 2798 11564 2812
rect 11482 2743 11506 2798
rect 11540 2743 11564 2798
rect 11660 2796 11694 2830
rect 14562 2796 14596 2830
rect 14740 2826 16033 2844
rect 14740 2810 15733 2826
rect 15767 2810 15819 2826
rect 15853 2810 15905 2826
rect 15939 2810 15991 2826
rect 11626 2780 11728 2796
rect 14528 2780 14630 2796
rect 11482 2726 11564 2743
rect 11482 2674 11506 2726
rect 11540 2674 11564 2726
rect 14740 2776 14774 2810
rect 14808 2776 14844 2810
rect 14878 2776 14914 2810
rect 14948 2776 14984 2810
rect 15018 2776 15054 2810
rect 15088 2776 15124 2810
rect 15158 2776 15194 2810
rect 15228 2776 15264 2810
rect 15298 2776 15334 2810
rect 15368 2776 15404 2810
rect 15438 2776 15474 2810
rect 15508 2776 15544 2810
rect 15578 2776 15614 2810
rect 15648 2776 15684 2810
rect 15718 2792 15733 2810
rect 15788 2792 15819 2810
rect 15718 2776 15754 2792
rect 15788 2776 15824 2792
rect 15858 2776 15894 2810
rect 15939 2792 15964 2810
rect 16025 2792 16033 2826
rect 15928 2776 15964 2792
rect 15998 2776 16033 2792
rect 14740 2754 16033 2776
rect 14740 2742 15733 2754
rect 15767 2742 15819 2754
rect 15853 2742 15905 2754
rect 15939 2742 15991 2754
rect 14740 2708 14774 2742
rect 14808 2708 14844 2742
rect 14878 2708 14914 2742
rect 14948 2708 14984 2742
rect 15018 2708 15054 2742
rect 15088 2708 15124 2742
rect 15158 2708 15194 2742
rect 15228 2708 15264 2742
rect 15298 2708 15334 2742
rect 15368 2708 15404 2742
rect 15438 2708 15474 2742
rect 15508 2708 15544 2742
rect 15578 2708 15614 2742
rect 15648 2708 15684 2742
rect 15718 2720 15733 2742
rect 15788 2720 15819 2742
rect 15718 2708 15754 2720
rect 15788 2708 15824 2720
rect 15858 2708 15894 2742
rect 15939 2720 15964 2742
rect 16025 2720 16033 2754
rect 15928 2708 15964 2720
rect 15998 2708 16033 2720
rect 11626 2676 11728 2692
rect 14528 2676 14630 2692
rect 14740 2681 16033 2708
rect 11482 2654 11564 2674
rect 11482 2605 11506 2654
rect 11540 2605 11564 2654
rect 11660 2642 11694 2676
rect 14562 2642 14596 2676
rect 14740 2674 15733 2681
rect 15767 2674 15819 2681
rect 15853 2674 15905 2681
rect 15939 2674 15991 2681
rect 11626 2626 11728 2642
rect 14528 2626 14630 2642
rect 14740 2640 14774 2674
rect 14808 2640 14844 2674
rect 14878 2640 14914 2674
rect 14948 2640 14984 2674
rect 15018 2640 15054 2674
rect 15088 2640 15124 2674
rect 15158 2640 15194 2674
rect 15228 2640 15264 2674
rect 15298 2640 15334 2674
rect 15368 2640 15404 2674
rect 15438 2640 15474 2674
rect 15508 2640 15544 2674
rect 15578 2640 15614 2674
rect 15648 2640 15684 2674
rect 15718 2647 15733 2674
rect 15788 2647 15819 2674
rect 15718 2640 15754 2647
rect 15788 2640 15824 2647
rect 15858 2640 15894 2674
rect 15939 2647 15964 2674
rect 16025 2647 16033 2681
rect 15928 2640 15964 2647
rect 15998 2640 16033 2647
rect 11482 2582 11564 2605
rect 11482 2536 11506 2582
rect 11540 2536 11564 2582
rect 14740 2608 16033 2640
rect 14740 2606 15733 2608
rect 15767 2606 15819 2608
rect 15853 2606 15905 2608
rect 15939 2606 15991 2608
rect 14740 2572 14774 2606
rect 14808 2572 14844 2606
rect 14878 2572 14914 2606
rect 14948 2572 14984 2606
rect 15018 2572 15054 2606
rect 15088 2572 15124 2606
rect 15158 2572 15194 2606
rect 15228 2572 15264 2606
rect 15298 2572 15334 2606
rect 15368 2572 15404 2606
rect 15438 2572 15474 2606
rect 15508 2572 15544 2606
rect 15578 2572 15614 2606
rect 15648 2572 15684 2606
rect 15718 2574 15733 2606
rect 15788 2574 15819 2606
rect 15718 2572 15754 2574
rect 15788 2572 15824 2574
rect 15858 2572 15894 2606
rect 15939 2574 15964 2606
rect 16025 2574 16033 2608
rect 15928 2572 15964 2574
rect 15998 2572 16033 2574
rect 14740 2538 16033 2572
rect 11482 2510 11564 2536
rect 11626 2522 11728 2538
rect 14528 2522 14630 2538
rect 11482 2467 11506 2510
rect 11540 2467 11564 2510
rect 11660 2488 11694 2522
rect 14562 2488 14596 2522
rect 14740 2504 14774 2538
rect 14808 2504 14844 2538
rect 14878 2504 14914 2538
rect 14948 2504 14984 2538
rect 15018 2504 15054 2538
rect 15088 2504 15124 2538
rect 15158 2504 15194 2538
rect 15228 2504 15264 2538
rect 15298 2504 15334 2538
rect 15368 2504 15404 2538
rect 15438 2504 15474 2538
rect 15508 2504 15544 2538
rect 15578 2504 15614 2538
rect 15648 2504 15684 2538
rect 15718 2535 15754 2538
rect 15788 2535 15824 2538
rect 15718 2504 15733 2535
rect 15788 2504 15819 2535
rect 15858 2504 15894 2538
rect 15928 2535 15964 2538
rect 15998 2535 16033 2538
rect 15939 2504 15964 2535
rect 14740 2501 15733 2504
rect 15767 2501 15819 2504
rect 15853 2501 15905 2504
rect 15939 2501 15991 2504
rect 16025 2501 16033 2535
rect 11626 2472 11728 2488
rect 14528 2472 14630 2488
rect 11482 2438 11564 2467
rect 11482 2397 11506 2438
rect 11540 2397 11564 2438
rect 11482 2366 11564 2397
rect 14740 2470 16033 2501
rect 14740 2436 14774 2470
rect 14808 2436 14844 2470
rect 14878 2436 14914 2470
rect 14948 2436 14984 2470
rect 15018 2436 15054 2470
rect 15088 2436 15124 2470
rect 15158 2436 15194 2470
rect 15228 2436 15264 2470
rect 15298 2436 15334 2470
rect 15368 2436 15404 2470
rect 15438 2436 15474 2470
rect 15508 2436 15544 2470
rect 15578 2436 15614 2470
rect 15648 2436 15684 2470
rect 15718 2462 15754 2470
rect 15788 2462 15824 2470
rect 15718 2436 15733 2462
rect 15788 2436 15819 2462
rect 15858 2436 15894 2470
rect 15928 2462 15964 2470
rect 15998 2462 16033 2470
rect 15939 2436 15964 2462
rect 14740 2428 15733 2436
rect 15767 2428 15819 2436
rect 15853 2428 15905 2436
rect 15939 2428 15991 2436
rect 16025 2428 16033 2462
rect 14740 2402 16033 2428
rect 11626 2368 11728 2384
rect 14528 2368 14630 2384
rect 14740 2368 14774 2402
rect 14808 2368 14844 2402
rect 14878 2368 14914 2402
rect 14948 2368 14984 2402
rect 15018 2368 15054 2402
rect 15088 2368 15124 2402
rect 15158 2368 15194 2402
rect 15228 2368 15264 2402
rect 15298 2368 15334 2402
rect 15368 2368 15404 2402
rect 15438 2368 15474 2402
rect 15508 2368 15544 2402
rect 15578 2368 15614 2402
rect 15648 2368 15684 2402
rect 15718 2389 15754 2402
rect 15788 2389 15824 2402
rect 15718 2368 15733 2389
rect 15788 2368 15819 2389
rect 15858 2368 15894 2402
rect 15928 2389 15964 2402
rect 15998 2389 16033 2402
rect 15939 2368 15964 2389
rect 11482 2327 11506 2366
rect 11540 2327 11564 2366
rect 11660 2334 11694 2368
rect 14562 2334 14596 2368
rect 14740 2355 15733 2368
rect 15767 2355 15819 2368
rect 15853 2355 15905 2368
rect 15939 2355 15991 2368
rect 16025 2355 16033 2389
rect 14740 2334 16033 2355
rect 11482 2294 11564 2327
rect 11626 2318 11728 2334
rect 14528 2318 14630 2334
rect 11482 2257 11506 2294
rect 11540 2257 11564 2294
rect 11482 2222 11564 2257
rect 14740 2300 14774 2334
rect 14808 2300 14844 2334
rect 14878 2300 14914 2334
rect 14948 2300 14984 2334
rect 15018 2300 15054 2334
rect 15088 2300 15124 2334
rect 15158 2300 15194 2334
rect 15228 2300 15264 2334
rect 15298 2300 15334 2334
rect 15368 2300 15404 2334
rect 15438 2300 15474 2334
rect 15508 2300 15544 2334
rect 15578 2300 15614 2334
rect 15648 2300 15684 2334
rect 15718 2316 15754 2334
rect 15788 2316 15824 2334
rect 15718 2300 15733 2316
rect 15788 2300 15819 2316
rect 15858 2300 15894 2334
rect 15928 2316 15964 2334
rect 15998 2316 16033 2334
rect 15939 2300 15964 2316
rect 14740 2282 15733 2300
rect 15767 2282 15819 2300
rect 15853 2282 15905 2300
rect 15939 2282 15991 2300
rect 16025 2282 16033 2316
rect 14740 2266 16033 2282
rect 14740 2232 14774 2266
rect 14808 2232 14844 2266
rect 14878 2232 14914 2266
rect 14948 2232 14984 2266
rect 15018 2232 15054 2266
rect 15088 2232 15124 2266
rect 15158 2232 15194 2266
rect 15228 2232 15264 2266
rect 15298 2232 15334 2266
rect 15368 2232 15404 2266
rect 15438 2232 15474 2266
rect 15508 2232 15544 2266
rect 15578 2232 15614 2266
rect 15648 2232 15684 2266
rect 15718 2243 15754 2266
rect 15788 2243 15824 2266
rect 15718 2232 15733 2243
rect 15788 2232 15819 2243
rect 15858 2232 15894 2266
rect 15928 2243 15964 2266
rect 15998 2243 16033 2266
rect 15939 2232 15964 2243
rect 11482 2187 11506 2222
rect 11540 2187 11564 2222
rect 11626 2214 11728 2230
rect 14528 2214 14630 2230
rect 11482 2151 11564 2187
rect 11660 2180 11694 2214
rect 14562 2180 14596 2214
rect 14740 2209 15733 2232
rect 15767 2209 15819 2232
rect 15853 2209 15905 2232
rect 15939 2209 15991 2232
rect 16025 2209 16033 2243
rect 14740 2198 16033 2209
rect 11626 2164 11728 2180
rect 14528 2164 14630 2180
rect 14740 2164 14774 2198
rect 14808 2164 14844 2198
rect 14878 2164 14914 2198
rect 14948 2164 14984 2198
rect 15018 2164 15054 2198
rect 15088 2164 15124 2198
rect 15158 2164 15194 2198
rect 15228 2164 15264 2198
rect 15298 2164 15334 2198
rect 15368 2164 15404 2198
rect 15438 2164 15474 2198
rect 15508 2164 15544 2198
rect 15578 2164 15614 2198
rect 15648 2164 15684 2198
rect 15718 2170 15754 2198
rect 15788 2170 15824 2198
rect 15718 2164 15733 2170
rect 15788 2164 15819 2170
rect 15858 2164 15894 2198
rect 15928 2170 15964 2198
rect 15998 2170 16033 2198
rect 15939 2164 15964 2170
rect 6659 2110 6698 2144
rect 6732 2110 6771 2144
rect 6805 2110 6844 2144
rect 6878 2110 6917 2144
rect 6951 2110 6990 2144
rect 7024 2110 7063 2144
rect 7097 2110 7136 2144
rect 7170 2110 7209 2144
rect 7243 2110 7282 2144
rect 7316 2110 7355 2144
rect 7389 2110 7428 2144
rect 7462 2110 7501 2144
rect 7535 2110 7574 2144
rect 7608 2110 7647 2144
rect 7681 2110 7720 2144
rect 7754 2110 7792 2144
rect 7826 2110 7864 2144
rect 7898 2110 7936 2144
rect 7970 2110 8008 2144
rect 8042 2110 8080 2144
rect 8114 2110 8152 2144
rect 8186 2110 8224 2144
rect 8258 2110 8296 2144
rect 8330 2110 8368 2144
rect 8402 2110 8440 2144
rect 8474 2110 8512 2144
rect 8546 2110 8584 2144
rect 8618 2110 8656 2144
rect 8690 2110 8728 2144
rect 8762 2110 8800 2144
rect 8834 2110 8872 2144
rect 8906 2110 8944 2144
rect 8978 2110 9016 2144
rect 9050 2110 9088 2144
rect 9122 2110 9160 2144
rect 9194 2110 9232 2144
rect 9266 2110 9304 2144
rect 9338 2110 9376 2144
rect 9410 2110 9448 2144
rect 9482 2110 9520 2144
rect 9554 2110 9592 2144
rect 9626 2110 9664 2144
rect 9698 2110 9736 2144
rect 9770 2110 9808 2144
rect 9842 2110 9880 2144
rect 9914 2110 9952 2144
rect 9986 2110 10024 2144
rect 10058 2110 10096 2144
rect 10130 2110 10168 2144
rect 10202 2110 10240 2144
rect 10274 2110 10312 2144
rect 10346 2110 10384 2144
rect 10418 2110 10456 2144
rect 10490 2110 10528 2144
rect 10562 2110 10600 2144
rect 10634 2110 10672 2144
rect 10706 2110 10744 2144
rect 10778 2110 10816 2144
rect 10850 2110 10888 2144
rect 11482 2116 11506 2151
rect 11540 2116 11564 2151
rect 11482 2093 11564 2116
rect 14740 2136 15733 2164
rect 15767 2136 15819 2164
rect 15853 2136 15905 2164
rect 15939 2136 15991 2164
rect 16025 2136 16033 2170
rect 14740 2130 16033 2136
rect 14740 2096 14774 2130
rect 14808 2096 14844 2130
rect 14878 2096 14914 2130
rect 14948 2096 14984 2130
rect 15018 2096 15054 2130
rect 15088 2096 15124 2130
rect 15158 2096 15194 2130
rect 15228 2096 15264 2130
rect 15298 2096 15334 2130
rect 15368 2096 15404 2130
rect 15438 2096 15474 2130
rect 15508 2096 15544 2130
rect 15578 2096 15614 2130
rect 15648 2096 15684 2130
rect 15718 2097 15754 2130
rect 15788 2097 15824 2130
rect 15718 2096 15733 2097
rect 15788 2096 15819 2097
rect 15858 2096 15894 2130
rect 15928 2097 15964 2130
rect 15998 2097 16033 2130
rect 15939 2096 15964 2097
rect 11506 2085 11540 2093
rect 14740 2085 15733 2096
rect 336 2078 15733 2085
rect 336 2069 11506 2078
rect 11540 2069 15733 2078
rect 370 2060 405 2069
rect 394 2035 405 2060
rect 439 2035 449 2069
rect 508 2035 521 2069
rect 577 2035 593 2069
rect 646 2035 665 2069
rect 715 2035 750 2069
rect 784 2035 819 2069
rect 853 2035 888 2069
rect 922 2035 957 2069
rect 991 2035 1026 2069
rect 1060 2035 1069 2069
rect 1129 2035 1141 2069
rect 1198 2035 1213 2069
rect 1267 2035 1302 2069
rect 1336 2035 1371 2069
rect 1405 2035 1440 2069
rect 1492 2035 1509 2069
rect 1564 2035 1578 2069
rect 1636 2035 1647 2069
rect 1681 2035 1716 2069
rect 1750 2035 1785 2069
rect 1819 2035 1854 2069
rect 1888 2035 1912 2069
rect 1957 2035 1984 2069
rect 2026 2035 2056 2069
rect 2095 2035 2130 2069
rect 2164 2035 2199 2069
rect 2233 2035 2268 2069
rect 2302 2035 2317 2069
rect 2371 2035 2389 2069
rect 2440 2035 2461 2069
rect 2509 2035 2544 2069
rect 2578 2035 2613 2069
rect 2647 2035 2682 2069
rect 2716 2035 2751 2069
rect 2815 2035 2820 2069
rect 2887 2035 2889 2069
rect 2923 2035 2925 2069
rect 2992 2035 3027 2069
rect 3061 2035 3096 2069
rect 3130 2035 3165 2069
rect 3199 2035 3219 2069
rect 3268 2035 3291 2069
rect 3337 2035 3363 2069
rect 3406 2035 3435 2069
rect 3475 2035 3507 2069
rect 3544 2035 3579 2069
rect 3613 2035 3648 2069
rect 3682 2035 3717 2069
rect 3751 2035 3786 2069
rect 3820 2035 3855 2069
rect 3889 2035 3924 2069
rect 3958 2035 3993 2069
rect 4027 2035 4062 2069
rect 4099 2035 4131 2069
rect 4171 2035 4200 2069
rect 4234 2035 4269 2069
rect 4303 2035 4338 2069
rect 4372 2035 4407 2069
rect 4441 2035 4475 2069
rect 4522 2035 4543 2069
rect 4594 2035 4611 2069
rect 4666 2035 4679 2069
rect 4713 2035 4747 2069
rect 4781 2035 4815 2069
rect 4849 2035 4882 2069
rect 4917 2035 4951 2069
rect 4988 2035 5019 2069
rect 5060 2035 5087 2069
rect 5121 2035 5155 2069
rect 5189 2035 5223 2069
rect 5257 2035 5291 2069
rect 5325 2035 5347 2069
rect 5393 2035 5419 2069
rect 5461 2035 5491 2069
rect 5529 2035 5563 2069
rect 5597 2035 5631 2069
rect 5665 2035 5699 2069
rect 5733 2035 5741 2069
rect 5801 2035 5813 2069
rect 5869 2035 5885 2069
rect 5937 2035 5971 2069
rect 6005 2035 6039 2069
rect 6073 2035 6107 2069
rect 6141 2035 6175 2069
rect 6209 2035 6211 2069
rect 6277 2035 6283 2069
rect 6345 2035 6355 2069
rect 6413 2035 6447 2069
rect 6481 2035 6515 2069
rect 6549 2035 6583 2069
rect 6617 2035 6629 2069
rect 6685 2035 6701 2069
rect 6753 2035 6773 2069
rect 6821 2035 6845 2069
rect 6889 2035 6917 2069
rect 6957 2035 6989 2069
rect 7025 2035 7059 2069
rect 7095 2035 7127 2069
rect 7167 2035 7195 2069
rect 7239 2035 7263 2069
rect 7311 2035 7331 2069
rect 7383 2035 7399 2069
rect 7455 2035 7467 2069
rect 7527 2035 7535 2069
rect 7599 2035 7603 2069
rect 7705 2035 7709 2069
rect 7773 2035 7781 2069
rect 7841 2035 7853 2069
rect 7909 2035 7925 2069
rect 7977 2035 7997 2069
rect 8045 2035 8069 2069
rect 8113 2035 8141 2069
rect 8181 2035 8213 2069
rect 8249 2035 8283 2069
rect 8319 2035 8351 2069
rect 8391 2035 8419 2069
rect 8463 2035 8487 2069
rect 8535 2035 8555 2069
rect 8607 2035 8623 2069
rect 8679 2035 8691 2069
rect 8751 2035 8759 2069
rect 8823 2035 8827 2069
rect 8929 2035 8933 2069
rect 8997 2035 9005 2069
rect 9065 2035 9077 2069
rect 9133 2035 9149 2069
rect 9201 2035 9221 2069
rect 9269 2035 9293 2069
rect 9337 2035 9365 2069
rect 9405 2035 9437 2069
rect 9473 2035 9507 2069
rect 9543 2035 9575 2069
rect 9615 2035 9643 2069
rect 9687 2035 9711 2069
rect 9759 2035 9779 2069
rect 9831 2035 9847 2069
rect 9903 2035 9915 2069
rect 9975 2035 9983 2069
rect 10047 2035 10051 2069
rect 10153 2035 10157 2069
rect 10221 2035 10229 2069
rect 10289 2035 10301 2069
rect 10357 2035 10373 2069
rect 10425 2035 10445 2069
rect 10493 2035 10517 2069
rect 10561 2035 10589 2069
rect 10629 2035 10661 2069
rect 10697 2035 10731 2069
rect 10767 2035 10799 2069
rect 10839 2035 10867 2069
rect 10911 2035 10935 2069
rect 10969 2035 11003 2069
rect 11037 2035 11071 2069
rect 11105 2035 11139 2069
rect 11173 2035 11207 2069
rect 11241 2035 11275 2069
rect 11309 2035 11343 2069
rect 11377 2035 11411 2069
rect 11445 2035 11479 2069
rect 11540 2044 11547 2069
rect 11513 2035 11547 2044
rect 11581 2035 11608 2069
rect 11649 2035 11680 2069
rect 11717 2035 11751 2069
rect 11786 2035 11819 2069
rect 11858 2035 11887 2069
rect 11930 2035 11955 2069
rect 12002 2035 12023 2069
rect 12074 2035 12091 2069
rect 12146 2035 12159 2069
rect 12218 2035 12227 2069
rect 12290 2035 12295 2069
rect 12362 2035 12363 2069
rect 12397 2035 12400 2069
rect 12465 2035 12472 2069
rect 12533 2035 12544 2069
rect 12601 2035 12616 2069
rect 12669 2035 12688 2069
rect 12737 2035 12760 2069
rect 12805 2035 12832 2069
rect 12873 2035 12904 2069
rect 12941 2035 12975 2069
rect 13010 2035 13043 2069
rect 13082 2035 13111 2069
rect 13154 2035 13179 2069
rect 13226 2035 13247 2069
rect 13298 2035 13315 2069
rect 13370 2035 13383 2069
rect 13442 2035 13451 2069
rect 13514 2035 13519 2069
rect 13586 2035 13587 2069
rect 13621 2035 13624 2069
rect 13689 2035 13696 2069
rect 13757 2035 13768 2069
rect 13825 2035 13840 2069
rect 13893 2035 13912 2069
rect 13961 2035 13984 2069
rect 14029 2035 14056 2069
rect 14097 2035 14128 2069
rect 14165 2035 14199 2069
rect 14234 2035 14267 2069
rect 14306 2035 14335 2069
rect 14378 2035 14403 2069
rect 14450 2035 14471 2069
rect 14522 2035 14539 2069
rect 14594 2035 14607 2069
rect 14666 2035 14675 2069
rect 14738 2063 15733 2069
rect 15767 2063 15819 2096
rect 15853 2063 15905 2096
rect 15939 2063 15991 2096
rect 16025 2063 16033 2097
rect 14738 2062 16033 2063
rect 14738 2035 14774 2062
rect 336 2026 360 2035
rect 394 2028 14774 2035
rect 14808 2028 14844 2062
rect 14878 2028 14914 2062
rect 14948 2028 14984 2062
rect 15018 2028 15054 2062
rect 15088 2028 15124 2062
rect 15158 2028 15194 2062
rect 15228 2028 15264 2062
rect 15298 2028 15334 2062
rect 15368 2028 15404 2062
rect 15438 2028 15474 2062
rect 15508 2028 15544 2062
rect 15578 2028 15614 2062
rect 15648 2028 15684 2062
rect 15718 2028 15754 2062
rect 15788 2028 15824 2062
rect 15858 2028 15894 2062
rect 15928 2028 15964 2062
rect 15998 2028 16033 2062
rect 394 2026 16033 2028
rect 336 2024 16033 2026
rect 336 2019 15733 2024
rect 344 1988 410 2019
rect 344 1925 360 1988
rect 394 1925 410 1988
rect 13152 2001 15733 2019
rect 13152 1967 13194 2001
rect 13228 1967 13264 2001
rect 13298 1967 13334 2001
rect 13368 1967 13404 2001
rect 13438 1967 13474 2001
rect 13508 1967 13544 2001
rect 13578 1967 13614 2001
rect 13648 1967 13684 2001
rect 13718 1967 13754 2001
rect 13788 1967 13824 2001
rect 13858 1967 13894 2001
rect 13928 1967 13964 2001
rect 13998 1967 14034 2001
rect 14068 1967 14104 2001
rect 14138 1967 14174 2001
rect 14208 1967 14244 2001
rect 14278 1967 14314 2001
rect 14348 1967 14384 2001
rect 14418 1967 14454 2001
rect 14488 1967 14524 2001
rect 14558 1967 14594 2001
rect 14628 1967 14664 2001
rect 14698 1994 15733 2001
rect 15767 1994 15819 2024
rect 15853 1994 15905 2024
rect 15939 1994 15991 2024
rect 14698 1967 14774 1994
rect 13152 1960 14774 1967
rect 14808 1960 14844 1994
rect 14878 1960 14914 1994
rect 14948 1960 14984 1994
rect 15018 1960 15054 1994
rect 15088 1960 15124 1994
rect 15158 1960 15194 1994
rect 15228 1960 15264 1994
rect 15298 1960 15334 1994
rect 15368 1960 15404 1994
rect 15438 1960 15474 1994
rect 15508 1960 15544 1994
rect 15578 1960 15614 1994
rect 15648 1960 15684 1994
rect 15718 1990 15733 1994
rect 15788 1990 15819 1994
rect 15718 1960 15754 1990
rect 15788 1960 15824 1990
rect 15858 1960 15894 1994
rect 15939 1990 15964 1994
rect 16025 1990 16033 2024
rect 15928 1960 15964 1990
rect 15998 1960 16033 1990
rect 13152 1951 16033 1960
rect 344 1916 410 1925
rect 480 1924 582 1940
rect 3382 1924 3484 1940
rect 12884 1924 12986 1940
rect 13152 1931 15733 1951
rect 344 1855 360 1916
rect 394 1855 410 1916
rect 514 1890 548 1924
rect 3416 1890 3450 1924
rect 12918 1890 12952 1924
rect 13152 1897 13194 1931
rect 13228 1897 13264 1931
rect 13298 1897 13334 1931
rect 13368 1897 13404 1931
rect 13438 1897 13474 1931
rect 13508 1897 13544 1931
rect 13578 1897 13614 1931
rect 13648 1897 13684 1931
rect 13718 1897 13754 1931
rect 13788 1897 13824 1931
rect 13858 1897 13894 1931
rect 13928 1897 13964 1931
rect 13998 1897 14034 1931
rect 14068 1897 14104 1931
rect 14138 1897 14174 1931
rect 14208 1897 14244 1931
rect 14278 1897 14314 1931
rect 14348 1897 14384 1931
rect 14418 1897 14454 1931
rect 14488 1897 14524 1931
rect 14558 1897 14594 1931
rect 14628 1897 14664 1931
rect 14698 1926 15733 1931
rect 15767 1926 15819 1951
rect 15853 1926 15905 1951
rect 15939 1926 15991 1951
rect 14698 1897 14774 1926
rect 13152 1892 14774 1897
rect 14808 1892 14844 1926
rect 14878 1892 14914 1926
rect 14948 1892 14984 1926
rect 15018 1892 15054 1926
rect 15088 1892 15124 1926
rect 15158 1892 15194 1926
rect 15228 1892 15264 1926
rect 15298 1892 15334 1926
rect 15368 1892 15404 1926
rect 15438 1892 15474 1926
rect 15508 1892 15544 1926
rect 15578 1892 15614 1926
rect 15648 1892 15684 1926
rect 15718 1917 15733 1926
rect 15788 1917 15819 1926
rect 15718 1892 15754 1917
rect 15788 1892 15824 1917
rect 15858 1892 15894 1926
rect 15939 1917 15964 1926
rect 16025 1917 16033 1951
rect 15928 1892 15964 1917
rect 15998 1892 16033 1917
rect 480 1874 582 1890
rect 3382 1874 3484 1890
rect 12884 1874 12986 1890
rect 13152 1878 16033 1892
rect 344 1844 410 1855
rect 344 1785 360 1844
rect 394 1785 410 1844
rect 13152 1861 15733 1878
rect 13152 1847 13194 1861
rect 13228 1847 13264 1861
rect 13298 1847 13334 1861
rect 13368 1847 13404 1861
rect 13438 1847 13474 1861
rect 13152 1813 13168 1847
rect 13228 1827 13244 1847
rect 13298 1827 13320 1847
rect 13368 1827 13396 1847
rect 13438 1827 13472 1847
rect 13508 1827 13544 1861
rect 13578 1847 13614 1861
rect 13648 1847 13684 1861
rect 13718 1847 13754 1861
rect 13788 1847 13824 1861
rect 13858 1847 13894 1861
rect 13928 1847 13964 1861
rect 13582 1827 13614 1847
rect 13658 1827 13684 1847
rect 13734 1827 13754 1847
rect 13810 1827 13824 1847
rect 13885 1827 13894 1847
rect 13960 1827 13964 1847
rect 13998 1847 14034 1861
rect 14068 1847 14104 1861
rect 14138 1847 14174 1861
rect 14208 1847 14244 1861
rect 14278 1847 14314 1861
rect 14348 1847 14384 1861
rect 14418 1847 14454 1861
rect 13998 1827 14001 1847
rect 14068 1827 14076 1847
rect 14138 1827 14151 1847
rect 14208 1827 14226 1847
rect 14278 1827 14301 1847
rect 14348 1827 14376 1847
rect 14418 1827 14451 1847
rect 14488 1827 14524 1861
rect 14558 1847 14594 1861
rect 14628 1847 14664 1861
rect 14560 1827 14594 1847
rect 14635 1827 14664 1847
rect 14698 1858 15733 1861
rect 15767 1858 15819 1878
rect 15853 1858 15905 1878
rect 15939 1858 15991 1878
rect 14698 1827 14774 1858
rect 13202 1813 13244 1827
rect 13278 1813 13320 1827
rect 13354 1813 13396 1827
rect 13430 1813 13472 1827
rect 13506 1813 13548 1827
rect 13582 1813 13624 1827
rect 13658 1813 13700 1827
rect 13734 1813 13776 1827
rect 13810 1813 13851 1827
rect 13885 1813 13926 1827
rect 13960 1813 14001 1827
rect 14035 1813 14076 1827
rect 14110 1813 14151 1827
rect 14185 1813 14226 1827
rect 14260 1813 14301 1827
rect 14335 1813 14376 1827
rect 14410 1813 14451 1827
rect 14485 1813 14526 1827
rect 14560 1813 14601 1827
rect 14635 1824 14774 1827
rect 14808 1824 14844 1858
rect 14878 1824 14914 1858
rect 14948 1824 14984 1858
rect 15018 1824 15054 1858
rect 15088 1824 15124 1858
rect 15158 1824 15194 1858
rect 15228 1824 15264 1858
rect 15298 1824 15334 1858
rect 15368 1824 15404 1858
rect 15438 1824 15474 1858
rect 15508 1824 15544 1858
rect 15578 1824 15614 1858
rect 15648 1824 15684 1858
rect 15718 1844 15733 1858
rect 15788 1844 15819 1858
rect 15718 1824 15754 1844
rect 15788 1824 15824 1844
rect 15858 1824 15894 1858
rect 15939 1844 15964 1858
rect 16025 1844 16033 1878
rect 15928 1824 15964 1844
rect 15998 1824 16033 1844
rect 14635 1813 16033 1824
rect 13152 1805 16033 1813
rect 13152 1791 15733 1805
rect 344 1772 410 1785
rect 344 1715 360 1772
rect 394 1715 410 1772
rect 480 1770 582 1786
rect 3382 1770 3484 1786
rect 12884 1770 12986 1786
rect 514 1736 548 1770
rect 3416 1736 3450 1770
rect 12918 1736 12952 1770
rect 13152 1757 13194 1791
rect 13228 1757 13264 1791
rect 13298 1757 13334 1791
rect 13368 1757 13404 1791
rect 13438 1757 13474 1791
rect 13508 1757 13544 1791
rect 13578 1757 13614 1791
rect 13648 1757 13684 1791
rect 13718 1757 13754 1791
rect 13788 1757 13824 1791
rect 13858 1757 13894 1791
rect 13928 1757 13964 1791
rect 13998 1757 14034 1791
rect 14068 1757 14104 1791
rect 14138 1757 14174 1791
rect 14208 1757 14244 1791
rect 14278 1757 14314 1791
rect 14348 1757 14384 1791
rect 14418 1757 14454 1791
rect 14488 1757 14524 1791
rect 14558 1757 14594 1791
rect 14628 1757 14664 1791
rect 14698 1790 15733 1791
rect 15767 1790 15819 1805
rect 15853 1790 15905 1805
rect 15939 1790 15991 1805
rect 14698 1757 14774 1790
rect 13152 1756 14774 1757
rect 14808 1756 14844 1790
rect 14878 1756 14914 1790
rect 14948 1756 14984 1790
rect 15018 1756 15054 1790
rect 15088 1756 15124 1790
rect 15158 1756 15194 1790
rect 15228 1756 15264 1790
rect 15298 1756 15334 1790
rect 15368 1756 15404 1790
rect 15438 1756 15474 1790
rect 15508 1756 15544 1790
rect 15578 1756 15614 1790
rect 15648 1756 15684 1790
rect 15718 1771 15733 1790
rect 15788 1771 15819 1790
rect 15718 1756 15754 1771
rect 15788 1756 15824 1771
rect 15858 1756 15894 1790
rect 15939 1771 15964 1790
rect 16025 1771 16033 1805
rect 15928 1756 15964 1771
rect 15998 1756 16033 1771
rect 480 1720 582 1736
rect 3382 1720 3484 1736
rect 12884 1720 12986 1736
rect 13152 1732 16033 1756
rect 13152 1722 15733 1732
rect 15767 1722 15819 1732
rect 15853 1722 15905 1732
rect 15939 1722 15991 1732
rect 13152 1721 14774 1722
rect 344 1700 410 1715
rect 344 1645 360 1700
rect 394 1645 410 1700
rect 344 1628 410 1645
rect 13152 1687 13194 1721
rect 13228 1687 13264 1721
rect 13298 1687 13334 1721
rect 13368 1687 13404 1721
rect 13438 1687 13474 1721
rect 13508 1687 13544 1721
rect 13578 1687 13614 1721
rect 13648 1687 13684 1721
rect 13718 1687 13754 1721
rect 13788 1687 13824 1721
rect 13858 1687 13894 1721
rect 13928 1687 13964 1721
rect 13998 1687 14034 1721
rect 14068 1687 14104 1721
rect 14138 1687 14174 1721
rect 14208 1687 14244 1721
rect 14278 1687 14314 1721
rect 14348 1687 14384 1721
rect 14418 1687 14454 1721
rect 14488 1687 14524 1721
rect 14558 1687 14594 1721
rect 14628 1687 14664 1721
rect 14698 1688 14774 1721
rect 14808 1688 14844 1722
rect 14878 1688 14914 1722
rect 14948 1688 14984 1722
rect 15018 1688 15054 1722
rect 15088 1688 15124 1722
rect 15158 1688 15194 1722
rect 15228 1688 15264 1722
rect 15298 1688 15334 1722
rect 15368 1688 15404 1722
rect 15438 1688 15474 1722
rect 15508 1688 15544 1722
rect 15578 1688 15614 1722
rect 15648 1688 15684 1722
rect 15718 1698 15733 1722
rect 15788 1698 15819 1722
rect 15718 1688 15754 1698
rect 15788 1688 15824 1698
rect 15858 1688 15894 1722
rect 15939 1698 15964 1722
rect 16025 1698 16033 1732
rect 15928 1688 15964 1698
rect 15998 1688 16033 1698
rect 14698 1687 16033 1688
rect 13152 1659 16033 1687
rect 13152 1654 15733 1659
rect 15767 1654 15819 1659
rect 15853 1654 15905 1659
rect 15939 1654 15991 1659
rect 13152 1651 14774 1654
rect 344 1575 360 1628
rect 394 1575 410 1628
rect 480 1616 582 1632
rect 3382 1616 3484 1632
rect 12884 1616 12986 1632
rect 13152 1617 13194 1651
rect 13228 1617 13264 1651
rect 13298 1617 13334 1651
rect 13368 1617 13404 1651
rect 13438 1617 13474 1651
rect 13508 1617 13544 1651
rect 13578 1617 13614 1651
rect 13648 1617 13684 1651
rect 13718 1617 13754 1651
rect 13788 1617 13824 1651
rect 13858 1617 13894 1651
rect 13928 1617 13964 1651
rect 13998 1617 14034 1651
rect 14068 1617 14104 1651
rect 14138 1617 14174 1651
rect 14208 1617 14244 1651
rect 14278 1617 14314 1651
rect 14348 1617 14384 1651
rect 14418 1617 14454 1651
rect 14488 1617 14524 1651
rect 14558 1617 14594 1651
rect 14628 1617 14664 1651
rect 14698 1620 14774 1651
rect 14808 1620 14844 1654
rect 14878 1620 14914 1654
rect 14948 1620 14984 1654
rect 15018 1620 15054 1654
rect 15088 1620 15124 1654
rect 15158 1620 15194 1654
rect 15228 1620 15264 1654
rect 15298 1620 15334 1654
rect 15368 1620 15404 1654
rect 15438 1620 15474 1654
rect 15508 1620 15544 1654
rect 15578 1620 15614 1654
rect 15648 1620 15684 1654
rect 15718 1625 15733 1654
rect 15788 1625 15819 1654
rect 15718 1620 15754 1625
rect 15788 1620 15824 1625
rect 15858 1620 15894 1654
rect 15939 1625 15964 1654
rect 16025 1625 16033 1659
rect 15928 1620 15964 1625
rect 15998 1620 16033 1625
rect 14698 1617 16033 1620
rect 514 1582 548 1616
rect 3416 1582 3450 1616
rect 12918 1582 12952 1616
rect 13152 1586 16033 1617
rect 344 1556 410 1575
rect 480 1566 582 1582
rect 3382 1566 3484 1582
rect 12884 1566 12986 1582
rect 13152 1581 14774 1586
rect 344 1505 360 1556
rect 394 1505 410 1556
rect 344 1484 410 1505
rect 344 1435 360 1484
rect 394 1435 410 1484
rect 13152 1547 13194 1581
rect 13228 1547 13264 1581
rect 13298 1547 13334 1581
rect 13368 1547 13404 1581
rect 13438 1547 13474 1581
rect 13508 1547 13544 1581
rect 13578 1547 13614 1581
rect 13648 1547 13684 1581
rect 13718 1547 13754 1581
rect 13788 1547 13824 1581
rect 13858 1547 13894 1581
rect 13928 1547 13964 1581
rect 13998 1547 14034 1581
rect 14068 1547 14104 1581
rect 14138 1547 14174 1581
rect 14208 1547 14244 1581
rect 14278 1547 14314 1581
rect 14348 1547 14384 1581
rect 14418 1547 14454 1581
rect 14488 1547 14524 1581
rect 14558 1547 14594 1581
rect 14628 1547 14664 1581
rect 14698 1552 14774 1581
rect 14808 1552 14844 1586
rect 14878 1552 14914 1586
rect 14948 1552 14984 1586
rect 15018 1552 15054 1586
rect 15088 1552 15124 1586
rect 15158 1552 15194 1586
rect 15228 1552 15264 1586
rect 15298 1552 15334 1586
rect 15368 1552 15404 1586
rect 15438 1552 15474 1586
rect 15508 1552 15544 1586
rect 15578 1552 15614 1586
rect 15648 1552 15684 1586
rect 15718 1552 15733 1586
rect 15788 1552 15819 1586
rect 15858 1552 15894 1586
rect 15939 1552 15964 1586
rect 16025 1552 16033 1586
rect 14698 1547 16033 1552
rect 13152 1518 16033 1547
rect 13152 1511 14774 1518
rect 480 1462 582 1478
rect 3382 1462 3484 1478
rect 12884 1462 12986 1478
rect 13152 1477 13194 1511
rect 13228 1477 13264 1511
rect 13298 1477 13334 1511
rect 13368 1477 13404 1511
rect 13438 1477 13474 1511
rect 13508 1477 13544 1511
rect 13578 1477 13614 1511
rect 13648 1477 13684 1511
rect 13718 1477 13754 1511
rect 13788 1477 13824 1511
rect 13858 1477 13894 1511
rect 13928 1477 13964 1511
rect 13998 1477 14034 1511
rect 14068 1477 14104 1511
rect 14138 1477 14174 1511
rect 14208 1477 14244 1511
rect 14278 1477 14314 1511
rect 14348 1477 14384 1511
rect 14418 1477 14454 1511
rect 14488 1477 14524 1511
rect 14558 1477 14594 1511
rect 14628 1477 14664 1511
rect 14698 1484 14774 1511
rect 14808 1484 14844 1518
rect 14878 1484 14914 1518
rect 14948 1484 14984 1518
rect 15018 1484 15054 1518
rect 15088 1484 15124 1518
rect 15158 1484 15194 1518
rect 15228 1484 15264 1518
rect 15298 1484 15334 1518
rect 15368 1484 15404 1518
rect 15438 1484 15474 1518
rect 15508 1484 15544 1518
rect 15578 1484 15614 1518
rect 15648 1484 15684 1518
rect 15718 1513 15754 1518
rect 15788 1513 15824 1518
rect 15718 1484 15733 1513
rect 15788 1484 15819 1513
rect 15858 1484 15894 1518
rect 15928 1513 15964 1518
rect 15998 1513 16033 1518
rect 15939 1484 15964 1513
rect 14698 1479 15733 1484
rect 15767 1479 15819 1484
rect 15853 1479 15905 1484
rect 15939 1479 15991 1484
rect 16025 1479 16033 1513
rect 14698 1477 16033 1479
rect 344 1412 410 1435
rect 514 1428 548 1462
rect 3416 1428 3450 1462
rect 12918 1428 12952 1462
rect 13152 1450 16033 1477
rect 13152 1441 14774 1450
rect 480 1412 582 1428
rect 3382 1412 3484 1428
rect 12884 1412 12986 1428
rect 344 1365 360 1412
rect 394 1365 410 1412
rect 344 1340 410 1365
rect 344 1295 360 1340
rect 394 1295 410 1340
rect 13152 1407 13194 1441
rect 13228 1407 13264 1441
rect 13298 1407 13334 1441
rect 13368 1407 13404 1441
rect 13438 1407 13474 1441
rect 13508 1407 13544 1441
rect 13578 1407 13614 1441
rect 13648 1407 13684 1441
rect 13718 1407 13754 1441
rect 13788 1407 13824 1441
rect 13858 1407 13894 1441
rect 13928 1407 13964 1441
rect 13998 1407 14034 1441
rect 14068 1407 14104 1441
rect 14138 1407 14174 1441
rect 14208 1407 14244 1441
rect 14278 1407 14314 1441
rect 14348 1407 14384 1441
rect 14418 1407 14454 1441
rect 14488 1407 14524 1441
rect 14558 1407 14594 1441
rect 14628 1407 14664 1441
rect 14698 1416 14774 1441
rect 14808 1416 14844 1450
rect 14878 1416 14914 1450
rect 14948 1416 14984 1450
rect 15018 1416 15054 1450
rect 15088 1416 15124 1450
rect 15158 1416 15194 1450
rect 15228 1416 15264 1450
rect 15298 1416 15334 1450
rect 15368 1416 15404 1450
rect 15438 1416 15474 1450
rect 15508 1416 15544 1450
rect 15578 1416 15614 1450
rect 15648 1416 15684 1450
rect 15718 1440 15754 1450
rect 15788 1440 15824 1450
rect 15718 1416 15733 1440
rect 15788 1416 15819 1440
rect 15858 1416 15894 1450
rect 15928 1440 15964 1450
rect 15998 1440 16033 1450
rect 15939 1416 15964 1440
rect 14698 1407 15733 1416
rect 13152 1406 15733 1407
rect 15767 1406 15819 1416
rect 15853 1406 15905 1416
rect 15939 1406 15991 1416
rect 16025 1406 16033 1440
rect 13152 1385 16033 1406
rect 13152 1351 13168 1385
rect 13202 1371 13244 1385
rect 13278 1371 13320 1385
rect 13354 1371 13396 1385
rect 13430 1371 13472 1385
rect 13506 1371 13548 1385
rect 13582 1371 13624 1385
rect 13658 1371 13700 1385
rect 13734 1371 13776 1385
rect 13810 1371 13851 1385
rect 13885 1371 13926 1385
rect 13960 1371 14001 1385
rect 14035 1371 14076 1385
rect 14110 1371 14151 1385
rect 14185 1371 14226 1385
rect 14260 1371 14301 1385
rect 14335 1371 14376 1385
rect 14410 1371 14451 1385
rect 14485 1371 14526 1385
rect 14560 1371 14601 1385
rect 14635 1382 16033 1385
rect 14635 1371 14774 1382
rect 13228 1351 13244 1371
rect 13298 1351 13320 1371
rect 13368 1351 13396 1371
rect 13438 1351 13472 1371
rect 13152 1337 13194 1351
rect 13228 1337 13264 1351
rect 13298 1337 13334 1351
rect 13368 1337 13404 1351
rect 13438 1337 13474 1351
rect 13508 1337 13544 1371
rect 13582 1351 13614 1371
rect 13658 1351 13684 1371
rect 13734 1351 13754 1371
rect 13810 1351 13824 1371
rect 13885 1351 13894 1371
rect 13960 1351 13964 1371
rect 13578 1337 13614 1351
rect 13648 1337 13684 1351
rect 13718 1337 13754 1351
rect 13788 1337 13824 1351
rect 13858 1337 13894 1351
rect 13928 1337 13964 1351
rect 13998 1351 14001 1371
rect 14068 1351 14076 1371
rect 14138 1351 14151 1371
rect 14208 1351 14226 1371
rect 14278 1351 14301 1371
rect 14348 1351 14376 1371
rect 14418 1351 14451 1371
rect 13998 1337 14034 1351
rect 14068 1337 14104 1351
rect 14138 1337 14174 1351
rect 14208 1337 14244 1351
rect 14278 1337 14314 1351
rect 14348 1337 14384 1351
rect 14418 1337 14454 1351
rect 14488 1337 14524 1371
rect 14560 1351 14594 1371
rect 14635 1351 14664 1371
rect 14558 1337 14594 1351
rect 14628 1337 14664 1351
rect 14698 1348 14774 1371
rect 14808 1348 14844 1382
rect 14878 1348 14914 1382
rect 14948 1348 14984 1382
rect 15018 1348 15054 1382
rect 15088 1348 15124 1382
rect 15158 1348 15194 1382
rect 15228 1348 15264 1382
rect 15298 1348 15334 1382
rect 15368 1348 15404 1382
rect 15438 1348 15474 1382
rect 15508 1348 15544 1382
rect 15578 1348 15614 1382
rect 15648 1348 15684 1382
rect 15718 1367 15754 1382
rect 15788 1367 15824 1382
rect 15718 1348 15733 1367
rect 15788 1348 15819 1367
rect 15858 1348 15894 1382
rect 15928 1367 15964 1382
rect 15998 1367 16033 1382
rect 15939 1348 15964 1367
rect 14698 1337 15733 1348
rect 13152 1333 15733 1337
rect 15767 1333 15819 1348
rect 15853 1333 15905 1348
rect 15939 1333 15991 1348
rect 16025 1333 16033 1367
rect 480 1308 582 1324
rect 3382 1308 3484 1324
rect 12884 1308 12986 1324
rect 13152 1314 16033 1333
rect 344 1268 410 1295
rect 514 1274 548 1308
rect 3416 1274 3450 1308
rect 12918 1274 12952 1308
rect 13152 1301 14774 1314
rect 344 1225 360 1268
rect 394 1225 410 1268
rect 480 1258 582 1274
rect 3382 1258 3484 1274
rect 12884 1258 12986 1274
rect 13152 1267 13194 1301
rect 13228 1267 13264 1301
rect 13298 1267 13334 1301
rect 13368 1267 13404 1301
rect 13438 1267 13474 1301
rect 13508 1267 13544 1301
rect 13578 1267 13614 1301
rect 13648 1267 13684 1301
rect 13718 1267 13754 1301
rect 13788 1267 13824 1301
rect 13858 1267 13894 1301
rect 13928 1267 13964 1301
rect 13998 1267 14034 1301
rect 14068 1267 14104 1301
rect 14138 1267 14174 1301
rect 14208 1267 14244 1301
rect 14278 1267 14314 1301
rect 14348 1267 14384 1301
rect 14418 1267 14454 1301
rect 14488 1267 14524 1301
rect 14558 1267 14594 1301
rect 14628 1267 14664 1301
rect 14698 1280 14774 1301
rect 14808 1280 14844 1314
rect 14878 1280 14914 1314
rect 14948 1280 14984 1314
rect 15018 1280 15054 1314
rect 15088 1280 15124 1314
rect 15158 1280 15194 1314
rect 15228 1280 15264 1314
rect 15298 1280 15334 1314
rect 15368 1280 15404 1314
rect 15438 1280 15474 1314
rect 15508 1280 15544 1314
rect 15578 1280 15614 1314
rect 15648 1280 15684 1314
rect 15718 1294 15754 1314
rect 15788 1294 15824 1314
rect 15718 1280 15733 1294
rect 15788 1280 15819 1294
rect 15858 1280 15894 1314
rect 15928 1294 15964 1314
rect 15998 1294 16033 1314
rect 15939 1280 15964 1294
rect 14698 1267 15733 1280
rect 13152 1260 15733 1267
rect 15767 1260 15819 1280
rect 15853 1260 15905 1280
rect 15939 1260 15991 1280
rect 16025 1260 16033 1294
rect 344 1196 410 1225
rect 344 1155 360 1196
rect 394 1155 410 1196
rect 13152 1246 16033 1260
rect 13152 1231 14774 1246
rect 13152 1197 13194 1231
rect 13228 1197 13264 1231
rect 13298 1197 13334 1231
rect 13368 1197 13404 1231
rect 13438 1197 13474 1231
rect 13508 1197 13544 1231
rect 13578 1197 13614 1231
rect 13648 1197 13684 1231
rect 13718 1197 13754 1231
rect 13788 1197 13824 1231
rect 13858 1197 13894 1231
rect 13928 1197 13964 1231
rect 13998 1197 14034 1231
rect 14068 1197 14104 1231
rect 14138 1197 14174 1231
rect 14208 1197 14244 1231
rect 14278 1197 14314 1231
rect 14348 1197 14384 1231
rect 14418 1197 14454 1231
rect 14488 1197 14524 1231
rect 14558 1197 14594 1231
rect 14628 1197 14664 1231
rect 14698 1212 14774 1231
rect 14808 1212 14844 1246
rect 14878 1212 14914 1246
rect 14948 1212 14984 1246
rect 15018 1212 15054 1246
rect 15088 1212 15124 1246
rect 15158 1212 15194 1246
rect 15228 1212 15264 1246
rect 15298 1212 15334 1246
rect 15368 1212 15404 1246
rect 15438 1212 15474 1246
rect 15508 1212 15544 1246
rect 15578 1212 15614 1246
rect 15648 1212 15684 1246
rect 15718 1221 15754 1246
rect 15788 1221 15824 1246
rect 15718 1212 15733 1221
rect 15788 1212 15819 1221
rect 15858 1212 15894 1246
rect 15928 1221 15964 1246
rect 15998 1221 16033 1246
rect 15939 1212 15964 1221
rect 14698 1197 15733 1212
rect 13152 1187 15733 1197
rect 15767 1187 15819 1212
rect 15853 1187 15905 1212
rect 15939 1187 15991 1212
rect 16025 1187 16033 1221
rect 13152 1178 16033 1187
rect 344 1124 410 1155
rect 480 1154 582 1170
rect 3382 1154 3484 1170
rect 12884 1154 12986 1170
rect 13152 1161 14774 1178
rect 344 1085 360 1124
rect 394 1085 410 1124
rect 514 1120 548 1154
rect 3416 1120 3450 1154
rect 12918 1120 12952 1154
rect 13152 1127 13194 1161
rect 13228 1127 13264 1161
rect 13298 1127 13334 1161
rect 13368 1127 13404 1161
rect 13438 1127 13474 1161
rect 13508 1127 13544 1161
rect 13578 1127 13614 1161
rect 13648 1127 13684 1161
rect 13718 1127 13754 1161
rect 13788 1127 13824 1161
rect 13858 1127 13894 1161
rect 13928 1127 13964 1161
rect 13998 1127 14034 1161
rect 14068 1127 14104 1161
rect 14138 1127 14174 1161
rect 14208 1127 14244 1161
rect 14278 1127 14314 1161
rect 14348 1127 14384 1161
rect 14418 1127 14454 1161
rect 14488 1127 14524 1161
rect 14558 1127 14594 1161
rect 14628 1127 14664 1161
rect 14698 1144 14774 1161
rect 14808 1144 14844 1178
rect 14878 1144 14914 1178
rect 14948 1144 14984 1178
rect 15018 1144 15054 1178
rect 15088 1144 15124 1178
rect 15158 1144 15194 1178
rect 15228 1144 15264 1178
rect 15298 1144 15334 1178
rect 15368 1144 15404 1178
rect 15438 1144 15474 1178
rect 15508 1144 15544 1178
rect 15578 1144 15614 1178
rect 15648 1144 15684 1178
rect 15718 1148 15754 1178
rect 15788 1148 15824 1178
rect 15718 1144 15733 1148
rect 15788 1144 15819 1148
rect 15858 1144 15894 1178
rect 15928 1148 15964 1178
rect 15998 1148 16033 1178
rect 15939 1144 15964 1148
rect 14698 1127 15733 1144
rect 480 1104 582 1120
rect 3382 1104 3484 1120
rect 12884 1104 12986 1120
rect 13152 1114 15733 1127
rect 15767 1114 15819 1144
rect 15853 1114 15905 1144
rect 15939 1114 15991 1144
rect 16025 1114 16033 1148
rect 13152 1110 16033 1114
rect 344 1052 410 1085
rect 344 1016 360 1052
rect 394 1016 410 1052
rect 13152 1091 14774 1110
rect 13152 1077 13194 1091
rect 13228 1077 13264 1091
rect 13298 1077 13334 1091
rect 13368 1077 13404 1091
rect 13438 1077 13474 1091
rect 13152 1043 13168 1077
rect 13228 1057 13244 1077
rect 13298 1057 13320 1077
rect 13368 1057 13396 1077
rect 13438 1057 13472 1077
rect 13508 1057 13544 1091
rect 13578 1077 13614 1091
rect 13648 1077 13684 1091
rect 13718 1077 13754 1091
rect 13788 1077 13824 1091
rect 13858 1077 13894 1091
rect 13928 1077 13964 1091
rect 13582 1057 13614 1077
rect 13658 1057 13684 1077
rect 13734 1057 13754 1077
rect 13810 1057 13824 1077
rect 13885 1057 13894 1077
rect 13960 1057 13964 1077
rect 13998 1077 14034 1091
rect 14068 1077 14104 1091
rect 14138 1077 14174 1091
rect 14208 1077 14244 1091
rect 14278 1077 14314 1091
rect 14348 1077 14384 1091
rect 14418 1077 14454 1091
rect 13998 1057 14001 1077
rect 14068 1057 14076 1077
rect 14138 1057 14151 1077
rect 14208 1057 14226 1077
rect 14278 1057 14301 1077
rect 14348 1057 14376 1077
rect 14418 1057 14451 1077
rect 14488 1057 14524 1091
rect 14558 1077 14594 1091
rect 14628 1077 14664 1091
rect 14560 1057 14594 1077
rect 14635 1057 14664 1077
rect 14698 1076 14774 1091
rect 14808 1076 14844 1110
rect 14878 1076 14914 1110
rect 14948 1076 14984 1110
rect 15018 1076 15054 1110
rect 15088 1076 15124 1110
rect 15158 1076 15194 1110
rect 15228 1076 15264 1110
rect 15298 1076 15334 1110
rect 15368 1076 15404 1110
rect 15438 1076 15474 1110
rect 15508 1076 15544 1110
rect 15578 1076 15614 1110
rect 15648 1076 15684 1110
rect 15718 1076 15754 1110
rect 15788 1076 15824 1110
rect 15858 1076 15894 1110
rect 15928 1076 15964 1110
rect 15998 1076 16033 1110
rect 14698 1075 16033 1076
rect 14698 1057 15733 1075
rect 13202 1043 13244 1057
rect 13278 1043 13320 1057
rect 13354 1043 13396 1057
rect 13430 1043 13472 1057
rect 13506 1043 13548 1057
rect 13582 1043 13624 1057
rect 13658 1043 13700 1057
rect 13734 1043 13776 1057
rect 13810 1043 13851 1057
rect 13885 1043 13926 1057
rect 13960 1043 14001 1057
rect 14035 1043 14076 1057
rect 14110 1043 14151 1057
rect 14185 1043 14226 1057
rect 14260 1043 14301 1057
rect 14335 1043 14376 1057
rect 14410 1043 14451 1057
rect 14485 1043 14526 1057
rect 14560 1043 14601 1057
rect 14635 1043 15733 1057
rect 13152 1042 15733 1043
rect 15767 1042 15819 1075
rect 15853 1042 15905 1075
rect 15939 1042 15991 1075
rect 13152 1021 14774 1042
rect 344 981 410 1016
rect 480 1000 582 1016
rect 3382 1000 3484 1016
rect 12884 1000 12986 1016
rect 344 946 360 981
rect 394 946 410 981
rect 514 966 548 1000
rect 3416 966 3450 1000
rect 12918 966 12952 1000
rect 13152 987 13194 1021
rect 13228 987 13264 1021
rect 13298 987 13334 1021
rect 13368 987 13404 1021
rect 13438 987 13474 1021
rect 13508 987 13544 1021
rect 13578 987 13614 1021
rect 13648 987 13684 1021
rect 13718 987 13754 1021
rect 13788 987 13824 1021
rect 13858 987 13894 1021
rect 13928 987 13964 1021
rect 13998 987 14034 1021
rect 14068 987 14104 1021
rect 14138 987 14174 1021
rect 14208 987 14244 1021
rect 14278 987 14314 1021
rect 14348 987 14384 1021
rect 14418 987 14454 1021
rect 14488 987 14524 1021
rect 14558 987 14594 1021
rect 14628 987 14664 1021
rect 14698 1008 14774 1021
rect 14808 1008 14844 1042
rect 14878 1008 14914 1042
rect 14948 1008 14984 1042
rect 15018 1008 15054 1042
rect 15088 1008 15124 1042
rect 15158 1008 15194 1042
rect 15228 1008 15264 1042
rect 15298 1008 15334 1042
rect 15368 1008 15404 1042
rect 15438 1008 15474 1042
rect 15508 1008 15544 1042
rect 15578 1008 15614 1042
rect 15648 1008 15684 1042
rect 15718 1041 15733 1042
rect 15788 1041 15819 1042
rect 15718 1008 15754 1041
rect 15788 1008 15824 1041
rect 15858 1008 15894 1042
rect 15939 1041 15964 1042
rect 16025 1041 16033 1075
rect 15928 1008 15964 1041
rect 15998 1008 16033 1041
rect 14698 1002 16033 1008
rect 14698 987 15733 1002
rect 13152 974 15733 987
rect 15767 974 15819 1002
rect 15853 974 15905 1002
rect 15939 974 15991 1002
rect 480 950 582 966
rect 3382 950 3484 966
rect 12884 950 12986 966
rect 13152 951 14774 974
rect 344 912 410 946
rect 344 874 360 912
rect 394 874 410 912
rect 344 843 410 874
rect 13152 917 13194 951
rect 13228 917 13264 951
rect 13298 917 13334 951
rect 13368 917 13404 951
rect 13438 917 13474 951
rect 13508 917 13544 951
rect 13578 917 13614 951
rect 13648 917 13684 951
rect 13718 917 13754 951
rect 13788 917 13824 951
rect 13858 917 13894 951
rect 13928 917 13964 951
rect 13998 917 14034 951
rect 14068 917 14104 951
rect 14138 917 14174 951
rect 14208 917 14244 951
rect 14278 917 14314 951
rect 14348 917 14384 951
rect 14418 917 14454 951
rect 14488 917 14524 951
rect 14558 917 14594 951
rect 14628 917 14664 951
rect 14698 940 14774 951
rect 14808 940 14844 974
rect 14878 940 14914 974
rect 14948 940 14984 974
rect 15018 940 15054 974
rect 15088 940 15124 974
rect 15158 940 15194 974
rect 15228 940 15264 974
rect 15298 940 15334 974
rect 15368 940 15404 974
rect 15438 940 15474 974
rect 15508 940 15544 974
rect 15578 940 15614 974
rect 15648 940 15684 974
rect 15718 968 15733 974
rect 15788 968 15819 974
rect 15718 940 15754 968
rect 15788 940 15824 968
rect 15858 940 15894 974
rect 15939 968 15964 974
rect 16025 968 16033 1002
rect 15928 940 15964 968
rect 15998 940 16033 968
rect 14698 929 16033 940
rect 14698 917 15733 929
rect 13152 906 15733 917
rect 15767 906 15819 929
rect 15853 906 15905 929
rect 15939 906 15991 929
rect 13152 881 14774 906
rect 480 846 582 862
rect 3382 846 3484 862
rect 12884 846 12986 862
rect 13152 847 13194 881
rect 13228 847 13264 881
rect 13298 847 13334 881
rect 13368 847 13404 881
rect 13438 847 13474 881
rect 13508 847 13544 881
rect 13578 847 13614 881
rect 13648 847 13684 881
rect 13718 847 13754 881
rect 13788 847 13824 881
rect 13858 847 13894 881
rect 13928 847 13964 881
rect 13998 847 14034 881
rect 14068 847 14104 881
rect 14138 847 14174 881
rect 14208 847 14244 881
rect 14278 847 14314 881
rect 14348 847 14384 881
rect 14418 847 14454 881
rect 14488 847 14524 881
rect 14558 847 14594 881
rect 14628 847 14664 881
rect 14698 872 14774 881
rect 14808 872 14844 906
rect 14878 872 14914 906
rect 14948 872 14984 906
rect 15018 872 15054 906
rect 15088 872 15124 906
rect 15158 872 15194 906
rect 15228 872 15264 906
rect 15298 872 15334 906
rect 15368 872 15404 906
rect 15438 872 15474 906
rect 15508 872 15544 906
rect 15578 872 15614 906
rect 15648 872 15684 906
rect 15718 895 15733 906
rect 15788 895 15819 906
rect 15718 872 15754 895
rect 15788 872 15824 895
rect 15858 872 15894 906
rect 15939 895 15964 906
rect 16025 895 16033 929
rect 15928 872 15964 895
rect 15998 872 16033 895
rect 14698 856 16033 872
rect 14698 847 15733 856
rect 344 802 360 843
rect 394 802 410 843
rect 514 812 548 846
rect 3416 812 3450 846
rect 12918 812 12952 846
rect 13152 838 15733 847
rect 15767 838 15819 856
rect 15853 838 15905 856
rect 15939 838 15991 856
rect 344 774 410 802
rect 480 796 582 812
rect 3382 796 3484 812
rect 12884 796 12986 812
rect 13152 811 14774 838
rect 344 730 360 774
rect 394 730 410 774
rect 344 705 410 730
rect 13152 777 13194 811
rect 13228 777 13264 811
rect 13298 777 13334 811
rect 13368 777 13404 811
rect 13438 777 13474 811
rect 13508 777 13544 811
rect 13578 777 13614 811
rect 13648 777 13684 811
rect 13718 777 13754 811
rect 13788 777 13824 811
rect 13858 777 13894 811
rect 13928 777 13964 811
rect 13998 777 14034 811
rect 14068 777 14104 811
rect 14138 777 14174 811
rect 14208 777 14244 811
rect 14278 777 14314 811
rect 14348 777 14384 811
rect 14418 777 14454 811
rect 14488 777 14524 811
rect 14558 777 14594 811
rect 14628 777 14664 811
rect 14698 804 14774 811
rect 14808 804 14844 838
rect 14878 804 14914 838
rect 14948 804 14984 838
rect 15018 804 15054 838
rect 15088 804 15124 838
rect 15158 804 15194 838
rect 15228 804 15264 838
rect 15298 804 15334 838
rect 15368 804 15404 838
rect 15438 804 15474 838
rect 15508 804 15544 838
rect 15578 804 15614 838
rect 15648 804 15684 838
rect 15718 822 15733 838
rect 15788 822 15819 838
rect 15718 804 15754 822
rect 15788 804 15824 822
rect 15858 804 15894 838
rect 15939 822 15964 838
rect 16025 822 16033 856
rect 15928 804 15964 822
rect 15998 804 16033 822
rect 14698 783 16033 804
rect 14698 777 15733 783
rect 13152 770 15733 777
rect 15767 770 15819 783
rect 15853 770 15905 783
rect 15939 770 15991 783
rect 13152 769 14774 770
rect 13152 735 13168 769
rect 13202 741 13244 769
rect 13278 741 13320 769
rect 13354 741 13396 769
rect 13430 741 13472 769
rect 13506 741 13548 769
rect 13582 741 13624 769
rect 13658 741 13700 769
rect 13734 741 13776 769
rect 13810 741 13851 769
rect 13885 741 13926 769
rect 13960 741 14001 769
rect 14035 741 14076 769
rect 14110 741 14151 769
rect 14185 741 14226 769
rect 14260 741 14301 769
rect 14335 741 14376 769
rect 14410 741 14451 769
rect 14485 741 14526 769
rect 14560 741 14601 769
rect 14635 741 14774 769
rect 13228 735 13244 741
rect 13298 735 13320 741
rect 13368 735 13396 741
rect 13438 735 13472 741
rect 344 658 360 705
rect 394 658 410 705
rect 480 692 582 708
rect 3382 692 3484 708
rect 12884 692 12986 708
rect 13152 707 13194 735
rect 13228 707 13264 735
rect 13298 707 13334 735
rect 13368 707 13404 735
rect 13438 707 13474 735
rect 13508 707 13544 741
rect 13582 735 13614 741
rect 13658 735 13684 741
rect 13734 735 13754 741
rect 13810 735 13824 741
rect 13885 735 13894 741
rect 13960 735 13964 741
rect 13578 707 13614 735
rect 13648 707 13684 735
rect 13718 707 13754 735
rect 13788 707 13824 735
rect 13858 707 13894 735
rect 13928 707 13964 735
rect 13998 735 14001 741
rect 14068 735 14076 741
rect 14138 735 14151 741
rect 14208 735 14226 741
rect 14278 735 14301 741
rect 14348 735 14376 741
rect 14418 735 14451 741
rect 13998 707 14034 735
rect 14068 707 14104 735
rect 14138 707 14174 735
rect 14208 707 14244 735
rect 14278 707 14314 735
rect 14348 707 14384 735
rect 14418 707 14454 735
rect 14488 707 14524 741
rect 14560 735 14594 741
rect 14635 735 14664 741
rect 14558 707 14594 735
rect 14628 707 14664 735
rect 14698 736 14774 741
rect 14808 736 14844 770
rect 14878 736 14914 770
rect 14948 736 14984 770
rect 15018 736 15054 770
rect 15088 736 15124 770
rect 15158 736 15194 770
rect 15228 736 15264 770
rect 15298 736 15334 770
rect 15368 736 15404 770
rect 15438 736 15474 770
rect 15508 736 15544 770
rect 15578 736 15614 770
rect 15648 736 15684 770
rect 15718 749 15733 770
rect 15788 749 15819 770
rect 15718 736 15754 749
rect 15788 736 15824 749
rect 15858 736 15894 770
rect 15939 749 15964 770
rect 16025 749 16033 783
rect 15928 736 15964 749
rect 15998 736 16033 749
rect 14698 710 16033 736
rect 14698 707 15733 710
rect 13152 702 15733 707
rect 15767 702 15819 710
rect 15853 702 15905 710
rect 15939 702 15991 710
rect 514 658 548 692
rect 3416 658 3450 692
rect 12918 658 12952 692
rect 13152 671 14774 702
rect 344 636 410 658
rect 480 642 582 658
rect 3382 642 3484 658
rect 12884 642 12986 658
rect 344 586 360 636
rect 394 586 410 636
rect 344 567 410 586
rect 344 514 360 567
rect 394 514 410 567
rect 13152 637 13194 671
rect 13228 637 13264 671
rect 13298 637 13334 671
rect 13368 637 13404 671
rect 13438 637 13474 671
rect 13508 637 13544 671
rect 13578 637 13614 671
rect 13648 637 13684 671
rect 13718 637 13754 671
rect 13788 637 13824 671
rect 13858 637 13894 671
rect 13928 637 13964 671
rect 13998 637 14034 671
rect 14068 637 14104 671
rect 14138 637 14174 671
rect 14208 637 14244 671
rect 14278 637 14314 671
rect 14348 637 14384 671
rect 14418 637 14454 671
rect 14488 637 14524 671
rect 14558 637 14594 671
rect 14628 637 14664 671
rect 14698 668 14774 671
rect 14808 668 14844 702
rect 14878 668 14914 702
rect 14948 668 14984 702
rect 15018 668 15054 702
rect 15088 668 15124 702
rect 15158 668 15194 702
rect 15228 668 15264 702
rect 15298 668 15334 702
rect 15368 668 15404 702
rect 15438 668 15474 702
rect 15508 668 15544 702
rect 15578 668 15614 702
rect 15648 668 15684 702
rect 15718 676 15733 702
rect 15788 676 15819 702
rect 15718 668 15754 676
rect 15788 668 15824 676
rect 15858 668 15894 702
rect 15939 676 15964 702
rect 16025 676 16033 710
rect 15928 668 15964 676
rect 15998 668 16033 676
rect 14698 637 16033 668
rect 13152 634 15733 637
rect 15767 634 15819 637
rect 15853 634 15905 637
rect 15939 634 15991 637
rect 13152 601 14774 634
rect 13152 567 13194 601
rect 13228 567 13264 601
rect 13298 567 13334 601
rect 13368 567 13404 601
rect 13438 567 13474 601
rect 13508 567 13544 601
rect 13578 567 13614 601
rect 13648 567 13684 601
rect 13718 567 13754 601
rect 13788 567 13824 601
rect 13858 567 13894 601
rect 13928 567 13964 601
rect 13998 567 14034 601
rect 14068 567 14104 601
rect 14138 567 14174 601
rect 14208 567 14244 601
rect 14278 567 14314 601
rect 14348 567 14384 601
rect 14418 567 14454 601
rect 14488 567 14524 601
rect 14558 567 14594 601
rect 14628 567 14664 601
rect 14698 600 14774 601
rect 14808 600 14844 634
rect 14878 600 14914 634
rect 14948 600 14984 634
rect 15018 600 15054 634
rect 15088 600 15124 634
rect 15158 600 15194 634
rect 15228 600 15264 634
rect 15298 600 15334 634
rect 15368 600 15404 634
rect 15438 600 15474 634
rect 15508 600 15544 634
rect 15578 600 15614 634
rect 15648 600 15684 634
rect 15718 603 15733 634
rect 15788 603 15819 634
rect 15718 600 15754 603
rect 15788 600 15824 603
rect 15858 600 15894 634
rect 15939 603 15964 634
rect 16025 603 16033 637
rect 15928 600 15964 603
rect 15998 600 16033 603
rect 14698 567 16033 600
rect 13152 566 16033 567
rect 480 538 582 554
rect 3382 538 3484 554
rect 12884 538 12986 554
rect 344 498 410 514
rect 514 504 548 538
rect 3416 504 3450 538
rect 12918 504 12952 538
rect 13152 532 14774 566
rect 14808 532 14844 566
rect 14878 532 14914 566
rect 14948 532 14984 566
rect 15018 532 15054 566
rect 15088 532 15124 566
rect 15158 532 15194 566
rect 15228 532 15264 566
rect 15298 532 15334 566
rect 15368 532 15404 566
rect 15438 532 15474 566
rect 15508 532 15544 566
rect 15578 532 15614 566
rect 15648 532 15684 566
rect 15718 564 15754 566
rect 15788 564 15824 566
rect 15718 532 15733 564
rect 15788 532 15819 564
rect 15858 532 15894 566
rect 15928 564 15964 566
rect 15998 564 16033 566
rect 15939 532 15964 564
rect 13152 531 15733 532
rect 344 442 360 498
rect 394 442 410 498
rect 480 488 582 504
rect 3382 488 3484 504
rect 12884 488 12986 504
rect 13152 497 13194 531
rect 13228 497 13264 531
rect 13298 497 13334 531
rect 13368 497 13404 531
rect 13438 497 13474 531
rect 13508 497 13544 531
rect 13578 497 13614 531
rect 13648 497 13684 531
rect 13718 497 13754 531
rect 13788 497 13824 531
rect 13858 497 13894 531
rect 13928 497 13964 531
rect 13998 497 14034 531
rect 14068 497 14104 531
rect 14138 497 14174 531
rect 14208 497 14244 531
rect 14278 497 14314 531
rect 14348 497 14384 531
rect 14418 497 14454 531
rect 14488 497 14524 531
rect 14558 497 14594 531
rect 14628 497 14664 531
rect 14698 530 15733 531
rect 15767 530 15819 532
rect 15853 530 15905 532
rect 15939 530 15991 532
rect 16025 530 16033 564
rect 14698 498 16033 530
rect 14698 497 14774 498
rect 344 429 410 442
rect 344 370 360 429
rect 394 370 410 429
rect 13152 464 14774 497
rect 14808 464 14844 498
rect 14878 464 14914 498
rect 14948 464 14984 498
rect 15018 464 15054 498
rect 15088 464 15124 498
rect 15158 464 15194 498
rect 15228 464 15264 498
rect 15298 464 15334 498
rect 15368 464 15404 498
rect 15438 464 15474 498
rect 15508 464 15544 498
rect 15578 464 15614 498
rect 15648 464 15684 498
rect 15718 491 15754 498
rect 15788 491 15824 498
rect 15718 464 15733 491
rect 15788 464 15819 491
rect 15858 464 15894 498
rect 15928 491 15964 498
rect 15998 491 16033 498
rect 15939 464 15964 491
rect 13152 461 15733 464
rect 13152 427 13168 461
rect 13228 427 13241 461
rect 13298 427 13314 461
rect 13368 427 13387 461
rect 13438 427 13460 461
rect 13508 427 13533 461
rect 13578 427 13606 461
rect 13648 427 13679 461
rect 13718 427 13752 461
rect 13788 427 13824 461
rect 13859 427 13894 461
rect 13932 427 13964 461
rect 14005 427 14034 461
rect 14078 427 14104 461
rect 14151 427 14174 461
rect 14224 427 14244 461
rect 14297 427 14314 461
rect 14370 427 14384 461
rect 14443 427 14454 461
rect 14516 427 14524 461
rect 14589 427 14594 461
rect 14662 427 14664 461
rect 14698 427 14701 461
rect 14735 427 14774 461
rect 14808 430 14847 461
rect 14881 430 14920 461
rect 14954 430 14993 461
rect 15027 430 15065 461
rect 15099 430 15137 461
rect 15171 430 15209 461
rect 15243 430 15281 461
rect 15315 430 15353 461
rect 15387 430 15425 461
rect 15459 430 15497 461
rect 15531 430 15569 461
rect 15603 430 15641 461
rect 15675 457 15733 461
rect 15767 457 15819 464
rect 15853 457 15905 464
rect 15939 457 15991 464
rect 16025 457 16033 491
rect 15675 430 16033 457
rect 480 384 582 400
rect 3382 384 3484 400
rect 12884 384 12986 400
rect 13152 396 14774 427
rect 14808 396 14844 430
rect 14881 427 14914 430
rect 14954 427 14984 430
rect 15027 427 15054 430
rect 15099 427 15124 430
rect 15171 427 15194 430
rect 15243 427 15264 430
rect 15315 427 15334 430
rect 15387 427 15404 430
rect 15459 427 15474 430
rect 15531 427 15544 430
rect 15603 427 15614 430
rect 15675 427 15684 430
rect 14878 396 14914 427
rect 14948 396 14984 427
rect 15018 396 15054 427
rect 15088 396 15124 427
rect 15158 396 15194 427
rect 15228 396 15264 427
rect 15298 396 15334 427
rect 15368 396 15404 427
rect 15438 396 15474 427
rect 15508 396 15544 427
rect 15578 396 15614 427
rect 15648 396 15684 427
rect 15718 418 15754 430
rect 15788 418 15824 430
rect 15718 396 15733 418
rect 15788 396 15819 418
rect 15858 396 15894 430
rect 15928 418 15964 430
rect 15998 418 16033 430
rect 15939 396 15964 418
rect 13152 391 15733 396
rect 344 360 410 370
rect 344 298 360 360
rect 394 298 410 360
rect 514 350 548 384
rect 3416 350 3450 384
rect 12918 350 12952 384
rect 13152 357 13194 391
rect 13228 357 13264 391
rect 13298 357 13334 391
rect 13368 357 13404 391
rect 13438 357 13474 391
rect 13508 357 13544 391
rect 13578 357 13614 391
rect 13648 357 13684 391
rect 13718 357 13754 391
rect 13788 357 13824 391
rect 13858 357 13894 391
rect 13928 357 13964 391
rect 13998 357 14034 391
rect 14068 357 14104 391
rect 14138 357 14174 391
rect 14208 357 14244 391
rect 14278 357 14314 391
rect 14348 357 14384 391
rect 14418 357 14454 391
rect 14488 357 14524 391
rect 14558 357 14594 391
rect 14628 357 14664 391
rect 14698 384 15733 391
rect 15767 384 15819 396
rect 15853 384 15905 396
rect 15939 384 15991 396
rect 16025 384 16033 418
rect 14698 362 16033 384
rect 14698 357 14774 362
rect 480 334 582 350
rect 3382 334 3484 350
rect 12884 334 12986 350
rect 344 291 410 298
rect 344 226 360 291
rect 394 226 410 291
rect 13152 328 14774 357
rect 14808 328 14844 362
rect 14878 328 14914 362
rect 14948 328 14984 362
rect 15018 328 15054 362
rect 15088 328 15124 362
rect 15158 328 15194 362
rect 15228 328 15264 362
rect 15298 328 15334 362
rect 15368 328 15404 362
rect 15438 328 15474 362
rect 15508 328 15544 362
rect 15578 328 15614 362
rect 15648 328 15684 362
rect 15718 345 15754 362
rect 15788 345 15824 362
rect 15718 328 15733 345
rect 15788 328 15819 345
rect 15858 328 15894 362
rect 15928 345 15964 362
rect 15998 345 16033 362
rect 15939 328 15964 345
rect 13152 321 15733 328
rect 13152 287 13194 321
rect 13228 287 13264 321
rect 13298 287 13334 321
rect 13368 287 13404 321
rect 13438 287 13474 321
rect 13508 287 13544 321
rect 13578 287 13614 321
rect 13648 287 13684 321
rect 13718 287 13754 321
rect 13788 287 13824 321
rect 13858 287 13894 321
rect 13928 287 13964 321
rect 13998 287 14034 321
rect 14068 287 14104 321
rect 14138 287 14174 321
rect 14208 287 14244 321
rect 14278 287 14314 321
rect 14348 287 14384 321
rect 14418 287 14454 321
rect 14488 287 14524 321
rect 14558 287 14594 321
rect 14628 287 14664 321
rect 14698 311 15733 321
rect 15767 311 15819 328
rect 15853 311 15905 328
rect 15939 311 15991 328
rect 16025 311 16033 345
rect 14698 294 16033 311
rect 14698 287 14774 294
rect 13152 260 14774 287
rect 14808 260 14844 294
rect 14878 260 14914 294
rect 14948 260 14984 294
rect 15018 260 15054 294
rect 15088 260 15124 294
rect 15158 260 15194 294
rect 15228 260 15264 294
rect 15298 260 15334 294
rect 15368 260 15404 294
rect 15438 260 15474 294
rect 15508 260 15544 294
rect 15578 260 15614 294
rect 15648 260 15684 294
rect 15718 272 15754 294
rect 15788 272 15824 294
rect 15718 260 15733 272
rect 15788 260 15819 272
rect 15858 260 15894 294
rect 15928 272 15964 294
rect 15998 272 16033 294
rect 15939 260 15964 272
rect 13152 251 15733 260
rect 480 230 582 246
rect 3382 230 3484 246
rect 12884 230 12986 246
rect 344 222 410 226
rect 344 154 360 222
rect 394 154 410 222
rect 514 196 548 230
rect 3416 196 3450 230
rect 12918 196 12952 230
rect 13152 217 13194 251
rect 13228 217 13264 251
rect 13298 217 13334 251
rect 13368 217 13404 251
rect 13438 217 13474 251
rect 13508 217 13544 251
rect 13578 217 13614 251
rect 13648 217 13684 251
rect 13718 217 13754 251
rect 13788 217 13824 251
rect 13858 217 13894 251
rect 13928 217 13964 251
rect 13998 217 14034 251
rect 14068 217 14104 251
rect 14138 217 14174 251
rect 14208 217 14244 251
rect 14278 217 14314 251
rect 14348 217 14384 251
rect 14418 217 14454 251
rect 14488 217 14524 251
rect 14558 217 14594 251
rect 14628 217 14664 251
rect 14698 238 15733 251
rect 15767 238 15819 260
rect 15853 238 15905 260
rect 15939 238 15991 260
rect 16025 238 16033 272
rect 14698 226 16033 238
rect 14698 217 14774 226
rect 480 180 582 196
rect 3382 180 3484 196
rect 12884 180 12986 196
rect 13152 192 14774 217
rect 14808 192 14844 226
rect 14878 192 14914 226
rect 14948 192 14984 226
rect 15018 192 15054 226
rect 15088 192 15124 226
rect 15158 192 15194 226
rect 15228 192 15264 226
rect 15298 192 15334 226
rect 15368 192 15404 226
rect 15438 192 15474 226
rect 15508 192 15544 226
rect 15578 192 15614 226
rect 15648 192 15684 226
rect 15718 199 15754 226
rect 15788 199 15824 226
rect 15718 192 15733 199
rect 15788 192 15819 199
rect 15858 192 15894 226
rect 15928 199 15964 226
rect 15998 199 16033 226
rect 15939 192 15964 199
rect 13152 181 15733 192
rect 344 153 410 154
rect 344 119 360 153
rect 394 119 410 153
rect 344 100 410 119
rect 13152 147 13194 181
rect 13228 147 13264 181
rect 13298 147 13334 181
rect 13368 147 13404 181
rect 13438 147 13474 181
rect 13508 147 13544 181
rect 13578 147 13614 181
rect 13648 147 13684 181
rect 13718 147 13754 181
rect 13788 147 13824 181
rect 13858 147 13894 181
rect 13928 147 13964 181
rect 13998 147 14034 181
rect 14068 147 14104 181
rect 14138 147 14174 181
rect 14208 147 14244 181
rect 14278 147 14314 181
rect 14348 147 14384 181
rect 14418 147 14454 181
rect 14488 147 14524 181
rect 14558 147 14594 181
rect 14628 147 14664 181
rect 14698 165 15733 181
rect 15767 165 15819 192
rect 15853 165 15905 192
rect 15939 165 15991 192
rect 16025 165 16033 199
rect 14698 158 16033 165
rect 14698 147 14774 158
rect 13152 124 14774 147
rect 14808 124 14844 158
rect 14878 124 14914 158
rect 14948 124 14984 158
rect 15018 124 15054 158
rect 15088 124 15124 158
rect 15158 124 15194 158
rect 15228 124 15264 158
rect 15298 124 15334 158
rect 15368 124 15404 158
rect 15438 124 15474 158
rect 15508 124 15544 158
rect 15578 124 15614 158
rect 15648 124 15684 158
rect 15718 126 15754 158
rect 15788 126 15824 158
rect 15718 124 15733 126
rect 15788 124 15819 126
rect 15858 124 15894 158
rect 15928 126 15964 158
rect 15998 126 16033 158
rect 15939 124 15964 126
rect 13152 100 15733 124
rect 344 92 15733 100
rect 15767 92 15819 124
rect 15853 92 15905 124
rect 15939 92 15991 124
rect 16025 92 16033 126
rect 344 84 16033 92
rect 344 50 360 84
rect 423 50 429 84
rect 495 50 498 84
rect 532 50 533 84
rect 601 50 605 84
rect 670 50 677 84
rect 739 50 774 84
rect 808 50 843 84
rect 877 50 912 84
rect 949 50 981 84
rect 1021 50 1050 84
rect 1093 50 1119 84
rect 1165 50 1188 84
rect 1237 50 1257 84
rect 1309 50 1326 84
rect 1381 50 1395 84
rect 1453 50 1464 84
rect 1525 50 1533 84
rect 1597 50 1602 84
rect 1669 50 1671 84
rect 1705 50 1707 84
rect 1774 50 1779 84
rect 1843 50 1851 84
rect 1912 50 1923 84
rect 1981 50 1995 84
rect 2050 50 2067 84
rect 2119 50 2139 84
rect 2188 50 2211 84
rect 2257 50 2283 84
rect 2326 50 2355 84
rect 2395 50 2427 84
rect 2464 50 2499 84
rect 2533 50 2568 84
rect 2605 50 2637 84
rect 2677 50 2706 84
rect 2749 50 2775 84
rect 2821 50 2844 84
rect 2893 50 2913 84
rect 2965 50 2982 84
rect 3037 50 3051 84
rect 3109 50 3120 84
rect 3181 50 3189 84
rect 3253 50 3258 84
rect 3325 50 3327 84
rect 3361 50 3363 84
rect 3430 50 3435 84
rect 3499 50 3507 84
rect 3568 50 3579 84
rect 3637 50 3651 84
rect 3706 50 3723 84
rect 3775 50 3795 84
rect 3844 50 3867 84
rect 3913 50 3939 84
rect 3982 50 4011 84
rect 4051 50 4083 84
rect 4120 50 4155 84
rect 4189 50 4224 84
rect 4261 50 4293 84
rect 4333 50 4362 84
rect 4405 50 4431 84
rect 4477 50 4500 84
rect 4549 50 4569 84
rect 4621 50 4638 84
rect 4693 50 4707 84
rect 4765 50 4776 84
rect 4837 50 4845 84
rect 4909 50 4914 84
rect 4981 50 4982 84
rect 5016 50 5019 84
rect 5084 50 5091 84
rect 5152 50 5163 84
rect 5220 50 5235 84
rect 5288 50 5307 84
rect 5356 50 5379 84
rect 5424 50 5451 84
rect 5492 50 5523 84
rect 5560 50 5594 84
rect 5629 50 5662 84
rect 5701 50 5730 84
rect 5773 50 5798 84
rect 5845 50 5866 84
rect 5917 50 5934 84
rect 5989 50 6002 84
rect 6061 50 6070 84
rect 6133 50 6138 84
rect 6205 50 6206 84
rect 6240 50 6243 84
rect 6308 50 6315 84
rect 6376 50 6387 84
rect 6444 50 6459 84
rect 6512 50 6531 84
rect 6580 50 6603 84
rect 6648 50 6675 84
rect 6716 50 6747 84
rect 6784 50 6818 84
rect 6853 50 6886 84
rect 6925 50 6954 84
rect 6997 50 7022 84
rect 7069 50 7090 84
rect 7141 50 7158 84
rect 7213 50 7226 84
rect 7285 50 7294 84
rect 7357 50 7362 84
rect 7429 50 7430 84
rect 7464 50 7467 84
rect 7532 50 7539 84
rect 7600 50 7611 84
rect 7668 50 7683 84
rect 7736 50 7755 84
rect 7804 50 7827 84
rect 7872 50 7899 84
rect 7940 50 7971 84
rect 8008 50 8042 84
rect 8077 50 8110 84
rect 8149 50 8178 84
rect 8221 50 8246 84
rect 8293 50 8314 84
rect 8365 50 8382 84
rect 8437 50 8450 84
rect 8509 50 8518 84
rect 8581 50 8586 84
rect 8653 50 8654 84
rect 8688 50 8691 84
rect 8756 50 8763 84
rect 8824 50 8835 84
rect 8892 50 8907 84
rect 8960 50 8979 84
rect 9028 50 9051 84
rect 9096 50 9123 84
rect 9164 50 9195 84
rect 9232 50 9266 84
rect 9301 50 9334 84
rect 9373 50 9402 84
rect 9445 50 9470 84
rect 9517 50 9538 84
rect 9589 50 9606 84
rect 9661 50 9674 84
rect 9733 50 9742 84
rect 9805 50 9810 84
rect 9877 50 9878 84
rect 9912 50 9915 84
rect 9980 50 9987 84
rect 10048 50 10059 84
rect 10116 50 10131 84
rect 10184 50 10203 84
rect 10252 50 10275 84
rect 10320 50 10347 84
rect 10388 50 10419 84
rect 10456 50 10490 84
rect 10525 50 10558 84
rect 10597 50 10626 84
rect 10669 50 10694 84
rect 10741 50 10762 84
rect 10813 50 10830 84
rect 10885 50 10898 84
rect 10957 50 10966 84
rect 11029 50 11034 84
rect 11101 50 11102 84
rect 11136 50 11139 84
rect 11204 50 11211 84
rect 11272 50 11283 84
rect 11340 50 11355 84
rect 11408 50 11427 84
rect 11476 50 11499 84
rect 11544 50 11571 84
rect 11612 50 11643 84
rect 11680 50 11714 84
rect 11749 50 11782 84
rect 11821 50 11850 84
rect 11893 50 11918 84
rect 11965 50 11986 84
rect 12037 50 12054 84
rect 12109 50 12122 84
rect 12181 50 12190 84
rect 12253 50 12258 84
rect 12325 50 12326 84
rect 12360 50 12363 84
rect 12428 50 12435 84
rect 12496 50 12507 84
rect 12564 50 12579 84
rect 12632 50 12651 84
rect 12700 50 12723 84
rect 12768 50 12795 84
rect 12836 50 12867 84
rect 12904 50 12938 84
rect 12973 50 13006 84
rect 13045 50 13074 84
rect 13117 50 13142 84
rect 13189 50 13210 84
rect 13261 50 13278 84
rect 13333 50 13346 84
rect 13405 50 13414 84
rect 13477 50 13482 84
rect 13549 50 13550 84
rect 13584 50 13587 84
rect 13652 50 13659 84
rect 13720 50 13731 84
rect 13788 50 13803 84
rect 13856 50 13875 84
rect 13924 50 13947 84
rect 13992 50 14019 84
rect 14060 50 14091 84
rect 14128 50 14162 84
rect 14197 50 14230 84
rect 14269 50 14298 84
rect 14341 50 14366 84
rect 14400 50 14434 84
rect 14468 50 14502 84
rect 14536 50 14570 84
rect 14604 50 14638 84
rect 14672 50 14706 84
rect 14740 50 14774 84
rect 14808 50 14842 84
rect 14876 50 14910 84
rect 14944 50 14978 84
rect 15012 50 15046 84
rect 15080 50 15114 84
rect 15148 50 15182 84
rect 15216 50 15250 84
rect 15284 50 15318 84
rect 15352 50 15386 84
rect 15420 50 15454 84
rect 15488 50 15522 84
rect 15556 50 15590 84
rect 15624 50 15658 84
rect 15692 50 15726 84
rect 15760 53 15794 84
rect 15828 53 15862 84
rect 15767 50 15794 53
rect 15853 50 15862 53
rect 15896 53 15930 84
rect 15964 53 15998 84
rect 15896 50 15905 53
rect 15964 50 15991 53
rect 16032 50 16033 84
rect 344 34 15733 50
rect 15725 19 15733 34
rect 15767 19 15819 50
rect 15853 19 15905 50
rect 15939 19 15991 50
rect 16025 19 16033 50
rect 15725 -13 16033 19
<< viali >>
rect 360 7984 370 8000
rect 370 7984 394 8000
rect 445 7984 474 8018
rect 474 7984 479 8018
rect 517 7984 543 8018
rect 543 7984 551 8018
rect 589 7984 612 8018
rect 612 7984 623 8018
rect 661 7984 681 8018
rect 681 7984 695 8018
rect 745 7984 750 8018
rect 750 7984 779 8018
rect 876 7984 888 8018
rect 888 7984 910 8018
rect 948 7984 957 8018
rect 957 7984 982 8018
rect 1020 7984 1026 8018
rect 1026 7984 1054 8018
rect 1092 7984 1095 8018
rect 1095 7984 1126 8018
rect 1164 7984 1198 8018
rect 1236 7984 1267 8018
rect 1267 7984 1270 8018
rect 1308 7984 1336 8018
rect 1336 7984 1342 8018
rect 1380 7984 1405 8018
rect 1405 7984 1414 8018
rect 1452 7984 1474 8018
rect 1474 7984 1486 8018
rect 1524 7984 1543 8018
rect 1543 7984 1558 8018
rect 1596 7984 1612 8018
rect 1612 7984 1630 8018
rect 1668 7984 1681 8018
rect 1681 7984 1702 8018
rect 1740 7984 1750 8018
rect 1750 7984 1774 8018
rect 1812 7984 1818 8018
rect 1818 7984 1846 8018
rect 1884 7984 1886 8018
rect 1886 7984 1918 8018
rect 1956 7984 1988 8018
rect 1988 7984 1990 8018
rect 2028 7984 2056 8018
rect 2056 7984 2062 8018
rect 2100 7984 2124 8018
rect 2124 7984 2134 8018
rect 2172 7984 2192 8018
rect 2192 7984 2206 8018
rect 2244 7984 2260 8018
rect 2260 7984 2278 8018
rect 2316 7984 2328 8018
rect 2328 7984 2350 8018
rect 2388 7984 2396 8018
rect 2396 7984 2422 8018
rect 2460 7984 2464 8018
rect 2464 7984 2494 8018
rect 2532 7984 2566 8018
rect 2604 7984 2634 8018
rect 2634 7984 2638 8018
rect 2676 7984 2702 8018
rect 2702 7984 2710 8018
rect 2748 7984 2770 8018
rect 2770 7984 2782 8018
rect 2820 7984 2838 8018
rect 2838 7984 2854 8018
rect 2892 7984 2906 8018
rect 2906 7984 2926 8018
rect 2964 7984 2974 8018
rect 2974 7984 2998 8018
rect 3036 7984 3042 8018
rect 3042 7984 3070 8018
rect 3108 7984 3110 8018
rect 3110 7984 3142 8018
rect 3180 7984 3212 8018
rect 3212 7984 3214 8018
rect 3252 7984 3280 8018
rect 3280 7984 3286 8018
rect 3324 7984 3348 8018
rect 3348 7984 3358 8018
rect 3396 7984 3416 8018
rect 3416 7984 3430 8018
rect 3468 7984 3484 8018
rect 3484 7984 3502 8018
rect 3540 7984 3552 8018
rect 3552 7984 3574 8018
rect 3612 7984 3620 8018
rect 3620 7984 3646 8018
rect 3684 7984 3688 8018
rect 3688 7984 3718 8018
rect 3756 7984 3790 8018
rect 3828 7984 3858 8018
rect 3858 7984 3862 8018
rect 3900 7984 3926 8018
rect 3926 7984 3934 8018
rect 3972 7984 3994 8018
rect 3994 7984 4006 8018
rect 4044 7984 4062 8018
rect 4062 7984 4078 8018
rect 4116 7984 4130 8018
rect 4130 7984 4150 8018
rect 4188 7984 4198 8018
rect 4198 7984 4222 8018
rect 4260 7984 4266 8018
rect 4266 7984 4294 8018
rect 4332 7984 4334 8018
rect 4334 7984 4366 8018
rect 4404 7984 4436 8018
rect 4436 7984 4438 8018
rect 4476 7984 4504 8018
rect 4504 7984 4510 8018
rect 4583 7984 4606 8018
rect 4606 7984 4617 8018
rect 4657 7984 4674 8018
rect 4674 7984 4691 8018
rect 4766 7984 4776 8018
rect 4776 7984 4800 8018
rect 4838 7984 4844 8018
rect 4844 7984 4872 8018
rect 4910 7984 4912 8018
rect 4912 7984 4944 8018
rect 4982 7984 5014 8018
rect 5014 7984 5016 8018
rect 5054 7984 5082 8018
rect 5082 7984 5088 8018
rect 5126 7984 5150 8018
rect 5150 7984 5160 8018
rect 5198 7984 5218 8018
rect 5218 7984 5232 8018
rect 5270 7984 5286 8018
rect 5286 7984 5304 8018
rect 5342 7984 5354 8018
rect 5354 7984 5376 8018
rect 5414 7984 5422 8018
rect 5422 7984 5448 8018
rect 5486 7984 5490 8018
rect 5490 7984 5520 8018
rect 5558 7984 5592 8018
rect 5630 7984 5660 8018
rect 5660 7984 5664 8018
rect 5702 7984 5728 8018
rect 5728 7984 5736 8018
rect 5774 7984 5796 8018
rect 5796 7984 5808 8018
rect 5846 7984 5864 8018
rect 5864 7984 5880 8018
rect 5918 7984 5932 8018
rect 5932 7984 5952 8018
rect 5990 7984 6000 8018
rect 6000 7984 6024 8018
rect 6062 7984 6068 8018
rect 6068 7984 6096 8018
rect 6134 7984 6136 8018
rect 6136 7984 6168 8018
rect 6206 7984 6238 8018
rect 6238 7984 6240 8018
rect 6278 7984 6306 8018
rect 6306 7984 6312 8018
rect 6350 7984 6374 8018
rect 6374 7984 6384 8018
rect 6422 7984 6442 8018
rect 6442 7984 6456 8018
rect 6494 7984 6510 8018
rect 6510 7984 6528 8018
rect 6566 7984 6578 8018
rect 6578 7984 6600 8018
rect 6667 7984 6680 8018
rect 6680 7984 6701 8018
rect 6741 7984 6748 8018
rect 6748 7984 6775 8018
rect 6850 7984 6884 8018
rect 6922 7984 6952 8018
rect 6952 7984 6956 8018
rect 6994 7984 7020 8018
rect 7020 7984 7028 8018
rect 7066 7984 7088 8018
rect 7088 7984 7100 8018
rect 7138 7984 7156 8018
rect 7156 7984 7172 8018
rect 7210 7984 7224 8018
rect 7224 7984 7244 8018
rect 7282 7984 7292 8018
rect 7292 7984 7316 8018
rect 7354 7984 7360 8018
rect 7360 7984 7388 8018
rect 7426 7984 7428 8018
rect 7428 7984 7460 8018
rect 7498 7984 7530 8018
rect 7530 7984 7532 8018
rect 7570 7984 7598 8018
rect 7598 7984 7604 8018
rect 7642 7984 7666 8018
rect 7666 7984 7676 8018
rect 7714 7984 7734 8018
rect 7734 7984 7748 8018
rect 7786 7984 7802 8018
rect 7802 7984 7820 8018
rect 7858 7984 7870 8018
rect 7870 7984 7892 8018
rect 7930 7984 7938 8018
rect 7938 7984 7964 8018
rect 8002 7984 8006 8018
rect 8006 7984 8036 8018
rect 8074 7984 8108 8018
rect 8146 7984 8176 8018
rect 8176 7984 8180 8018
rect 8218 7984 8244 8018
rect 8244 7984 8252 8018
rect 8290 7984 8312 8018
rect 8312 7984 8324 8018
rect 8362 7984 8380 8018
rect 8380 7984 8396 8018
rect 8434 7984 8448 8018
rect 8448 7984 8468 8018
rect 8506 7984 8516 8018
rect 8516 7984 8540 8018
rect 8578 7984 8584 8018
rect 8584 7984 8612 8018
rect 8650 7984 8652 8018
rect 8652 7984 8684 8018
rect 8722 7984 8754 8018
rect 8754 7984 8756 8018
rect 8794 7984 8822 8018
rect 8822 7984 8828 8018
rect 8866 7984 8890 8018
rect 8890 7984 8900 8018
rect 8938 7984 8958 8018
rect 8958 7984 8972 8018
rect 9010 7984 9026 8018
rect 9026 7984 9044 8018
rect 9082 7984 9094 8018
rect 9094 7984 9116 8018
rect 9154 7984 9162 8018
rect 9162 7984 9188 8018
rect 9226 7984 9230 8018
rect 9230 7984 9260 8018
rect 9298 7984 9332 8018
rect 9370 7984 9400 8018
rect 9400 7984 9404 8018
rect 9442 7984 9468 8018
rect 9468 7984 9476 8018
rect 9514 7984 9536 8018
rect 9536 7984 9548 8018
rect 9586 7984 9604 8018
rect 9604 7984 9620 8018
rect 9658 7984 9672 8018
rect 9672 7984 9692 8018
rect 9730 7984 9740 8018
rect 9740 7984 9764 8018
rect 9802 7984 9808 8018
rect 9808 7984 9836 8018
rect 9874 7984 9876 8018
rect 9876 7984 9908 8018
rect 9946 7984 9978 8018
rect 9978 7984 9980 8018
rect 10018 7984 10046 8018
rect 10046 7984 10052 8018
rect 10090 7984 10114 8018
rect 10114 7984 10124 8018
rect 10162 7984 10182 8018
rect 10182 7984 10196 8018
rect 10234 7984 10250 8018
rect 10250 7984 10268 8018
rect 10306 7984 10318 8018
rect 10318 7984 10340 8018
rect 10378 7984 10386 8018
rect 10386 7984 10412 8018
rect 10450 7984 10454 8018
rect 10454 7984 10484 8018
rect 10522 7984 10556 8018
rect 10594 7984 10624 8018
rect 10624 7984 10628 8018
rect 10666 7984 10692 8018
rect 10692 7984 10700 8018
rect 10738 7984 10760 8018
rect 10760 7984 10772 8018
rect 10810 7984 10828 8018
rect 10828 7984 10844 8018
rect 10882 7984 10896 8018
rect 10896 7984 10916 8018
rect 10954 7984 10964 8018
rect 10964 7984 10988 8018
rect 11026 7984 11032 8018
rect 11032 7984 11060 8018
rect 11098 7984 11100 8018
rect 11100 7984 11132 8018
rect 11170 7984 11202 8018
rect 11202 7984 11204 8018
rect 11242 7984 11270 8018
rect 11270 7984 11276 8018
rect 11314 7984 11338 8018
rect 11338 7984 11348 8018
rect 11386 7984 11406 8018
rect 11406 7984 11420 8018
rect 11458 7984 11474 8018
rect 11474 7984 11492 8018
rect 11530 7984 11542 8018
rect 11542 7984 11564 8018
rect 11602 7984 11610 8018
rect 11610 7984 11636 8018
rect 11674 7984 11678 8018
rect 11678 7984 11708 8018
rect 11746 7984 11780 8018
rect 11818 7984 11848 8018
rect 11848 7984 11852 8018
rect 11890 7984 11916 8018
rect 11916 7984 11924 8018
rect 11962 7984 11984 8018
rect 11984 7984 11996 8018
rect 12034 7984 12052 8018
rect 12052 7984 12068 8018
rect 12106 7984 12120 8018
rect 12120 7984 12140 8018
rect 12178 7984 12188 8018
rect 12188 7984 12212 8018
rect 12250 7984 12256 8018
rect 12256 7984 12284 8018
rect 12322 7984 12324 8018
rect 12324 7984 12356 8018
rect 12394 7984 12426 8018
rect 12426 7984 12428 8018
rect 12466 7984 12494 8018
rect 12494 7984 12500 8018
rect 12538 7984 12562 8018
rect 12562 7984 12572 8018
rect 12610 7984 12630 8018
rect 12630 7984 12644 8018
rect 12682 7984 12698 8018
rect 12698 7984 12716 8018
rect 12754 7984 12766 8018
rect 12766 7984 12788 8018
rect 12826 7984 12834 8018
rect 12834 7984 12860 8018
rect 12898 7984 12902 8018
rect 12902 7984 12932 8018
rect 12970 7984 13004 8018
rect 13042 7984 13072 8018
rect 13072 7984 13076 8018
rect 13114 7984 13140 8018
rect 13140 7984 13148 8018
rect 13186 7984 13208 8018
rect 13208 7984 13220 8018
rect 13258 7984 13276 8018
rect 13276 7984 13292 8018
rect 13330 7984 13344 8018
rect 13344 7984 13364 8018
rect 13402 7984 13412 8018
rect 13412 7984 13436 8018
rect 13474 7984 13480 8018
rect 13480 7984 13508 8018
rect 13546 7984 13548 8018
rect 13548 7984 13580 8018
rect 15733 7984 15754 8010
rect 15754 7984 15767 8010
rect 15819 7984 15824 8010
rect 15824 7984 15853 8010
rect 15905 7984 15928 8010
rect 15928 7984 15939 8010
rect 15991 7984 15998 8010
rect 15998 7984 16025 8010
rect 360 7966 394 7984
rect 15733 7976 15767 7984
rect 15819 7976 15853 7984
rect 15905 7976 15939 7984
rect 15991 7976 16025 7984
rect 360 7908 394 7928
rect 360 7894 394 7908
rect 15733 7915 15754 7938
rect 15754 7915 15767 7938
rect 15819 7915 15824 7938
rect 15824 7915 15853 7938
rect 15905 7915 15928 7938
rect 15928 7915 15939 7938
rect 15991 7915 15998 7938
rect 15998 7915 16025 7938
rect 15733 7904 15767 7915
rect 15819 7904 15853 7915
rect 15905 7904 15939 7915
rect 15991 7904 16025 7915
rect 360 7838 394 7856
rect 360 7822 394 7838
rect 478 7839 480 7873
rect 480 7839 512 7873
rect 550 7839 582 7873
rect 582 7839 584 7873
rect 3380 7839 3382 7873
rect 3382 7839 3414 7873
rect 3452 7839 3484 7873
rect 3484 7839 3486 7873
rect 12882 7839 12884 7873
rect 12884 7839 12916 7873
rect 12954 7839 12986 7873
rect 12986 7839 12988 7873
rect 15733 7846 15754 7866
rect 15754 7846 15767 7866
rect 15819 7846 15824 7866
rect 15824 7846 15853 7866
rect 15905 7846 15928 7866
rect 15928 7846 15939 7866
rect 15991 7846 15998 7866
rect 15998 7846 16025 7866
rect 15733 7832 15767 7846
rect 15819 7832 15853 7846
rect 15905 7832 15939 7846
rect 15991 7832 16025 7846
rect 360 7768 394 7784
rect 360 7750 394 7768
rect 15733 7777 15754 7794
rect 15754 7777 15767 7794
rect 15819 7777 15824 7794
rect 15824 7777 15853 7794
rect 15905 7777 15928 7794
rect 15928 7777 15939 7794
rect 15991 7777 15998 7794
rect 15998 7777 16025 7794
rect 15733 7760 15767 7777
rect 15819 7760 15853 7777
rect 15905 7760 15939 7777
rect 15991 7760 16025 7777
rect 360 7698 394 7712
rect 360 7678 394 7698
rect 478 7685 480 7719
rect 480 7685 512 7719
rect 550 7685 582 7719
rect 582 7685 584 7719
rect 3380 7685 3382 7719
rect 3382 7685 3414 7719
rect 3452 7685 3484 7719
rect 3484 7685 3486 7719
rect 12882 7685 12884 7719
rect 12884 7685 12916 7719
rect 12954 7685 12986 7719
rect 12986 7685 12988 7719
rect 15733 7708 15754 7722
rect 15754 7708 15767 7722
rect 15819 7708 15824 7722
rect 15824 7708 15853 7722
rect 15905 7708 15928 7722
rect 15928 7708 15939 7722
rect 15991 7708 15998 7722
rect 15998 7708 16025 7722
rect 15733 7688 15767 7708
rect 15819 7688 15853 7708
rect 15905 7688 15939 7708
rect 15991 7688 16025 7708
rect 360 7628 394 7640
rect 360 7606 394 7628
rect 15733 7639 15754 7650
rect 15754 7639 15767 7650
rect 15819 7639 15824 7650
rect 15824 7639 15853 7650
rect 15905 7639 15928 7650
rect 15928 7639 15939 7650
rect 15991 7639 15998 7650
rect 15998 7639 16025 7650
rect 15733 7616 15767 7639
rect 15819 7616 15853 7639
rect 15905 7616 15939 7639
rect 15991 7616 16025 7639
rect 360 7558 394 7568
rect 360 7534 394 7558
rect 478 7531 480 7565
rect 480 7531 512 7565
rect 550 7531 582 7565
rect 582 7531 584 7565
rect 3380 7531 3382 7565
rect 3382 7531 3414 7565
rect 3452 7531 3484 7565
rect 3484 7531 3486 7565
rect 12882 7531 12884 7565
rect 12884 7531 12916 7565
rect 12954 7531 12986 7565
rect 12986 7531 12988 7565
rect 15733 7570 15754 7578
rect 15754 7570 15767 7578
rect 15819 7570 15824 7578
rect 15824 7570 15853 7578
rect 15905 7570 15928 7578
rect 15928 7570 15939 7578
rect 15991 7570 15998 7578
rect 15998 7570 16025 7578
rect 15733 7544 15767 7570
rect 15819 7544 15853 7570
rect 15905 7544 15939 7570
rect 15991 7544 16025 7570
rect 360 7488 394 7496
rect 360 7462 394 7488
rect 15733 7501 15754 7506
rect 15754 7501 15767 7506
rect 15819 7501 15824 7506
rect 15824 7501 15853 7506
rect 15905 7501 15928 7506
rect 15928 7501 15939 7506
rect 15991 7501 15998 7506
rect 15998 7501 16025 7506
rect 15733 7472 15767 7501
rect 15819 7472 15853 7501
rect 15905 7472 15939 7501
rect 15991 7472 16025 7501
rect 360 7418 394 7424
rect 360 7390 394 7418
rect 478 7377 480 7411
rect 480 7377 512 7411
rect 550 7377 582 7411
rect 582 7377 584 7411
rect 3380 7377 3382 7411
rect 3382 7377 3414 7411
rect 3452 7377 3484 7411
rect 3484 7377 3486 7411
rect 12882 7377 12884 7411
rect 12884 7377 12916 7411
rect 12954 7377 12986 7411
rect 12986 7377 12988 7411
rect 15733 7432 15754 7434
rect 15754 7432 15767 7434
rect 15819 7432 15824 7434
rect 15824 7432 15853 7434
rect 15905 7432 15928 7434
rect 15928 7432 15939 7434
rect 15991 7432 15998 7434
rect 15998 7432 16025 7434
rect 15733 7400 15767 7432
rect 15819 7400 15853 7432
rect 15905 7400 15939 7432
rect 15991 7400 16025 7432
rect 360 7348 394 7352
rect 360 7318 394 7348
rect 360 7278 394 7280
rect 360 7246 394 7278
rect 15733 7328 15767 7362
rect 15819 7328 15853 7362
rect 15905 7328 15939 7362
rect 15991 7328 16025 7362
rect 15733 7259 15767 7290
rect 15819 7259 15853 7290
rect 15905 7259 15939 7290
rect 15991 7259 16025 7290
rect 478 7223 480 7257
rect 480 7223 512 7257
rect 550 7223 582 7257
rect 582 7223 584 7257
rect 3380 7223 3382 7257
rect 3382 7223 3414 7257
rect 3452 7223 3484 7257
rect 3484 7223 3486 7257
rect 12882 7223 12884 7257
rect 12884 7223 12916 7257
rect 12954 7223 12986 7257
rect 12986 7223 12988 7257
rect 360 7174 394 7208
rect 360 7104 394 7136
rect 360 7102 394 7104
rect 15733 7256 15754 7259
rect 15754 7256 15767 7259
rect 15819 7256 15824 7259
rect 15824 7256 15853 7259
rect 15905 7256 15928 7259
rect 15928 7256 15939 7259
rect 15991 7256 15998 7259
rect 15998 7256 16025 7259
rect 15733 7190 15767 7218
rect 15819 7190 15853 7218
rect 15905 7190 15939 7218
rect 15991 7190 16025 7218
rect 15733 7184 15754 7190
rect 15754 7184 15767 7190
rect 15819 7184 15824 7190
rect 15824 7184 15853 7190
rect 15905 7184 15928 7190
rect 15928 7184 15939 7190
rect 15991 7184 15998 7190
rect 15998 7184 16025 7190
rect 15733 7121 15767 7146
rect 15819 7121 15853 7146
rect 15905 7121 15939 7146
rect 15991 7121 16025 7146
rect 478 7069 480 7103
rect 480 7069 512 7103
rect 550 7069 582 7103
rect 582 7069 584 7103
rect 3380 7069 3382 7103
rect 3382 7069 3414 7103
rect 3452 7069 3484 7103
rect 3484 7069 3486 7103
rect 12882 7069 12884 7103
rect 12884 7069 12916 7103
rect 12954 7069 12986 7103
rect 12986 7069 12988 7103
rect 360 7034 394 7064
rect 360 7030 394 7034
rect 15733 7112 15754 7121
rect 15754 7112 15767 7121
rect 15819 7112 15824 7121
rect 15824 7112 15853 7121
rect 15905 7112 15928 7121
rect 15928 7112 15939 7121
rect 15991 7112 15998 7121
rect 15998 7112 16025 7121
rect 360 6965 394 6992
rect 360 6958 394 6965
rect 15733 7052 15767 7074
rect 15819 7052 15853 7074
rect 15905 7052 15939 7074
rect 15991 7052 16025 7074
rect 15733 7040 15754 7052
rect 15754 7040 15767 7052
rect 15819 7040 15824 7052
rect 15824 7040 15853 7052
rect 15905 7040 15928 7052
rect 15928 7040 15939 7052
rect 15991 7040 15998 7052
rect 15998 7040 16025 7052
rect 15733 6983 15767 7002
rect 15819 6983 15853 7002
rect 15905 6983 15939 7002
rect 15991 6983 16025 7002
rect 15733 6968 15754 6983
rect 15754 6968 15767 6983
rect 15819 6968 15824 6983
rect 15824 6968 15853 6983
rect 15905 6968 15928 6983
rect 15928 6968 15939 6983
rect 15991 6968 15998 6983
rect 15998 6968 16025 6983
rect 360 6896 394 6920
rect 360 6886 394 6896
rect 478 6915 480 6949
rect 480 6915 512 6949
rect 550 6915 582 6949
rect 582 6915 584 6949
rect 3380 6915 3382 6949
rect 3382 6915 3414 6949
rect 3452 6915 3484 6949
rect 3484 6915 3486 6949
rect 12882 6915 12884 6949
rect 12884 6915 12916 6949
rect 12954 6915 12986 6949
rect 12986 6915 12988 6949
rect 15733 6914 15767 6930
rect 15819 6914 15853 6930
rect 15905 6914 15939 6930
rect 15991 6914 16025 6930
rect 360 6827 394 6848
rect 360 6814 394 6827
rect 15733 6896 15754 6914
rect 15754 6896 15767 6914
rect 15819 6896 15824 6914
rect 15824 6896 15853 6914
rect 15905 6896 15928 6914
rect 15928 6896 15939 6914
rect 15991 6896 15998 6914
rect 15998 6896 16025 6914
rect 15733 6845 15767 6858
rect 15819 6845 15853 6858
rect 15905 6845 15939 6858
rect 15991 6845 16025 6858
rect 15733 6824 15754 6845
rect 15754 6824 15767 6845
rect 15819 6824 15824 6845
rect 15824 6824 15853 6845
rect 15905 6824 15928 6845
rect 15928 6824 15939 6845
rect 15991 6824 15998 6845
rect 15998 6824 16025 6845
rect 360 6758 394 6776
rect 360 6742 394 6758
rect 478 6761 480 6795
rect 480 6761 512 6795
rect 550 6761 582 6795
rect 582 6761 584 6795
rect 3380 6761 3382 6795
rect 3382 6761 3414 6795
rect 3452 6761 3484 6795
rect 3484 6761 3486 6795
rect 12882 6761 12884 6795
rect 12884 6761 12916 6795
rect 12954 6761 12986 6795
rect 12986 6761 12988 6795
rect 15733 6776 15767 6786
rect 15819 6776 15853 6786
rect 15905 6776 15939 6786
rect 15991 6776 16025 6786
rect 360 6689 394 6704
rect 360 6670 394 6689
rect 15733 6752 15754 6776
rect 15754 6752 15767 6776
rect 15819 6752 15824 6776
rect 15824 6752 15853 6776
rect 15905 6752 15928 6776
rect 15928 6752 15939 6776
rect 15991 6752 15998 6776
rect 15998 6752 16025 6776
rect 15733 6707 15767 6714
rect 15819 6707 15853 6714
rect 15905 6707 15939 6714
rect 15991 6707 16025 6714
rect 15733 6680 15754 6707
rect 15754 6680 15767 6707
rect 15819 6680 15824 6707
rect 15824 6680 15853 6707
rect 15905 6680 15928 6707
rect 15928 6680 15939 6707
rect 15991 6680 15998 6707
rect 15998 6680 16025 6707
rect 360 6620 394 6632
rect 360 6598 394 6620
rect 478 6607 480 6641
rect 480 6607 512 6641
rect 550 6607 582 6641
rect 582 6607 584 6641
rect 3380 6607 3382 6641
rect 3382 6607 3414 6641
rect 3452 6607 3484 6641
rect 3484 6607 3486 6641
rect 12882 6607 12884 6641
rect 12884 6607 12916 6641
rect 12954 6607 12986 6641
rect 12986 6607 12988 6641
rect 15733 6638 15767 6642
rect 15819 6638 15853 6642
rect 15905 6638 15939 6642
rect 15991 6638 16025 6642
rect 15733 6608 15754 6638
rect 15754 6608 15767 6638
rect 15819 6608 15824 6638
rect 15824 6608 15853 6638
rect 15905 6608 15928 6638
rect 15928 6608 15939 6638
rect 15991 6608 15998 6638
rect 15998 6608 16025 6638
rect 360 6551 394 6560
rect 360 6526 394 6551
rect 360 6482 394 6488
rect 360 6454 394 6482
rect 15733 6569 15767 6570
rect 15819 6569 15853 6570
rect 15905 6569 15939 6570
rect 15991 6569 16025 6570
rect 15733 6536 15754 6569
rect 15754 6536 15767 6569
rect 15819 6536 15824 6569
rect 15824 6536 15853 6569
rect 15905 6536 15928 6569
rect 15928 6536 15939 6569
rect 15991 6536 15998 6569
rect 15998 6536 16025 6569
rect 478 6453 480 6487
rect 480 6453 512 6487
rect 550 6453 582 6487
rect 582 6453 584 6487
rect 3380 6453 3382 6487
rect 3382 6453 3414 6487
rect 3452 6453 3484 6487
rect 3484 6453 3486 6487
rect 12882 6453 12884 6487
rect 12884 6453 12916 6487
rect 12954 6453 12986 6487
rect 12986 6453 12988 6487
rect 15733 6466 15754 6498
rect 15754 6466 15767 6498
rect 15819 6466 15824 6498
rect 15824 6466 15853 6498
rect 15905 6466 15928 6498
rect 15928 6466 15939 6498
rect 15991 6466 15998 6498
rect 15998 6466 16025 6498
rect 15733 6464 15767 6466
rect 15819 6464 15853 6466
rect 15905 6464 15939 6466
rect 15991 6464 16025 6466
rect 360 6413 394 6416
rect 360 6382 394 6413
rect 360 6310 394 6344
rect 15733 6397 15754 6426
rect 15754 6397 15767 6426
rect 15819 6397 15824 6426
rect 15824 6397 15853 6426
rect 15905 6397 15928 6426
rect 15928 6397 15939 6426
rect 15991 6397 15998 6426
rect 15998 6397 16025 6426
rect 15733 6392 15767 6397
rect 15819 6392 15853 6397
rect 15905 6392 15939 6397
rect 15991 6392 16025 6397
rect 478 6299 480 6333
rect 480 6299 512 6333
rect 550 6299 582 6333
rect 582 6299 584 6333
rect 3380 6299 3382 6333
rect 3382 6299 3414 6333
rect 3452 6299 3484 6333
rect 3484 6299 3486 6333
rect 12882 6299 12884 6333
rect 12884 6299 12916 6333
rect 12954 6299 12986 6333
rect 12986 6299 12988 6333
rect 15733 6328 15754 6354
rect 15754 6328 15767 6354
rect 15819 6328 15824 6354
rect 15824 6328 15853 6354
rect 15905 6328 15928 6354
rect 15928 6328 15939 6354
rect 15991 6328 15998 6354
rect 15998 6328 16025 6354
rect 15733 6320 15767 6328
rect 15819 6320 15853 6328
rect 15905 6320 15939 6328
rect 15991 6320 16025 6328
rect 360 6240 394 6272
rect 360 6238 394 6240
rect 360 6171 394 6200
rect 360 6166 394 6171
rect 15733 6259 15754 6282
rect 15754 6259 15767 6282
rect 15819 6259 15824 6282
rect 15824 6259 15853 6282
rect 15905 6259 15928 6282
rect 15928 6259 15939 6282
rect 15991 6259 15998 6282
rect 15998 6259 16025 6282
rect 15733 6248 15767 6259
rect 15819 6248 15853 6259
rect 15905 6248 15939 6259
rect 15991 6248 16025 6259
rect 15733 6190 15754 6210
rect 15754 6190 15767 6210
rect 15819 6190 15824 6210
rect 15824 6190 15853 6210
rect 15905 6190 15928 6210
rect 15928 6190 15939 6210
rect 15991 6190 15998 6210
rect 15998 6190 16025 6210
rect 478 6145 480 6179
rect 480 6145 512 6179
rect 550 6145 582 6179
rect 582 6145 584 6179
rect 3380 6145 3382 6179
rect 3382 6145 3414 6179
rect 3452 6145 3484 6179
rect 3484 6145 3486 6179
rect 12882 6145 12884 6179
rect 12884 6145 12916 6179
rect 12954 6145 12986 6179
rect 12986 6145 12988 6179
rect 15733 6176 15767 6190
rect 15819 6176 15853 6190
rect 15905 6176 15939 6190
rect 15991 6176 16025 6190
rect 360 6102 394 6128
rect 360 6094 394 6102
rect 15733 6121 15754 6138
rect 15754 6121 15767 6138
rect 15819 6121 15824 6138
rect 15824 6121 15853 6138
rect 15905 6121 15928 6138
rect 15928 6121 15939 6138
rect 15991 6121 15998 6138
rect 15998 6121 16025 6138
rect 15733 6104 15767 6121
rect 15819 6104 15853 6121
rect 15905 6104 15939 6121
rect 15991 6104 16025 6121
rect 15733 6052 15754 6066
rect 15754 6052 15767 6066
rect 15819 6052 15824 6066
rect 15824 6052 15853 6066
rect 15905 6052 15928 6066
rect 15928 6052 15939 6066
rect 15991 6052 15998 6066
rect 15998 6052 16025 6066
rect 389 5999 394 6033
rect 394 5999 423 6033
rect 461 5999 463 6033
rect 463 5999 495 6033
rect 533 5999 567 6033
rect 605 5999 636 6033
rect 636 5999 639 6033
rect 677 5999 705 6033
rect 705 5999 711 6033
rect 765 5999 774 6032
rect 774 5999 799 6032
rect 837 5999 843 6032
rect 843 5999 871 6032
rect 914 5999 946 6033
rect 946 5999 948 6033
rect 986 5999 1015 6033
rect 1015 5999 1020 6033
rect 1058 5999 1084 6033
rect 1084 5999 1092 6033
rect 1130 5999 1153 6033
rect 1153 5999 1164 6033
rect 1202 5999 1222 6033
rect 1222 5999 1236 6033
rect 1274 5999 1291 6033
rect 1291 5999 1308 6033
rect 1346 5999 1360 6033
rect 1360 5999 1380 6033
rect 1418 5999 1429 6033
rect 1429 5999 1452 6033
rect 1490 5999 1498 6033
rect 1498 5999 1524 6033
rect 1562 5999 1567 6033
rect 1567 5999 1596 6033
rect 1634 5999 1636 6033
rect 1636 5999 1668 6033
rect 1706 5999 1740 6033
rect 1778 5999 1809 6033
rect 1809 5999 1812 6033
rect 1850 5999 1878 6033
rect 1878 5999 1884 6033
rect 1922 5999 1947 6033
rect 1947 5999 1956 6033
rect 1994 5999 2016 6033
rect 2016 5999 2028 6033
rect 2066 5999 2085 6033
rect 2085 5999 2100 6033
rect 2138 5999 2154 6033
rect 2154 5999 2172 6033
rect 2210 5999 2223 6033
rect 2223 5999 2244 6033
rect 2282 5999 2292 6033
rect 2292 5999 2316 6033
rect 2354 5999 2361 6033
rect 2361 5999 2388 6033
rect 2426 5999 2430 6033
rect 2430 5999 2460 6033
rect 2498 5999 2499 6033
rect 2499 5999 2532 6033
rect 2570 5999 2602 6033
rect 2602 5999 2604 6033
rect 2642 5999 2671 6033
rect 2671 5999 2676 6033
rect 2714 5999 2740 6033
rect 2740 5999 2748 6033
rect 2786 5999 2809 6033
rect 2809 5999 2820 6033
rect 2858 5999 2878 6033
rect 2878 5999 2892 6033
rect 2930 5999 2947 6033
rect 2947 5999 2964 6033
rect 3002 5999 3016 6033
rect 3016 5999 3036 6033
rect 3074 5999 3085 6033
rect 3085 5999 3108 6033
rect 3146 5999 3154 6033
rect 3154 5999 3180 6033
rect 3218 5999 3223 6033
rect 3223 5999 3252 6033
rect 3290 5999 3291 6033
rect 3291 5999 3324 6033
rect 3362 5999 3393 6033
rect 3393 5999 3396 6033
rect 3434 5999 3461 6033
rect 3461 5999 3468 6033
rect 3506 5999 3529 6033
rect 3529 5999 3540 6033
rect 3578 5999 3597 6033
rect 3597 5999 3612 6033
rect 3650 5999 3665 6033
rect 3665 5999 3684 6033
rect 3722 5999 3733 6033
rect 3733 5999 3756 6033
rect 3794 5999 3801 6033
rect 3801 5999 3828 6033
rect 3866 5999 3869 6033
rect 3869 5999 3900 6033
rect 3938 5999 3971 6033
rect 3971 5999 3972 6033
rect 4010 5999 4039 6033
rect 4039 5999 4044 6033
rect 4082 5999 4107 6033
rect 4107 5999 4116 6033
rect 4154 5999 4175 6033
rect 4175 5999 4188 6033
rect 4226 5999 4243 6033
rect 4243 5999 4260 6033
rect 4298 5999 4311 6033
rect 4311 5999 4332 6033
rect 4370 5999 4379 6033
rect 4379 5999 4404 6033
rect 4442 5999 4447 6033
rect 4447 5999 4476 6033
rect 4514 5999 4515 6033
rect 4515 5999 4548 6033
rect 4618 5999 4651 6032
rect 4651 5999 4652 6032
rect 4690 5999 4719 6032
rect 4719 5999 4724 6032
rect 4773 5999 4787 6033
rect 4787 5999 4807 6033
rect 4845 5999 4855 6033
rect 4855 5999 4879 6033
rect 4917 5999 4923 6033
rect 4923 5999 4951 6033
rect 4989 5999 4991 6033
rect 4991 5999 5023 6033
rect 5061 5999 5093 6033
rect 5093 5999 5095 6033
rect 5133 5999 5161 6033
rect 5161 5999 5167 6033
rect 5205 5999 5229 6033
rect 5229 5999 5239 6033
rect 5277 5999 5297 6033
rect 5297 5999 5311 6033
rect 5349 5999 5365 6033
rect 5365 5999 5383 6033
rect 5421 5999 5433 6033
rect 5433 5999 5455 6033
rect 5493 5999 5501 6033
rect 5501 5999 5527 6033
rect 5565 5999 5569 6033
rect 5569 5999 5599 6033
rect 5637 5999 5671 6033
rect 5709 5999 5739 6033
rect 5739 5999 5743 6033
rect 5781 5999 5807 6033
rect 5807 5999 5815 6033
rect 5853 5999 5875 6033
rect 5875 5999 5887 6033
rect 6195 5999 6215 6033
rect 6215 5999 6229 6033
rect 6269 5999 6283 6033
rect 6283 5999 6303 6033
rect 6342 5999 6351 6033
rect 6351 5999 6376 6033
rect 6415 5999 6419 6033
rect 6419 5999 6449 6033
rect 6488 5999 6521 6033
rect 6521 5999 6522 6033
rect 6561 5999 6589 6033
rect 6589 5999 6595 6033
rect 6634 5999 6657 6033
rect 6657 5999 6668 6033
rect 6707 5999 6725 6033
rect 6725 5999 6741 6033
rect 6780 5999 6793 6033
rect 6793 5999 6814 6033
rect 7069 5999 7099 6033
rect 7099 5999 7103 6033
rect 7141 5999 7167 6033
rect 7167 5999 7175 6033
rect 7213 5999 7235 6033
rect 7235 5999 7247 6033
rect 7285 5999 7303 6033
rect 7303 5999 7319 6033
rect 7357 5999 7371 6033
rect 7371 5999 7391 6033
rect 7429 5999 7439 6033
rect 7439 5999 7463 6033
rect 7501 5999 7507 6033
rect 7507 5999 7535 6033
rect 7573 5999 7575 6033
rect 7575 5999 7607 6033
rect 7932 5999 7949 6033
rect 7949 5999 7966 6033
rect 8004 5999 8017 6033
rect 8017 5999 8038 6033
rect 8076 5999 8085 6033
rect 8085 5999 8110 6033
rect 8148 5999 8153 6033
rect 8153 5999 8182 6033
rect 8220 5999 8221 6033
rect 8221 5999 8254 6033
rect 8292 5999 8323 6033
rect 8323 5999 8326 6033
rect 8364 5999 8391 6033
rect 8391 5999 8398 6033
rect 8436 5999 8459 6033
rect 8459 5999 8470 6033
rect 8790 5999 8799 6033
rect 8799 5999 8824 6033
rect 8862 5999 8867 6033
rect 8867 5999 8896 6033
rect 8934 5999 8935 6033
rect 8935 5999 8968 6033
rect 9006 5999 9037 6033
rect 9037 5999 9040 6033
rect 9078 5999 9105 6033
rect 9105 5999 9112 6033
rect 9150 5999 9173 6033
rect 9173 5999 9184 6033
rect 9222 5999 9241 6033
rect 9241 5999 9256 6033
rect 9294 5999 9309 6033
rect 9309 5999 9328 6033
rect 9628 5999 9649 6033
rect 9649 5999 9662 6033
rect 9700 5999 9717 6033
rect 9717 5999 9734 6033
rect 9772 5999 9785 6033
rect 9785 5999 9806 6033
rect 9844 5999 9853 6033
rect 9853 5999 9878 6033
rect 9916 5999 9921 6033
rect 9921 5999 9950 6033
rect 9988 5999 9989 6033
rect 9989 5999 10022 6033
rect 10060 5999 10091 6033
rect 10091 5999 10094 6033
rect 10132 5999 10159 6033
rect 10159 5999 10166 6033
rect 10538 5999 10567 6033
rect 10567 5999 10572 6033
rect 10610 5999 10635 6033
rect 10635 5999 10644 6033
rect 10682 5999 10703 6033
rect 10703 5999 10716 6033
rect 10754 5999 10771 6033
rect 10771 5999 10788 6033
rect 10826 5999 10839 6033
rect 10839 5999 10860 6033
rect 10898 5999 10907 6033
rect 10907 5999 10932 6033
rect 10970 5999 10975 6033
rect 10975 5999 11004 6033
rect 11042 5999 11043 6033
rect 11043 5999 11076 6033
rect 11114 5999 11145 6033
rect 11145 5999 11148 6033
rect 11186 5999 11213 6033
rect 11213 5999 11220 6033
rect 11258 5999 11281 6033
rect 11281 5999 11292 6033
rect 11330 5999 11349 6033
rect 11349 5999 11364 6033
rect 11402 5999 11417 6033
rect 11417 5999 11436 6033
rect 11474 5999 11485 6033
rect 11485 5999 11508 6033
rect 11546 5999 11553 6033
rect 11553 5999 11580 6033
rect 11618 5999 11621 6033
rect 11621 5999 11652 6033
rect 11690 5999 11723 6033
rect 11723 5999 11724 6033
rect 11762 5999 11791 6033
rect 11791 5999 11796 6033
rect 11834 5999 11859 6033
rect 11859 5999 11868 6033
rect 11906 5999 11927 6033
rect 11927 5999 11940 6033
rect 11978 5999 11995 6033
rect 11995 5999 12012 6033
rect 12050 5999 12063 6033
rect 12063 5999 12084 6033
rect 12122 5999 12131 6033
rect 12131 5999 12156 6033
rect 12194 5999 12199 6033
rect 12199 5999 12228 6033
rect 12266 5999 12267 6033
rect 12267 5999 12300 6033
rect 12338 5999 12369 6033
rect 12369 5999 12372 6033
rect 12410 5999 12437 6033
rect 12437 5999 12444 6033
rect 12482 5999 12505 6033
rect 12505 5999 12516 6033
rect 12554 5999 12573 6033
rect 12573 5999 12588 6033
rect 12626 5999 12641 6033
rect 12641 5999 12660 6033
rect 12698 5999 12709 6033
rect 12709 5999 12732 6033
rect 12770 5999 12777 6033
rect 12777 5999 12804 6033
rect 12842 5999 12845 6033
rect 12845 5999 12876 6033
rect 12914 5999 12947 6033
rect 12947 5999 12948 6033
rect 12986 5999 13015 6033
rect 13015 5999 13020 6033
rect 13058 5999 13083 6033
rect 13083 5999 13092 6033
rect 13165 5999 13185 6033
rect 13185 5999 13199 6033
rect 13240 5999 13253 6033
rect 13253 5999 13274 6033
rect 13315 5999 13321 6033
rect 13321 5999 13349 6033
rect 13390 5999 13423 6033
rect 13423 5999 13424 6033
rect 13465 5999 13491 6033
rect 13491 5999 13499 6033
rect 13540 5999 13559 6033
rect 13559 5999 13574 6033
rect 13615 5999 13627 6033
rect 13627 5999 13649 6033
rect 13690 5999 13695 6033
rect 13695 5999 13724 6033
rect 13765 5999 13797 6033
rect 13797 5999 13799 6033
rect 13840 5999 13865 6033
rect 13865 5999 13874 6033
rect 13915 5999 13933 6033
rect 13933 5999 13949 6033
rect 13990 5999 14001 6033
rect 14001 5999 14024 6033
rect 14065 5999 14069 6033
rect 14069 5999 14099 6033
rect 14140 5999 14171 6033
rect 14171 5999 14174 6033
rect 14215 5999 14239 6033
rect 14239 5999 14249 6033
rect 14290 5999 14307 6033
rect 14307 5999 14324 6033
rect 14365 5999 14375 6033
rect 14375 5999 14399 6033
rect 14440 5999 14443 6033
rect 14443 5999 14474 6033
rect 14515 5999 14545 6033
rect 14545 5999 14549 6033
rect 765 5998 799 5999
rect 837 5998 871 5999
rect 4618 5998 4652 5999
rect 4690 5998 4724 5999
rect 15733 6032 15767 6052
rect 15819 6032 15853 6052
rect 15905 6032 15939 6052
rect 15991 6032 16025 6052
rect 15733 5983 15754 5994
rect 15754 5983 15767 5994
rect 15819 5983 15824 5994
rect 15824 5983 15853 5994
rect 15905 5983 15928 5994
rect 15928 5983 15939 5994
rect 15991 5983 15998 5994
rect 15998 5983 16025 5994
rect 15733 5960 15767 5983
rect 15819 5960 15853 5983
rect 15905 5960 15939 5983
rect 15991 5960 16025 5983
rect 15733 5914 15754 5922
rect 15754 5914 15767 5922
rect 15819 5914 15824 5922
rect 15824 5914 15853 5922
rect 15905 5914 15928 5922
rect 15928 5914 15939 5922
rect 15991 5914 15998 5922
rect 15998 5914 16025 5922
rect 15733 5888 15767 5914
rect 15819 5888 15853 5914
rect 15905 5888 15939 5914
rect 15991 5888 16025 5914
rect 434 5765 462 5799
rect 462 5765 468 5799
rect 506 5765 530 5799
rect 530 5765 540 5799
rect 578 5765 598 5799
rect 598 5765 612 5799
rect 650 5765 666 5799
rect 666 5765 684 5799
rect 722 5765 734 5799
rect 734 5765 756 5799
rect 794 5765 802 5799
rect 802 5765 828 5799
rect 866 5765 870 5799
rect 870 5765 900 5799
rect 938 5765 972 5799
rect 1010 5765 1040 5799
rect 1040 5765 1044 5799
rect 1082 5765 1108 5799
rect 1108 5765 1116 5799
rect 1154 5765 1176 5799
rect 1176 5765 1188 5799
rect 1226 5765 1244 5799
rect 1244 5765 1260 5799
rect 1298 5765 1312 5799
rect 1312 5765 1332 5799
rect 1370 5765 1380 5799
rect 1380 5765 1404 5799
rect 1442 5765 1448 5799
rect 1448 5765 1476 5799
rect 1514 5765 1516 5799
rect 1516 5765 1548 5799
rect 1586 5765 1618 5799
rect 1618 5765 1620 5799
rect 1658 5765 1686 5799
rect 1686 5765 1692 5799
rect 1730 5765 1754 5799
rect 1754 5765 1764 5799
rect 1802 5765 1822 5799
rect 1822 5765 1836 5799
rect 1874 5765 1890 5799
rect 1890 5765 1908 5799
rect 1946 5765 1958 5799
rect 1958 5765 1980 5799
rect 2018 5765 2026 5799
rect 2026 5765 2052 5799
rect 2090 5765 2094 5799
rect 2094 5765 2124 5799
rect 2162 5765 2196 5799
rect 2234 5765 2264 5799
rect 2264 5765 2268 5799
rect 2306 5765 2332 5799
rect 2332 5765 2340 5799
rect 2378 5765 2400 5799
rect 2400 5765 2412 5799
rect 2450 5765 2468 5799
rect 2468 5765 2484 5799
rect 2522 5765 2536 5799
rect 2536 5765 2556 5799
rect 2594 5765 2604 5799
rect 2604 5765 2628 5799
rect 2666 5765 2672 5799
rect 2672 5765 2700 5799
rect 2738 5765 2740 5799
rect 2740 5765 2772 5799
rect 2810 5765 2842 5799
rect 2842 5765 2844 5799
rect 2882 5765 2910 5799
rect 2910 5765 2916 5799
rect 2954 5765 2978 5799
rect 2978 5765 2988 5799
rect 3026 5765 3046 5799
rect 3046 5765 3060 5799
rect 3098 5765 3114 5799
rect 3114 5765 3132 5799
rect 3170 5765 3182 5799
rect 3182 5765 3204 5799
rect 3242 5765 3250 5799
rect 3250 5765 3276 5799
rect 3314 5765 3318 5799
rect 3318 5765 3348 5799
rect 3386 5765 3420 5799
rect 3458 5765 3488 5799
rect 3488 5765 3492 5799
rect 3530 5765 3556 5799
rect 3556 5765 3564 5799
rect 3602 5765 3624 5799
rect 3624 5765 3636 5799
rect 3674 5765 3692 5799
rect 3692 5765 3708 5799
rect 3746 5765 3760 5799
rect 3760 5765 3780 5799
rect 3818 5765 3828 5799
rect 3828 5765 3852 5799
rect 3890 5765 3896 5799
rect 3896 5765 3924 5799
rect 3962 5765 3964 5799
rect 3964 5765 3996 5799
rect 4034 5765 4066 5799
rect 4066 5765 4068 5799
rect 4106 5765 4134 5799
rect 4134 5765 4140 5799
rect 4178 5765 4202 5799
rect 4202 5765 4212 5799
rect 4250 5765 4270 5799
rect 4270 5765 4284 5799
rect 4322 5765 4338 5799
rect 4338 5765 4356 5799
rect 4394 5765 4406 5799
rect 4406 5765 4428 5799
rect 4466 5765 4474 5799
rect 4474 5765 4500 5799
rect 4538 5765 4542 5799
rect 4542 5765 4572 5799
rect 4610 5765 4644 5799
rect 4682 5765 4712 5799
rect 4712 5765 4716 5799
rect 4754 5765 4780 5799
rect 4780 5765 4788 5799
rect 4826 5765 4848 5799
rect 4848 5765 4860 5799
rect 4898 5765 4916 5799
rect 4916 5765 4932 5799
rect 4970 5765 4984 5799
rect 4984 5765 5004 5799
rect 5042 5765 5052 5799
rect 5052 5765 5076 5799
rect 5114 5765 5120 5799
rect 5120 5765 5148 5799
rect 5186 5765 5188 5799
rect 5188 5765 5220 5799
rect 5258 5765 5290 5799
rect 5290 5765 5292 5799
rect 5330 5765 5358 5799
rect 5358 5765 5364 5799
rect 5402 5765 5426 5799
rect 5426 5765 5436 5799
rect 5474 5765 5494 5799
rect 5494 5765 5508 5799
rect 5546 5765 5562 5799
rect 5562 5765 5580 5799
rect 5618 5765 5630 5799
rect 5630 5765 5652 5799
rect 5690 5765 5698 5799
rect 5698 5765 5724 5799
rect 5763 5765 5766 5799
rect 5766 5765 5797 5799
rect 5836 5765 5868 5799
rect 5868 5765 5870 5799
rect 5909 5765 5936 5799
rect 5936 5765 5943 5799
rect 6195 5765 6208 5799
rect 6208 5765 6229 5799
rect 6269 5765 6276 5799
rect 6276 5765 6303 5799
rect 6342 5765 6344 5799
rect 6344 5765 6376 5799
rect 6415 5765 6446 5799
rect 6446 5765 6449 5799
rect 6488 5765 6514 5799
rect 6514 5765 6522 5799
rect 6561 5765 6582 5799
rect 6582 5765 6595 5799
rect 6634 5765 6650 5799
rect 6650 5765 6668 5799
rect 6707 5765 6718 5799
rect 6718 5765 6741 5799
rect 6780 5765 6786 5799
rect 6786 5765 6814 5799
rect 7069 5765 7092 5799
rect 7092 5765 7103 5799
rect 7141 5765 7160 5799
rect 7160 5765 7175 5799
rect 7213 5765 7228 5799
rect 7228 5765 7247 5799
rect 7285 5765 7296 5799
rect 7296 5765 7319 5799
rect 7357 5765 7364 5799
rect 7364 5765 7391 5799
rect 7429 5765 7432 5799
rect 7432 5765 7463 5799
rect 7501 5765 7534 5799
rect 7534 5765 7535 5799
rect 7573 5765 7602 5799
rect 7602 5765 7607 5799
rect 7932 5765 7942 5799
rect 7942 5765 7966 5799
rect 8004 5765 8010 5799
rect 8010 5765 8038 5799
rect 8076 5765 8078 5799
rect 8078 5765 8110 5799
rect 8148 5765 8181 5799
rect 8181 5765 8182 5799
rect 8220 5765 8250 5799
rect 8250 5765 8254 5799
rect 8292 5765 8319 5799
rect 8319 5765 8326 5799
rect 8364 5765 8388 5799
rect 8388 5765 8398 5799
rect 8436 5765 8457 5799
rect 8457 5765 8470 5799
rect 8790 5765 8802 5799
rect 8802 5765 8824 5799
rect 8862 5765 8871 5799
rect 8871 5765 8896 5799
rect 8934 5765 8940 5799
rect 8940 5765 8968 5799
rect 9006 5765 9009 5799
rect 9009 5765 9040 5799
rect 9078 5765 9112 5799
rect 9150 5765 9181 5799
rect 9181 5765 9184 5799
rect 9222 5765 9250 5799
rect 9250 5765 9256 5799
rect 9294 5765 9319 5799
rect 9319 5765 9328 5799
rect 9628 5765 9630 5799
rect 9630 5765 9662 5799
rect 9700 5765 9733 5799
rect 9733 5765 9734 5799
rect 9772 5765 9802 5799
rect 9802 5765 9806 5799
rect 9844 5765 9871 5799
rect 9871 5765 9878 5799
rect 9916 5765 9940 5799
rect 9940 5765 9950 5799
rect 9988 5765 10009 5799
rect 10009 5765 10022 5799
rect 10060 5765 10078 5799
rect 10078 5765 10094 5799
rect 10132 5765 10147 5799
rect 10147 5765 10166 5799
rect 10487 5765 10492 5799
rect 10492 5765 10521 5799
rect 10559 5765 10561 5799
rect 10561 5765 10593 5799
rect 10631 5765 10665 5799
rect 10703 5765 10734 5799
rect 10734 5765 10737 5799
rect 10775 5765 10803 5799
rect 10803 5765 10809 5799
rect 10847 5765 10872 5799
rect 10872 5765 10881 5799
rect 360 5731 394 5765
rect 360 5690 394 5693
rect 360 5659 394 5690
rect 360 5615 394 5621
rect 360 5587 394 5615
rect 10872 5696 10906 5710
rect 10872 5676 10906 5696
rect 360 5541 394 5549
rect 360 5515 394 5541
rect 360 5467 394 5477
rect 360 5443 394 5467
rect 360 5393 394 5405
rect 360 5371 394 5393
rect 360 5321 394 5333
rect 360 5299 394 5321
rect 360 5251 394 5261
rect 360 5227 394 5251
rect 360 5181 394 5189
rect 360 5155 394 5181
rect 360 5111 394 5117
rect 360 5083 394 5111
rect 360 5041 394 5045
rect 360 5011 394 5041
rect 360 4971 394 4973
rect 360 4939 394 4971
rect 360 4868 394 4901
rect 360 4867 394 4868
rect 360 4799 394 4829
rect 360 4795 394 4799
rect 360 4730 394 4757
rect 360 4723 394 4730
rect 360 4661 394 4685
rect 360 4651 394 4661
rect 360 4592 394 4613
rect 360 4579 394 4592
rect 360 4523 394 4541
rect 360 4507 394 4523
rect 360 4454 394 4469
rect 360 4435 394 4454
rect 360 4385 394 4397
rect 360 4363 394 4385
rect 360 4316 394 4325
rect 360 4291 394 4316
rect 480 5387 514 5411
rect 480 5377 514 5387
rect 480 5319 514 5339
rect 480 5305 514 5319
rect 480 5251 514 5267
rect 480 5233 514 5251
rect 480 5183 514 5195
rect 480 5161 514 5183
rect 480 5115 514 5123
rect 480 5089 514 5115
rect 480 5047 514 5051
rect 480 5017 514 5047
rect 480 4945 514 4979
rect 480 4877 514 4907
rect 480 4873 514 4877
rect 480 4809 514 4835
rect 480 4801 514 4809
rect 480 4741 514 4763
rect 480 4729 514 4741
rect 480 4673 514 4691
rect 480 4657 514 4673
rect 480 4605 514 4619
rect 480 4585 514 4605
rect 480 4537 514 4547
rect 480 4513 514 4537
rect 1336 5387 1370 5411
rect 1336 5377 1370 5387
rect 1336 5319 1370 5339
rect 1336 5305 1370 5319
rect 1336 5251 1370 5267
rect 1336 5233 1370 5251
rect 1336 5183 1370 5195
rect 1336 5161 1370 5183
rect 1336 5115 1370 5123
rect 1336 5089 1370 5115
rect 1336 5047 1370 5051
rect 1336 5017 1370 5047
rect 1336 4945 1370 4979
rect 1336 4877 1370 4907
rect 1336 4873 1370 4877
rect 1336 4809 1370 4835
rect 1336 4801 1370 4809
rect 1336 4741 1370 4763
rect 1336 4729 1370 4741
rect 1336 4673 1370 4691
rect 1336 4657 1370 4673
rect 1336 4605 1370 4619
rect 1336 4585 1370 4605
rect 1336 4537 1370 4547
rect 1336 4513 1370 4537
rect 2192 5387 2226 5411
rect 2192 5377 2226 5387
rect 2192 5319 2226 5339
rect 2192 5305 2226 5319
rect 2192 5251 2226 5267
rect 2192 5233 2226 5251
rect 2192 5183 2226 5195
rect 2192 5161 2226 5183
rect 2192 5115 2226 5123
rect 2192 5089 2226 5115
rect 2192 5047 2226 5051
rect 2192 5017 2226 5047
rect 2192 4945 2226 4979
rect 2192 4877 2226 4907
rect 2192 4873 2226 4877
rect 2192 4809 2226 4835
rect 2192 4801 2226 4809
rect 2192 4741 2226 4763
rect 2192 4729 2226 4741
rect 2192 4673 2226 4691
rect 2192 4657 2226 4673
rect 2192 4605 2226 4619
rect 2192 4585 2226 4605
rect 2192 4537 2226 4547
rect 2192 4513 2226 4537
rect 3048 5387 3082 5411
rect 3048 5377 3082 5387
rect 3048 5319 3082 5339
rect 3048 5305 3082 5319
rect 3048 5251 3082 5267
rect 3048 5233 3082 5251
rect 3048 5183 3082 5195
rect 3048 5161 3082 5183
rect 3048 5115 3082 5123
rect 3048 5089 3082 5115
rect 3048 5047 3082 5051
rect 3048 5017 3082 5047
rect 3048 4945 3082 4979
rect 3048 4877 3082 4907
rect 3048 4873 3082 4877
rect 3048 4809 3082 4835
rect 3048 4801 3082 4809
rect 3048 4741 3082 4763
rect 3048 4729 3082 4741
rect 3048 4673 3082 4691
rect 3048 4657 3082 4673
rect 3048 4605 3082 4619
rect 3048 4585 3082 4605
rect 3048 4537 3082 4547
rect 3048 4513 3082 4537
rect 3904 5387 3938 5411
rect 3904 5377 3938 5387
rect 3904 5319 3938 5339
rect 3904 5305 3938 5319
rect 3904 5251 3938 5267
rect 3904 5233 3938 5251
rect 3904 5183 3938 5195
rect 3904 5161 3938 5183
rect 3904 5115 3938 5123
rect 3904 5089 3938 5115
rect 3904 5047 3938 5051
rect 3904 5017 3938 5047
rect 3904 4945 3938 4979
rect 3904 4877 3938 4907
rect 3904 4873 3938 4877
rect 3904 4809 3938 4835
rect 3904 4801 3938 4809
rect 3904 4741 3938 4763
rect 3904 4729 3938 4741
rect 3904 4673 3938 4691
rect 3904 4657 3938 4673
rect 3904 4605 3938 4619
rect 3904 4585 3938 4605
rect 3904 4537 3938 4547
rect 3904 4513 3938 4537
rect 4760 5387 4794 5411
rect 4760 5377 4794 5387
rect 4760 5319 4794 5339
rect 4760 5305 4794 5319
rect 4760 5251 4794 5267
rect 4760 5233 4794 5251
rect 4760 5183 4794 5195
rect 4760 5161 4794 5183
rect 4760 5115 4794 5123
rect 4760 5089 4794 5115
rect 4760 5047 4794 5051
rect 4760 5017 4794 5047
rect 4760 4945 4794 4979
rect 4760 4877 4794 4907
rect 4760 4873 4794 4877
rect 4760 4809 4794 4835
rect 4760 4801 4794 4809
rect 4760 4741 4794 4763
rect 4760 4729 4794 4741
rect 4760 4673 4794 4691
rect 4760 4657 4794 4673
rect 4760 4605 4794 4619
rect 4760 4585 4794 4605
rect 4760 4537 4794 4547
rect 4760 4513 4794 4537
rect 5616 5387 5650 5411
rect 5616 5377 5650 5387
rect 5616 5319 5650 5339
rect 5616 5305 5650 5319
rect 5616 5251 5650 5267
rect 5616 5233 5650 5251
rect 5616 5183 5650 5195
rect 5616 5161 5650 5183
rect 5616 5115 5650 5123
rect 5616 5089 5650 5115
rect 5616 5047 5650 5051
rect 5616 5017 5650 5047
rect 5616 4945 5650 4979
rect 5616 4877 5650 4907
rect 5616 4873 5650 4877
rect 5616 4809 5650 4835
rect 5616 4801 5650 4809
rect 5616 4741 5650 4763
rect 5616 4729 5650 4741
rect 5616 4673 5650 4691
rect 5616 4657 5650 4673
rect 5616 4605 5650 4619
rect 5616 4585 5650 4605
rect 5616 4537 5650 4547
rect 5616 4513 5650 4537
rect 6472 5387 6506 5411
rect 6472 5377 6506 5387
rect 6472 5319 6506 5339
rect 6472 5305 6506 5319
rect 6472 5251 6506 5267
rect 6472 5233 6506 5251
rect 6472 5183 6506 5195
rect 6472 5161 6506 5183
rect 6472 5115 6506 5123
rect 6472 5089 6506 5115
rect 6472 5047 6506 5051
rect 6472 5017 6506 5047
rect 6472 4945 6506 4979
rect 6472 4877 6506 4907
rect 6472 4873 6506 4877
rect 6472 4809 6506 4835
rect 6472 4801 6506 4809
rect 6472 4741 6506 4763
rect 6472 4729 6506 4741
rect 6472 4673 6506 4691
rect 6472 4657 6506 4673
rect 6472 4605 6506 4619
rect 6472 4585 6506 4605
rect 6472 4537 6506 4547
rect 6472 4513 6506 4537
rect 7328 5387 7362 5411
rect 7328 5377 7362 5387
rect 7328 5319 7362 5339
rect 7328 5305 7362 5319
rect 7328 5251 7362 5267
rect 7328 5233 7362 5251
rect 7328 5183 7362 5195
rect 7328 5161 7362 5183
rect 7328 5115 7362 5123
rect 7328 5089 7362 5115
rect 7328 5047 7362 5051
rect 7328 5017 7362 5047
rect 7328 4945 7362 4979
rect 7328 4877 7362 4907
rect 7328 4873 7362 4877
rect 7328 4809 7362 4835
rect 7328 4801 7362 4809
rect 7328 4741 7362 4763
rect 7328 4729 7362 4741
rect 7328 4673 7362 4691
rect 7328 4657 7362 4673
rect 7328 4605 7362 4619
rect 7328 4585 7362 4605
rect 7328 4537 7362 4547
rect 7328 4513 7362 4537
rect 8184 5387 8218 5411
rect 8184 5377 8218 5387
rect 8184 5319 8218 5339
rect 8184 5305 8218 5319
rect 8184 5251 8218 5267
rect 8184 5233 8218 5251
rect 8184 5183 8218 5195
rect 8184 5161 8218 5183
rect 8184 5115 8218 5123
rect 8184 5089 8218 5115
rect 8184 5047 8218 5051
rect 8184 5017 8218 5047
rect 8184 4945 8218 4979
rect 8184 4877 8218 4907
rect 8184 4873 8218 4877
rect 8184 4809 8218 4835
rect 8184 4801 8218 4809
rect 8184 4741 8218 4763
rect 8184 4729 8218 4741
rect 8184 4673 8218 4691
rect 8184 4657 8218 4673
rect 8184 4605 8218 4619
rect 8184 4585 8218 4605
rect 8184 4537 8218 4547
rect 8184 4513 8218 4537
rect 9040 5387 9074 5411
rect 9040 5377 9074 5387
rect 9040 5319 9074 5339
rect 9040 5305 9074 5319
rect 9040 5251 9074 5267
rect 9040 5233 9074 5251
rect 9040 5183 9074 5195
rect 9040 5161 9074 5183
rect 9040 5115 9074 5123
rect 9040 5089 9074 5115
rect 9040 5047 9074 5051
rect 9040 5017 9074 5047
rect 9040 4945 9074 4979
rect 9040 4877 9074 4907
rect 9040 4873 9074 4877
rect 9040 4809 9074 4835
rect 9040 4801 9074 4809
rect 9040 4741 9074 4763
rect 9040 4729 9074 4741
rect 9040 4673 9074 4691
rect 9040 4657 9074 4673
rect 9040 4605 9074 4619
rect 9040 4585 9074 4605
rect 9040 4537 9074 4547
rect 9040 4513 9074 4537
rect 9896 5387 9930 5411
rect 9896 5377 9930 5387
rect 9896 5319 9930 5339
rect 9896 5305 9930 5319
rect 9896 5251 9930 5267
rect 9896 5233 9930 5251
rect 9896 5183 9930 5195
rect 9896 5161 9930 5183
rect 9896 5115 9930 5123
rect 9896 5089 9930 5115
rect 9896 5047 9930 5051
rect 9896 5017 9930 5047
rect 9896 4945 9930 4979
rect 9896 4877 9930 4907
rect 9896 4873 9930 4877
rect 9896 4809 9930 4835
rect 9896 4801 9930 4809
rect 9896 4741 9930 4763
rect 9896 4729 9930 4741
rect 9896 4673 9930 4691
rect 9896 4657 9930 4673
rect 9896 4605 9930 4619
rect 9896 4585 9930 4605
rect 9896 4537 9930 4547
rect 9896 4513 9930 4537
rect 10752 5387 10786 5411
rect 10752 5377 10786 5387
rect 10752 5319 10786 5339
rect 10752 5305 10786 5319
rect 10752 5251 10786 5267
rect 10752 5233 10786 5251
rect 10752 5183 10786 5195
rect 10752 5161 10786 5183
rect 10752 5115 10786 5123
rect 10752 5089 10786 5115
rect 10752 5047 10786 5051
rect 10752 5017 10786 5047
rect 10752 4945 10786 4979
rect 10752 4877 10786 4907
rect 10752 4873 10786 4877
rect 10752 4809 10786 4835
rect 10752 4801 10786 4809
rect 10752 4741 10786 4763
rect 10752 4729 10786 4741
rect 10752 4673 10786 4691
rect 10752 4657 10786 4673
rect 10752 4605 10786 4619
rect 10752 4585 10786 4605
rect 10752 4537 10786 4547
rect 10752 4513 10786 4537
rect 10872 5627 10906 5638
rect 10872 5604 10906 5627
rect 10872 5558 10906 5566
rect 10872 5532 10906 5558
rect 10872 5489 10906 5494
rect 10872 5460 10906 5489
rect 10872 5420 10906 5422
rect 10872 5388 10906 5420
rect 10872 5316 10906 5350
rect 10872 5247 10906 5278
rect 10872 5244 10906 5247
rect 10872 5178 10906 5206
rect 10872 5172 10906 5178
rect 10872 5109 10906 5134
rect 10872 5100 10906 5109
rect 10872 5040 10906 5062
rect 10872 5028 10906 5040
rect 10872 4971 10906 4990
rect 10872 4956 10906 4971
rect 10872 4902 10906 4918
rect 10872 4884 10906 4902
rect 10872 4833 10906 4846
rect 10872 4812 10906 4833
rect 10872 4764 10906 4774
rect 10872 4740 10906 4764
rect 10872 4695 10906 4702
rect 10872 4668 10906 4695
rect 10872 4626 10906 4630
rect 10872 4596 10906 4626
rect 10872 4557 10906 4558
rect 10872 4524 10906 4557
rect 10872 4454 10906 4486
rect 10872 4452 10906 4454
rect 10872 4385 10906 4414
rect 10872 4380 10906 4385
rect 10872 4316 10906 4342
rect 10872 4308 10906 4316
rect 360 4247 394 4253
rect 360 4219 394 4247
rect 552 4205 568 4239
rect 568 4205 586 4239
rect 632 4205 636 4239
rect 636 4205 666 4239
rect 711 4205 738 4239
rect 738 4205 745 4239
rect 790 4205 806 4239
rect 806 4205 824 4239
rect 869 4205 874 4239
rect 874 4205 903 4239
rect 948 4205 976 4239
rect 976 4205 982 4239
rect 1027 4205 1044 4239
rect 1044 4205 1061 4239
rect 1106 4205 1112 4239
rect 1112 4205 1140 4239
rect 1185 4205 1214 4239
rect 1214 4205 1219 4239
rect 1264 4205 1282 4239
rect 1282 4205 1298 4239
rect 1408 4205 1424 4239
rect 1424 4205 1442 4239
rect 1488 4205 1492 4239
rect 1492 4205 1522 4239
rect 1567 4205 1594 4239
rect 1594 4205 1601 4239
rect 1646 4205 1662 4239
rect 1662 4205 1680 4239
rect 1725 4205 1730 4239
rect 1730 4205 1759 4239
rect 1804 4205 1832 4239
rect 1832 4205 1838 4239
rect 1883 4205 1900 4239
rect 1900 4205 1917 4239
rect 1962 4205 1968 4239
rect 1968 4205 1996 4239
rect 2041 4205 2070 4239
rect 2070 4205 2075 4239
rect 2120 4205 2138 4239
rect 2138 4205 2154 4239
rect 2264 4205 2280 4239
rect 2280 4205 2298 4239
rect 2344 4205 2348 4239
rect 2348 4205 2378 4239
rect 2423 4205 2450 4239
rect 2450 4205 2457 4239
rect 2502 4205 2518 4239
rect 2518 4205 2536 4239
rect 2581 4205 2586 4239
rect 2586 4205 2615 4239
rect 2660 4205 2688 4239
rect 2688 4205 2694 4239
rect 2739 4205 2756 4239
rect 2756 4205 2773 4239
rect 2818 4205 2824 4239
rect 2824 4205 2852 4239
rect 2897 4205 2926 4239
rect 2926 4205 2931 4239
rect 2976 4205 2994 4239
rect 2994 4205 3010 4239
rect 3120 4205 3136 4239
rect 3136 4205 3154 4239
rect 3200 4205 3204 4239
rect 3204 4205 3234 4239
rect 3279 4205 3306 4239
rect 3306 4205 3313 4239
rect 3358 4205 3374 4239
rect 3374 4205 3392 4239
rect 3437 4205 3442 4239
rect 3442 4205 3471 4239
rect 3516 4205 3544 4239
rect 3544 4205 3550 4239
rect 3595 4205 3612 4239
rect 3612 4205 3629 4239
rect 3674 4205 3680 4239
rect 3680 4205 3708 4239
rect 3753 4205 3782 4239
rect 3782 4205 3787 4239
rect 3832 4205 3850 4239
rect 3850 4205 3866 4239
rect 3976 4205 3992 4239
rect 3992 4205 4010 4239
rect 4056 4205 4060 4239
rect 4060 4205 4090 4239
rect 4135 4205 4162 4239
rect 4162 4205 4169 4239
rect 4214 4205 4230 4239
rect 4230 4205 4248 4239
rect 4293 4205 4298 4239
rect 4298 4205 4327 4239
rect 4372 4205 4400 4239
rect 4400 4205 4406 4239
rect 4451 4205 4468 4239
rect 4468 4205 4485 4239
rect 4530 4205 4536 4239
rect 4536 4205 4564 4239
rect 4609 4205 4638 4239
rect 4638 4205 4643 4239
rect 4688 4205 4706 4239
rect 4706 4205 4722 4239
rect 4832 4205 4848 4239
rect 4848 4205 4866 4239
rect 4912 4205 4916 4239
rect 4916 4205 4946 4239
rect 4991 4205 5018 4239
rect 5018 4205 5025 4239
rect 5070 4205 5086 4239
rect 5086 4205 5104 4239
rect 5149 4205 5154 4239
rect 5154 4205 5183 4239
rect 5228 4205 5256 4239
rect 5256 4205 5262 4239
rect 5307 4205 5324 4239
rect 5324 4205 5341 4239
rect 5386 4205 5392 4239
rect 5392 4205 5420 4239
rect 5465 4205 5494 4239
rect 5494 4205 5499 4239
rect 5544 4205 5562 4239
rect 5562 4205 5578 4239
rect 5688 4205 5704 4239
rect 5704 4205 5722 4239
rect 5768 4205 5772 4239
rect 5772 4205 5802 4239
rect 5847 4205 5874 4239
rect 5874 4205 5881 4239
rect 5926 4205 5942 4239
rect 5942 4205 5960 4239
rect 6005 4205 6010 4239
rect 6010 4205 6039 4239
rect 6084 4205 6112 4239
rect 6112 4205 6118 4239
rect 6163 4205 6180 4239
rect 6180 4205 6197 4239
rect 6242 4205 6248 4239
rect 6248 4205 6276 4239
rect 6321 4205 6350 4239
rect 6350 4205 6355 4239
rect 6400 4205 6418 4239
rect 6418 4205 6434 4239
rect 6544 4205 6560 4239
rect 6560 4205 6578 4239
rect 6624 4205 6628 4239
rect 6628 4205 6658 4239
rect 6703 4205 6730 4239
rect 6730 4205 6737 4239
rect 6782 4205 6798 4239
rect 6798 4205 6816 4239
rect 6861 4205 6866 4239
rect 6866 4205 6895 4239
rect 6940 4205 6968 4239
rect 6968 4205 6974 4239
rect 7019 4205 7036 4239
rect 7036 4205 7053 4239
rect 7098 4205 7104 4239
rect 7104 4205 7132 4239
rect 7177 4205 7206 4239
rect 7206 4205 7211 4239
rect 7256 4205 7274 4239
rect 7274 4205 7290 4239
rect 7400 4205 7416 4239
rect 7416 4205 7434 4239
rect 7480 4205 7484 4239
rect 7484 4205 7514 4239
rect 7559 4205 7586 4239
rect 7586 4205 7593 4239
rect 7638 4205 7654 4239
rect 7654 4205 7672 4239
rect 7717 4205 7722 4239
rect 7722 4205 7751 4239
rect 7796 4205 7824 4239
rect 7824 4205 7830 4239
rect 7875 4205 7892 4239
rect 7892 4205 7909 4239
rect 7954 4205 7960 4239
rect 7960 4205 7988 4239
rect 8033 4205 8062 4239
rect 8062 4205 8067 4239
rect 8112 4205 8130 4239
rect 8130 4205 8146 4239
rect 8256 4205 8272 4239
rect 8272 4205 8290 4239
rect 8336 4205 8340 4239
rect 8340 4205 8370 4239
rect 8415 4205 8442 4239
rect 8442 4205 8449 4239
rect 8494 4205 8510 4239
rect 8510 4205 8528 4239
rect 8573 4205 8578 4239
rect 8578 4205 8607 4239
rect 8652 4205 8680 4239
rect 8680 4205 8686 4239
rect 8731 4205 8748 4239
rect 8748 4205 8765 4239
rect 8810 4205 8816 4239
rect 8816 4205 8844 4239
rect 8889 4205 8918 4239
rect 8918 4205 8923 4239
rect 8968 4205 8986 4239
rect 8986 4205 9002 4239
rect 9112 4205 9128 4239
rect 9128 4205 9146 4239
rect 9192 4205 9196 4239
rect 9196 4205 9226 4239
rect 9271 4205 9298 4239
rect 9298 4205 9305 4239
rect 9350 4205 9366 4239
rect 9366 4205 9384 4239
rect 9429 4205 9434 4239
rect 9434 4205 9463 4239
rect 9508 4205 9536 4239
rect 9536 4205 9542 4239
rect 9587 4205 9604 4239
rect 9604 4205 9621 4239
rect 9666 4205 9672 4239
rect 9672 4205 9700 4239
rect 9745 4205 9774 4239
rect 9774 4205 9779 4239
rect 9824 4205 9842 4239
rect 9842 4205 9858 4239
rect 9968 4205 9984 4239
rect 9984 4205 10002 4239
rect 10048 4205 10052 4239
rect 10052 4205 10082 4239
rect 10127 4205 10154 4239
rect 10154 4205 10161 4239
rect 10206 4205 10222 4239
rect 10222 4205 10240 4239
rect 10285 4205 10290 4239
rect 10290 4205 10319 4239
rect 10364 4205 10392 4239
rect 10392 4205 10398 4239
rect 10443 4205 10460 4239
rect 10460 4205 10477 4239
rect 10522 4205 10528 4239
rect 10528 4205 10556 4239
rect 10601 4205 10630 4239
rect 10630 4205 10635 4239
rect 10680 4205 10698 4239
rect 10698 4205 10714 4239
rect 10872 4247 10906 4270
rect 10872 4236 10906 4247
rect 379 4109 394 4139
rect 394 4109 413 4139
rect 452 4109 463 4139
rect 463 4109 486 4139
rect 525 4109 532 4139
rect 532 4109 559 4139
rect 598 4109 601 4139
rect 601 4109 632 4139
rect 379 4105 413 4109
rect 452 4105 486 4109
rect 525 4105 559 4109
rect 598 4105 632 4109
rect 671 4105 705 4139
rect 744 4109 774 4139
rect 774 4109 778 4139
rect 817 4109 843 4139
rect 843 4109 851 4139
rect 890 4109 912 4139
rect 912 4109 924 4139
rect 963 4109 981 4139
rect 981 4109 997 4139
rect 1036 4109 1050 4139
rect 1050 4109 1070 4139
rect 1109 4109 1119 4139
rect 1119 4109 1143 4139
rect 1182 4109 1188 4139
rect 1188 4109 1216 4139
rect 1255 4109 1257 4139
rect 1257 4109 1289 4139
rect 1328 4109 1360 4139
rect 1360 4109 1362 4139
rect 1401 4109 1429 4139
rect 1429 4109 1435 4139
rect 1474 4109 1498 4139
rect 1498 4109 1508 4139
rect 1547 4109 1567 4139
rect 1567 4109 1581 4139
rect 1620 4109 1636 4139
rect 1636 4109 1654 4139
rect 1693 4109 1705 4139
rect 1705 4109 1727 4139
rect 1766 4109 1774 4139
rect 1774 4109 1800 4139
rect 1839 4109 1843 4139
rect 1843 4109 1873 4139
rect 744 4105 778 4109
rect 817 4105 851 4109
rect 890 4105 924 4109
rect 963 4105 997 4109
rect 1036 4105 1070 4109
rect 1109 4105 1143 4109
rect 1182 4105 1216 4109
rect 1255 4105 1289 4109
rect 1328 4105 1362 4109
rect 1401 4105 1435 4109
rect 1474 4105 1508 4109
rect 1547 4105 1581 4109
rect 1620 4105 1654 4109
rect 1693 4105 1727 4109
rect 1766 4105 1800 4109
rect 1839 4105 1873 4109
rect 1912 4105 1946 4139
rect 1985 4109 2016 4139
rect 2016 4109 2019 4139
rect 2058 4109 2085 4139
rect 2085 4109 2092 4139
rect 2131 4109 2154 4139
rect 2154 4109 2165 4139
rect 2204 4109 2223 4139
rect 2223 4109 2238 4139
rect 2277 4109 2292 4139
rect 2292 4109 2311 4139
rect 2350 4109 2361 4139
rect 2361 4109 2384 4139
rect 2423 4109 2430 4139
rect 2430 4109 2457 4139
rect 2496 4109 2499 4139
rect 2499 4109 2530 4139
rect 2569 4109 2602 4139
rect 2602 4109 2603 4139
rect 2642 4109 2671 4139
rect 2671 4109 2676 4139
rect 2715 4109 2740 4139
rect 2740 4109 2749 4139
rect 2788 4109 2809 4139
rect 2809 4109 2822 4139
rect 2861 4109 2878 4139
rect 2878 4109 2895 4139
rect 2934 4109 2947 4139
rect 2947 4109 2968 4139
rect 3007 4109 3016 4139
rect 3016 4109 3041 4139
rect 3080 4109 3085 4139
rect 3085 4109 3114 4139
rect 3153 4109 3154 4139
rect 3154 4109 3187 4139
rect 3226 4109 3256 4139
rect 3256 4109 3260 4139
rect 3299 4109 3324 4139
rect 3324 4109 3333 4139
rect 3372 4109 3392 4139
rect 3392 4109 3406 4139
rect 3444 4109 3460 4139
rect 3460 4109 3478 4139
rect 3516 4109 3528 4139
rect 3528 4109 3550 4139
rect 3588 4109 3596 4139
rect 3596 4109 3622 4139
rect 3660 4109 3664 4139
rect 3664 4109 3694 4139
rect 3732 4109 3766 4139
rect 3804 4109 3834 4139
rect 3834 4109 3838 4139
rect 3876 4109 3902 4139
rect 3902 4109 3910 4139
rect 3948 4109 3970 4139
rect 3970 4109 3982 4139
rect 4020 4109 4038 4139
rect 4038 4109 4054 4139
rect 4092 4109 4106 4139
rect 4106 4109 4126 4139
rect 4164 4109 4174 4139
rect 4174 4109 4198 4139
rect 4236 4109 4242 4139
rect 4242 4109 4270 4139
rect 4308 4109 4310 4139
rect 4310 4109 4342 4139
rect 4380 4109 4412 4139
rect 4412 4109 4414 4139
rect 4452 4109 4480 4139
rect 4480 4109 4486 4139
rect 4524 4109 4548 4139
rect 4548 4109 4558 4139
rect 4596 4109 4616 4139
rect 4616 4109 4630 4139
rect 4668 4109 4684 4139
rect 4684 4109 4702 4139
rect 4740 4109 4752 4139
rect 4752 4109 4774 4139
rect 4812 4109 4820 4139
rect 4820 4109 4846 4139
rect 4884 4109 4888 4139
rect 4888 4109 4918 4139
rect 4956 4109 4990 4139
rect 5028 4109 5058 4139
rect 5058 4109 5062 4139
rect 5100 4109 5126 4139
rect 5126 4109 5134 4139
rect 5172 4109 5194 4139
rect 5194 4109 5206 4139
rect 5244 4109 5262 4139
rect 5262 4109 5278 4139
rect 5316 4109 5330 4139
rect 5330 4109 5350 4139
rect 5388 4109 5398 4139
rect 5398 4109 5422 4139
rect 5460 4109 5466 4139
rect 5466 4109 5494 4139
rect 5532 4109 5534 4139
rect 5534 4109 5566 4139
rect 5604 4109 5636 4139
rect 5636 4109 5638 4139
rect 5676 4109 5704 4139
rect 5704 4109 5710 4139
rect 5748 4109 5772 4139
rect 5772 4109 5782 4139
rect 5820 4109 5840 4139
rect 5840 4109 5854 4139
rect 5892 4109 5908 4139
rect 5908 4109 5926 4139
rect 5964 4109 5976 4139
rect 5976 4109 5998 4139
rect 6036 4109 6044 4139
rect 6044 4109 6070 4139
rect 6108 4109 6112 4139
rect 6112 4109 6142 4139
rect 6180 4109 6214 4139
rect 6252 4109 6282 4139
rect 6282 4109 6286 4139
rect 6324 4109 6350 4139
rect 6350 4109 6358 4139
rect 6396 4109 6418 4139
rect 6418 4109 6430 4139
rect 6468 4109 6486 4139
rect 6486 4109 6502 4139
rect 6540 4109 6554 4139
rect 6554 4109 6574 4139
rect 6612 4109 6622 4139
rect 6622 4109 6646 4139
rect 6684 4109 6690 4139
rect 6690 4109 6718 4139
rect 6756 4109 6758 4139
rect 6758 4109 6790 4139
rect 6828 4109 6860 4139
rect 6860 4109 6862 4139
rect 6900 4109 6928 4139
rect 6928 4109 6934 4139
rect 6972 4109 6996 4139
rect 6996 4109 7006 4139
rect 7044 4109 7064 4139
rect 7064 4109 7078 4139
rect 7116 4109 7132 4139
rect 7132 4109 7150 4139
rect 7188 4109 7200 4139
rect 7200 4109 7222 4139
rect 7260 4109 7268 4139
rect 7268 4109 7294 4139
rect 7332 4109 7336 4139
rect 7336 4109 7366 4139
rect 7404 4109 7438 4139
rect 7476 4109 7506 4139
rect 7506 4109 7510 4139
rect 7548 4109 7574 4139
rect 7574 4109 7582 4139
rect 7620 4109 7642 4139
rect 7642 4109 7654 4139
rect 7692 4109 7710 4139
rect 7710 4109 7726 4139
rect 7764 4109 7778 4139
rect 7778 4109 7798 4139
rect 7836 4109 7846 4139
rect 7846 4109 7870 4139
rect 7908 4109 7914 4139
rect 7914 4109 7942 4139
rect 7980 4109 7982 4139
rect 7982 4109 8014 4139
rect 8052 4109 8084 4139
rect 8084 4109 8086 4139
rect 8124 4109 8152 4139
rect 8152 4109 8158 4139
rect 8196 4109 8220 4139
rect 8220 4109 8230 4139
rect 8268 4109 8288 4139
rect 8288 4109 8302 4139
rect 8340 4109 8356 4139
rect 8356 4109 8374 4139
rect 8412 4109 8424 4139
rect 8424 4109 8446 4139
rect 8484 4109 8492 4139
rect 8492 4109 8518 4139
rect 8556 4109 8560 4139
rect 8560 4109 8590 4139
rect 8628 4109 8662 4139
rect 8700 4109 8730 4139
rect 8730 4109 8734 4139
rect 8772 4109 8798 4139
rect 8798 4109 8806 4139
rect 8844 4109 8866 4139
rect 8866 4109 8878 4139
rect 8916 4109 8934 4139
rect 8934 4109 8950 4139
rect 8988 4109 9002 4139
rect 9002 4109 9022 4139
rect 9060 4109 9070 4139
rect 9070 4109 9094 4139
rect 9132 4109 9138 4139
rect 9138 4109 9166 4139
rect 9204 4109 9206 4139
rect 9206 4109 9238 4139
rect 9276 4109 9308 4139
rect 9308 4109 9310 4139
rect 9348 4109 9376 4139
rect 9376 4109 9382 4139
rect 9420 4109 9444 4139
rect 9444 4109 9454 4139
rect 9492 4109 9512 4139
rect 9512 4109 9526 4139
rect 9564 4109 9580 4139
rect 9580 4109 9598 4139
rect 9636 4109 9648 4139
rect 9648 4109 9670 4139
rect 9708 4109 9716 4139
rect 9716 4109 9742 4139
rect 9780 4109 9784 4139
rect 9784 4109 9814 4139
rect 9852 4109 9886 4139
rect 9924 4109 9954 4139
rect 9954 4109 9958 4139
rect 9996 4109 10022 4139
rect 10022 4109 10030 4139
rect 10068 4109 10090 4139
rect 10090 4109 10102 4139
rect 10140 4109 10158 4139
rect 10158 4109 10174 4139
rect 10212 4109 10226 4139
rect 10226 4109 10246 4139
rect 10284 4109 10294 4139
rect 10294 4109 10318 4139
rect 10356 4109 10362 4139
rect 10362 4109 10390 4139
rect 10428 4109 10430 4139
rect 10430 4109 10462 4139
rect 10500 4109 10532 4139
rect 10532 4109 10534 4139
rect 10572 4109 10600 4139
rect 10600 4109 10606 4139
rect 10644 4109 10668 4139
rect 10668 4109 10678 4139
rect 10716 4109 10736 4139
rect 10736 4109 10750 4139
rect 10788 4109 10804 4139
rect 10804 4109 10822 4139
rect 10860 4109 10872 4139
rect 10872 4109 10894 4139
rect 1985 4105 2019 4109
rect 2058 4105 2092 4109
rect 2131 4105 2165 4109
rect 2204 4105 2238 4109
rect 2277 4105 2311 4109
rect 2350 4105 2384 4109
rect 2423 4105 2457 4109
rect 2496 4105 2530 4109
rect 2569 4105 2603 4109
rect 2642 4105 2676 4109
rect 2715 4105 2749 4109
rect 2788 4105 2822 4109
rect 2861 4105 2895 4109
rect 2934 4105 2968 4109
rect 3007 4105 3041 4109
rect 3080 4105 3114 4109
rect 3153 4105 3187 4109
rect 3226 4105 3260 4109
rect 3299 4105 3333 4109
rect 3372 4105 3406 4109
rect 3444 4105 3478 4109
rect 3516 4105 3550 4109
rect 3588 4105 3622 4109
rect 3660 4105 3694 4109
rect 3732 4105 3766 4109
rect 3804 4105 3838 4109
rect 3876 4105 3910 4109
rect 3948 4105 3982 4109
rect 4020 4105 4054 4109
rect 4092 4105 4126 4109
rect 4164 4105 4198 4109
rect 4236 4105 4270 4109
rect 4308 4105 4342 4109
rect 4380 4105 4414 4109
rect 4452 4105 4486 4109
rect 4524 4105 4558 4109
rect 4596 4105 4630 4109
rect 4668 4105 4702 4109
rect 4740 4105 4774 4109
rect 4812 4105 4846 4109
rect 4884 4105 4918 4109
rect 4956 4105 4990 4109
rect 5028 4105 5062 4109
rect 5100 4105 5134 4109
rect 5172 4105 5206 4109
rect 5244 4105 5278 4109
rect 5316 4105 5350 4109
rect 5388 4105 5422 4109
rect 5460 4105 5494 4109
rect 5532 4105 5566 4109
rect 5604 4105 5638 4109
rect 5676 4105 5710 4109
rect 5748 4105 5782 4109
rect 5820 4105 5854 4109
rect 5892 4105 5926 4109
rect 5964 4105 5998 4109
rect 6036 4105 6070 4109
rect 6108 4105 6142 4109
rect 6180 4105 6214 4109
rect 6252 4105 6286 4109
rect 6324 4105 6358 4109
rect 6396 4105 6430 4109
rect 6468 4105 6502 4109
rect 6540 4105 6574 4109
rect 6612 4105 6646 4109
rect 6684 4105 6718 4109
rect 6756 4105 6790 4109
rect 6828 4105 6862 4109
rect 6900 4105 6934 4109
rect 6972 4105 7006 4109
rect 7044 4105 7078 4109
rect 7116 4105 7150 4109
rect 7188 4105 7222 4109
rect 7260 4105 7294 4109
rect 7332 4105 7366 4109
rect 7404 4105 7438 4109
rect 7476 4105 7510 4109
rect 7548 4105 7582 4109
rect 7620 4105 7654 4109
rect 7692 4105 7726 4109
rect 7764 4105 7798 4109
rect 7836 4105 7870 4109
rect 7908 4105 7942 4109
rect 7980 4105 8014 4109
rect 8052 4105 8086 4109
rect 8124 4105 8158 4109
rect 8196 4105 8230 4109
rect 8268 4105 8302 4109
rect 8340 4105 8374 4109
rect 8412 4105 8446 4109
rect 8484 4105 8518 4109
rect 8556 4105 8590 4109
rect 8628 4105 8662 4109
rect 8700 4105 8734 4109
rect 8772 4105 8806 4109
rect 8844 4105 8878 4109
rect 8916 4105 8950 4109
rect 8988 4105 9022 4109
rect 9060 4105 9094 4109
rect 9132 4105 9166 4109
rect 9204 4105 9238 4109
rect 9276 4105 9310 4109
rect 9348 4105 9382 4109
rect 9420 4105 9454 4109
rect 9492 4105 9526 4109
rect 9564 4105 9598 4109
rect 9636 4105 9670 4109
rect 9708 4105 9742 4109
rect 9780 4105 9814 4109
rect 9852 4105 9886 4109
rect 9924 4105 9958 4109
rect 9996 4105 10030 4109
rect 10068 4105 10102 4109
rect 10140 4105 10174 4109
rect 10212 4105 10246 4109
rect 10284 4105 10318 4109
rect 10356 4105 10390 4109
rect 10428 4105 10462 4109
rect 10500 4105 10534 4109
rect 10572 4105 10606 4109
rect 10644 4105 10678 4109
rect 10716 4105 10750 4109
rect 10788 4105 10822 4109
rect 10860 4105 10894 4109
rect 11624 5854 11626 5872
rect 11626 5854 11658 5872
rect 11696 5854 11728 5872
rect 11728 5854 11730 5872
rect 14526 5854 14528 5888
rect 14528 5854 14560 5888
rect 14598 5854 14630 5888
rect 14630 5854 14632 5888
rect 11624 5838 11658 5854
rect 11696 5838 11730 5854
rect 15733 5845 15754 5850
rect 15754 5845 15767 5850
rect 15819 5845 15824 5850
rect 15824 5845 15853 5850
rect 15905 5845 15928 5850
rect 15928 5845 15939 5850
rect 15991 5845 15998 5850
rect 15998 5845 16025 5850
rect 15733 5816 15767 5845
rect 15819 5816 15853 5845
rect 15905 5816 15939 5845
rect 15991 5816 16025 5845
rect 15733 5776 15754 5778
rect 15754 5776 15767 5778
rect 15819 5776 15824 5778
rect 15824 5776 15853 5778
rect 15905 5776 15928 5778
rect 15928 5776 15939 5778
rect 15991 5776 15998 5778
rect 15998 5776 16025 5778
rect 15733 5744 15767 5776
rect 15819 5744 15853 5776
rect 15905 5744 15939 5776
rect 15991 5744 16025 5776
rect 11624 5700 11626 5734
rect 11626 5700 11658 5734
rect 11696 5700 11728 5734
rect 11728 5700 11730 5734
rect 14526 5700 14528 5734
rect 14528 5700 14560 5734
rect 14598 5700 14630 5734
rect 14630 5700 14632 5734
rect 11500 5572 11506 5599
rect 11506 5572 11534 5599
rect 15733 5672 15767 5706
rect 15819 5672 15853 5706
rect 15905 5672 15939 5706
rect 15991 5672 16025 5706
rect 15733 5603 15767 5634
rect 15819 5603 15853 5634
rect 15905 5603 15939 5634
rect 15991 5603 16025 5634
rect 11500 5565 11534 5572
rect 11624 5546 11626 5580
rect 11626 5546 11658 5580
rect 11696 5546 11728 5580
rect 11728 5546 11730 5580
rect 14526 5546 14528 5580
rect 14528 5546 14560 5580
rect 14598 5546 14630 5580
rect 14630 5546 14632 5580
rect 15733 5600 15754 5603
rect 15754 5600 15767 5603
rect 15819 5600 15824 5603
rect 15824 5600 15853 5603
rect 15905 5600 15928 5603
rect 15928 5600 15939 5603
rect 15991 5600 15998 5603
rect 15998 5600 16025 5603
rect 11500 5503 11506 5525
rect 11506 5503 11534 5525
rect 15733 5534 15767 5562
rect 15819 5534 15853 5562
rect 15905 5534 15939 5562
rect 15991 5534 16025 5562
rect 11500 5491 11534 5503
rect 11500 5434 11506 5451
rect 11506 5434 11534 5451
rect 15733 5528 15754 5534
rect 15754 5528 15767 5534
rect 15819 5528 15824 5534
rect 15824 5528 15853 5534
rect 15905 5528 15928 5534
rect 15928 5528 15939 5534
rect 15991 5528 15998 5534
rect 15998 5528 16025 5534
rect 15733 5465 15767 5490
rect 15819 5465 15853 5490
rect 15905 5465 15939 5490
rect 15991 5465 16025 5490
rect 11500 5417 11534 5434
rect 15733 5456 15754 5465
rect 15754 5456 15767 5465
rect 15819 5456 15824 5465
rect 15824 5456 15853 5465
rect 15905 5456 15928 5465
rect 15928 5456 15939 5465
rect 15991 5456 15998 5465
rect 15998 5456 16025 5465
rect 11500 5365 11506 5377
rect 11506 5365 11534 5377
rect 11624 5392 11626 5426
rect 11626 5392 11658 5426
rect 11696 5392 11728 5426
rect 11728 5392 11730 5426
rect 14526 5392 14528 5426
rect 14528 5392 14560 5426
rect 14598 5392 14630 5426
rect 14630 5392 14632 5426
rect 15733 5396 15767 5418
rect 15819 5396 15853 5418
rect 15905 5396 15939 5418
rect 15991 5396 16025 5418
rect 11500 5343 11534 5365
rect 11500 5296 11506 5303
rect 11506 5296 11534 5303
rect 11500 5269 11534 5296
rect 15733 5384 15754 5396
rect 15754 5384 15767 5396
rect 15819 5384 15824 5396
rect 15824 5384 15853 5396
rect 15905 5384 15928 5396
rect 15928 5384 15939 5396
rect 15991 5384 15998 5396
rect 15998 5384 16025 5396
rect 15733 5327 15767 5346
rect 15819 5327 15853 5346
rect 15905 5327 15939 5346
rect 15991 5327 16025 5346
rect 15733 5312 15754 5327
rect 15754 5312 15767 5327
rect 15819 5312 15824 5327
rect 15824 5312 15853 5327
rect 15905 5312 15928 5327
rect 15928 5312 15939 5327
rect 15991 5312 15998 5327
rect 15998 5312 16025 5327
rect 11500 5227 11506 5229
rect 11506 5227 11534 5229
rect 11624 5238 11626 5272
rect 11626 5238 11658 5272
rect 11696 5238 11728 5272
rect 11728 5238 11730 5272
rect 14526 5238 14528 5272
rect 14528 5238 14560 5272
rect 14598 5238 14630 5272
rect 14630 5238 14632 5272
rect 15733 5258 15767 5274
rect 15819 5258 15853 5274
rect 15905 5258 15939 5274
rect 15991 5258 16025 5274
rect 11500 5195 11534 5227
rect 15733 5240 15754 5258
rect 15754 5240 15767 5258
rect 15819 5240 15824 5258
rect 15824 5240 15853 5258
rect 15905 5240 15928 5258
rect 15928 5240 15939 5258
rect 15991 5240 15998 5258
rect 15998 5240 16025 5258
rect 11500 5123 11534 5155
rect 15733 5190 15767 5202
rect 15819 5190 15853 5202
rect 15905 5190 15939 5202
rect 15991 5190 16025 5202
rect 15733 5168 15754 5190
rect 15754 5168 15767 5190
rect 15819 5168 15824 5190
rect 15824 5168 15853 5190
rect 15905 5168 15928 5190
rect 15928 5168 15939 5190
rect 15991 5168 15998 5190
rect 15998 5168 16025 5190
rect 11500 5121 11506 5123
rect 11506 5121 11534 5123
rect 15733 5122 15767 5130
rect 15819 5122 15853 5130
rect 15905 5122 15939 5130
rect 15991 5122 16025 5130
rect 11624 5084 11626 5118
rect 11626 5084 11658 5118
rect 11696 5084 11728 5118
rect 11728 5084 11730 5118
rect 14526 5084 14528 5118
rect 14528 5084 14560 5118
rect 14598 5084 14630 5118
rect 14630 5084 14632 5118
rect 15733 5096 15754 5122
rect 15754 5096 15767 5122
rect 15819 5096 15824 5122
rect 15824 5096 15853 5122
rect 15905 5096 15928 5122
rect 15928 5096 15939 5122
rect 15991 5096 15998 5122
rect 15998 5096 16025 5122
rect 11500 5054 11534 5081
rect 11500 5047 11506 5054
rect 11506 5047 11534 5054
rect 11500 4985 11534 5007
rect 11500 4973 11506 4985
rect 11506 4973 11534 4985
rect 15733 5054 15767 5058
rect 15819 5054 15853 5058
rect 15905 5054 15939 5058
rect 15991 5054 16025 5058
rect 15733 5024 15754 5054
rect 15754 5024 15767 5054
rect 15819 5024 15824 5054
rect 15824 5024 15853 5054
rect 15905 5024 15928 5054
rect 15928 5024 15939 5054
rect 15991 5024 15998 5054
rect 15998 5024 16025 5054
rect 11500 4916 11534 4933
rect 11624 4930 11626 4964
rect 11626 4930 11658 4964
rect 11696 4930 11728 4964
rect 11728 4930 11730 4964
rect 14526 4930 14528 4964
rect 14528 4930 14560 4964
rect 14598 4930 14630 4964
rect 14630 4930 14632 4964
rect 15733 4952 15754 4986
rect 15754 4952 15767 4986
rect 15819 4952 15824 4986
rect 15824 4952 15853 4986
rect 15905 4952 15928 4986
rect 15928 4952 15939 4986
rect 15991 4952 15998 4986
rect 15998 4952 16025 4986
rect 11500 4899 11506 4916
rect 11506 4899 11534 4916
rect 11500 4847 11534 4859
rect 11500 4825 11506 4847
rect 11506 4825 11534 4847
rect 15733 4884 15754 4914
rect 15754 4884 15767 4914
rect 15819 4884 15824 4914
rect 15824 4884 15853 4914
rect 15905 4884 15928 4914
rect 15928 4884 15939 4914
rect 15991 4884 15998 4914
rect 15998 4884 16025 4914
rect 15733 4880 15767 4884
rect 15819 4880 15853 4884
rect 15905 4880 15939 4884
rect 15991 4880 16025 4884
rect 15733 4816 15754 4842
rect 15754 4816 15767 4842
rect 15819 4816 15824 4842
rect 15824 4816 15853 4842
rect 15905 4816 15928 4842
rect 15928 4816 15939 4842
rect 15991 4816 15998 4842
rect 15998 4816 16025 4842
rect 11500 4778 11534 4786
rect 11500 4752 11506 4778
rect 11506 4752 11534 4778
rect 11624 4776 11626 4810
rect 11626 4776 11658 4810
rect 11696 4776 11728 4810
rect 11728 4776 11730 4810
rect 14526 4776 14528 4810
rect 14528 4776 14560 4810
rect 14598 4776 14630 4810
rect 14630 4776 14632 4810
rect 15733 4808 15767 4816
rect 15819 4808 15853 4816
rect 15905 4808 15939 4816
rect 15991 4808 16025 4816
rect 11500 4709 11534 4713
rect 11500 4679 11506 4709
rect 11506 4679 11534 4709
rect 15733 4748 15754 4770
rect 15754 4748 15767 4770
rect 15819 4748 15824 4770
rect 15824 4748 15853 4770
rect 15905 4748 15928 4770
rect 15928 4748 15939 4770
rect 15991 4748 15998 4770
rect 15998 4748 16025 4770
rect 15733 4736 15767 4748
rect 15819 4736 15853 4748
rect 15905 4736 15939 4748
rect 15991 4736 16025 4748
rect 15733 4680 15754 4698
rect 15754 4680 15767 4698
rect 15819 4680 15824 4698
rect 15824 4680 15853 4698
rect 15905 4680 15928 4698
rect 15928 4680 15939 4698
rect 15991 4680 15998 4698
rect 15998 4680 16025 4698
rect 15733 4664 15767 4680
rect 15819 4664 15853 4680
rect 15905 4664 15939 4680
rect 15991 4664 16025 4680
rect 11500 4606 11506 4640
rect 11506 4606 11534 4640
rect 11624 4622 11626 4656
rect 11626 4622 11658 4656
rect 11696 4622 11728 4656
rect 11728 4622 11730 4656
rect 14526 4622 14528 4656
rect 14528 4622 14560 4656
rect 14598 4622 14630 4656
rect 14630 4622 14632 4656
rect 15733 4612 15754 4626
rect 15754 4612 15767 4626
rect 15819 4612 15824 4626
rect 15824 4612 15853 4626
rect 15905 4612 15928 4626
rect 15928 4612 15939 4626
rect 15991 4612 15998 4626
rect 15998 4612 16025 4626
rect 11500 4537 11506 4567
rect 11506 4537 11534 4567
rect 11500 4533 11534 4537
rect 15733 4592 15767 4612
rect 15819 4592 15853 4612
rect 15905 4592 15939 4612
rect 15991 4592 16025 4612
rect 15733 4544 15754 4554
rect 15754 4544 15767 4554
rect 15819 4544 15824 4554
rect 15824 4544 15853 4554
rect 15905 4544 15928 4554
rect 15928 4544 15939 4554
rect 15991 4544 15998 4554
rect 15998 4544 16025 4554
rect 15733 4520 15767 4544
rect 15819 4520 15853 4544
rect 15905 4520 15939 4544
rect 15991 4520 16025 4544
rect 11500 4468 11506 4494
rect 11506 4468 11534 4494
rect 11624 4468 11626 4502
rect 11626 4468 11658 4502
rect 11696 4468 11728 4502
rect 11728 4468 11730 4502
rect 14526 4468 14528 4502
rect 14528 4468 14560 4502
rect 14598 4468 14630 4502
rect 14630 4468 14632 4502
rect 15733 4476 15754 4482
rect 15754 4476 15767 4482
rect 15819 4476 15824 4482
rect 15824 4476 15853 4482
rect 15905 4476 15928 4482
rect 15928 4476 15939 4482
rect 15991 4476 15998 4482
rect 15998 4476 16025 4482
rect 11500 4460 11534 4468
rect 11500 4399 11506 4421
rect 11506 4399 11534 4421
rect 11500 4387 11534 4399
rect 15733 4448 15767 4476
rect 15819 4448 15853 4476
rect 15905 4448 15939 4476
rect 15991 4448 16025 4476
rect 15733 4408 15754 4410
rect 15754 4408 15767 4410
rect 15819 4408 15824 4410
rect 15824 4408 15853 4410
rect 15905 4408 15928 4410
rect 15928 4408 15939 4410
rect 15991 4408 15998 4410
rect 15998 4408 16025 4410
rect 15733 4376 15767 4408
rect 15819 4376 15853 4408
rect 15905 4376 15939 4408
rect 15991 4376 16025 4408
rect 11500 4330 11506 4348
rect 11506 4330 11534 4348
rect 11500 4314 11534 4330
rect 11624 4314 11626 4348
rect 11626 4314 11658 4348
rect 11696 4314 11728 4348
rect 11728 4314 11730 4348
rect 14526 4314 14528 4348
rect 14528 4314 14560 4348
rect 14598 4314 14630 4348
rect 14630 4314 14632 4348
rect 15733 4306 15767 4338
rect 15819 4306 15853 4338
rect 15905 4306 15939 4338
rect 15991 4306 16025 4338
rect 11500 4261 11506 4275
rect 11506 4261 11534 4275
rect 11500 4241 11534 4261
rect 11500 4192 11506 4202
rect 11506 4192 11534 4202
rect 15733 4304 15754 4306
rect 15754 4304 15767 4306
rect 15819 4304 15824 4306
rect 15824 4304 15853 4306
rect 15905 4304 15928 4306
rect 15928 4304 15939 4306
rect 15991 4304 15998 4306
rect 15998 4304 16025 4306
rect 15554 4238 15588 4246
rect 15626 4238 15660 4246
rect 15733 4238 15767 4266
rect 15819 4238 15853 4266
rect 15905 4238 15939 4266
rect 15991 4238 16025 4266
rect 15554 4212 15578 4238
rect 15578 4212 15588 4238
rect 15626 4212 15648 4238
rect 15648 4212 15660 4238
rect 15733 4232 15754 4238
rect 15754 4232 15767 4238
rect 15819 4232 15824 4238
rect 15824 4232 15853 4238
rect 15905 4232 15928 4238
rect 15928 4232 15939 4238
rect 15991 4232 15998 4238
rect 15998 4232 16025 4238
rect 11500 4168 11534 4192
rect 11624 4160 11626 4194
rect 11626 4160 11658 4194
rect 11696 4160 11728 4194
rect 11728 4160 11730 4194
rect 14526 4160 14528 4194
rect 14528 4160 14560 4194
rect 14598 4160 14630 4194
rect 14630 4160 14632 4194
rect 15484 4170 15518 4173
rect 15560 4170 15594 4173
rect 15636 4170 15670 4173
rect 15733 4170 15767 4194
rect 15819 4170 15853 4194
rect 15905 4170 15939 4194
rect 15991 4170 16025 4194
rect 11500 4123 11506 4129
rect 11506 4123 11534 4129
rect 11500 4095 11534 4123
rect 11500 4054 11506 4056
rect 11506 4054 11534 4056
rect 11500 4022 11534 4054
rect 15484 4139 15508 4170
rect 15508 4139 15518 4170
rect 15560 4139 15578 4170
rect 15578 4139 15594 4170
rect 15636 4139 15648 4170
rect 15648 4139 15670 4170
rect 15733 4160 15754 4170
rect 15754 4160 15767 4170
rect 15819 4160 15824 4170
rect 15824 4160 15853 4170
rect 15905 4160 15928 4170
rect 15928 4160 15939 4170
rect 15991 4160 15998 4170
rect 15998 4160 16025 4170
rect 15733 4102 15767 4122
rect 15819 4102 15853 4122
rect 15905 4102 15939 4122
rect 15991 4102 16025 4122
rect 15405 4068 15438 4088
rect 15438 4068 15439 4088
rect 15484 4068 15508 4092
rect 15508 4068 15518 4092
rect 15560 4068 15578 4092
rect 15578 4068 15594 4092
rect 15636 4068 15648 4092
rect 15648 4068 15670 4092
rect 15733 4088 15754 4102
rect 15754 4088 15767 4102
rect 15819 4088 15824 4102
rect 15824 4088 15853 4102
rect 15905 4088 15928 4102
rect 15928 4088 15939 4102
rect 15991 4088 15998 4102
rect 15998 4088 16025 4102
rect 15405 4054 15439 4068
rect 15484 4058 15518 4068
rect 15560 4058 15594 4068
rect 15636 4058 15670 4068
rect 11583 4017 11588 4051
rect 11588 4017 11617 4051
rect 11656 4017 11657 4051
rect 11657 4017 11690 4051
rect 11729 4017 11760 4051
rect 11760 4017 11763 4051
rect 11801 4017 11829 4051
rect 11829 4017 11835 4051
rect 11873 4017 11898 4051
rect 11898 4017 11907 4051
rect 11945 4017 11967 4051
rect 11967 4017 11979 4051
rect 12017 4017 12036 4051
rect 12036 4017 12051 4051
rect 12089 4017 12105 4051
rect 12105 4017 12123 4051
rect 12161 4017 12174 4051
rect 12174 4017 12195 4051
rect 12233 4017 12243 4051
rect 12243 4017 12267 4051
rect 12305 4017 12312 4051
rect 12312 4017 12339 4051
rect 12377 4017 12381 4051
rect 12381 4017 12411 4051
rect 12449 4017 12450 4051
rect 12450 4017 12483 4051
rect 12521 4017 12554 4051
rect 12554 4017 12555 4051
rect 12593 4017 12623 4051
rect 12623 4017 12627 4051
rect 12665 4017 12692 4051
rect 12692 4017 12699 4051
rect 12737 4017 12761 4051
rect 12761 4017 12771 4051
rect 12809 4017 12830 4051
rect 12830 4017 12843 4051
rect 12881 4017 12899 4051
rect 12899 4017 12915 4051
rect 12953 4017 12968 4051
rect 12968 4017 12987 4051
rect 13025 4017 13037 4051
rect 13037 4017 13059 4051
rect 13097 4017 13106 4051
rect 13106 4017 13131 4051
rect 13169 4017 13175 4051
rect 13175 4017 13203 4051
rect 13241 4017 13244 4051
rect 13244 4017 13275 4051
rect 13313 4017 13347 4051
rect 13385 4017 13416 4051
rect 13416 4017 13419 4051
rect 13457 4017 13485 4051
rect 13485 4017 13491 4051
rect 13529 4017 13554 4051
rect 13554 4017 13563 4051
rect 13601 4017 13623 4051
rect 13623 4017 13635 4051
rect 13673 4017 13692 4051
rect 13692 4017 13707 4051
rect 13745 4017 13761 4051
rect 13761 4017 13779 4051
rect 13817 4017 13830 4051
rect 13830 4017 13851 4051
rect 13889 4017 13899 4051
rect 13899 4017 13923 4051
rect 13961 4017 13968 4051
rect 13968 4017 13995 4051
rect 14033 4017 14036 4051
rect 14036 4017 14067 4051
rect 14105 4017 14138 4051
rect 14138 4017 14139 4051
rect 14177 4017 14206 4051
rect 14206 4017 14211 4051
rect 14249 4017 14274 4051
rect 14274 4017 14283 4051
rect 14321 4017 14342 4051
rect 14342 4017 14355 4051
rect 14393 4017 14410 4051
rect 14410 4017 14427 4051
rect 14465 4017 14478 4051
rect 14478 4017 14499 4051
rect 14537 4017 14546 4051
rect 14546 4017 14571 4051
rect 14609 4017 14614 4051
rect 14614 4017 14643 4051
rect 14681 4017 14682 4051
rect 14682 4017 14715 4051
rect 14753 4034 14787 4051
rect 14825 4034 14859 4051
rect 14897 4034 14931 4051
rect 14969 4034 15003 4051
rect 15041 4034 15075 4051
rect 15113 4034 15147 4051
rect 15185 4034 15219 4051
rect 15257 4034 15291 4051
rect 15329 4034 15363 4051
rect 15733 4034 15767 4050
rect 15819 4034 15853 4050
rect 15905 4034 15939 4050
rect 15991 4034 16025 4050
rect 14753 4017 14774 4034
rect 14774 4017 14787 4034
rect 14825 4017 14844 4034
rect 14844 4017 14859 4034
rect 14897 4017 14914 4034
rect 14914 4017 14931 4034
rect 14969 4017 14984 4034
rect 14984 4017 15003 4034
rect 15041 4017 15054 4034
rect 15054 4017 15075 4034
rect 15113 4017 15124 4034
rect 15124 4017 15147 4034
rect 15185 4017 15194 4034
rect 15194 4017 15219 4034
rect 15257 4017 15264 4034
rect 15264 4017 15291 4034
rect 15329 4017 15334 4034
rect 15334 4017 15363 4034
rect 379 3906 413 3907
rect 379 3873 394 3906
rect 394 3873 413 3906
rect 452 3875 470 3907
rect 470 3875 486 3907
rect 525 3875 538 3907
rect 538 3875 559 3907
rect 598 3875 606 3907
rect 606 3875 632 3907
rect 671 3875 674 3907
rect 674 3875 705 3907
rect 744 3875 776 3907
rect 776 3875 778 3907
rect 817 3875 844 3907
rect 844 3875 851 3907
rect 890 3875 912 3907
rect 912 3875 924 3907
rect 963 3875 980 3907
rect 980 3875 997 3907
rect 1036 3875 1048 3907
rect 1048 3875 1070 3907
rect 1109 3875 1116 3907
rect 1116 3875 1143 3907
rect 1182 3875 1184 3907
rect 1184 3875 1216 3907
rect 1255 3875 1286 3907
rect 1286 3875 1289 3907
rect 1328 3875 1354 3907
rect 1354 3875 1362 3907
rect 1401 3875 1422 3907
rect 1422 3875 1435 3907
rect 1474 3875 1490 3907
rect 1490 3875 1508 3907
rect 1547 3875 1558 3907
rect 1558 3875 1581 3907
rect 1620 3875 1626 3907
rect 1626 3875 1654 3907
rect 1693 3875 1694 3907
rect 1694 3875 1727 3907
rect 1766 3875 1796 3907
rect 1796 3875 1800 3907
rect 1839 3875 1864 3907
rect 1864 3875 1873 3907
rect 1912 3875 1932 3907
rect 1932 3875 1946 3907
rect 1985 3875 2000 3907
rect 2000 3875 2019 3907
rect 2058 3875 2068 3907
rect 2068 3875 2092 3907
rect 2131 3875 2136 3907
rect 2136 3875 2165 3907
rect 452 3873 486 3875
rect 525 3873 559 3875
rect 598 3873 632 3875
rect 671 3873 705 3875
rect 744 3873 778 3875
rect 817 3873 851 3875
rect 890 3873 924 3875
rect 963 3873 997 3875
rect 1036 3873 1070 3875
rect 1109 3873 1143 3875
rect 1182 3873 1216 3875
rect 1255 3873 1289 3875
rect 1328 3873 1362 3875
rect 1401 3873 1435 3875
rect 1474 3873 1508 3875
rect 1547 3873 1581 3875
rect 1620 3873 1654 3875
rect 1693 3873 1727 3875
rect 1766 3873 1800 3875
rect 1839 3873 1873 3875
rect 1912 3873 1946 3875
rect 1985 3873 2019 3875
rect 2058 3873 2092 3875
rect 2131 3873 2165 3875
rect 2204 3873 2238 3907
rect 2277 3875 2306 3907
rect 2306 3875 2311 3907
rect 2350 3875 2374 3907
rect 2374 3875 2384 3907
rect 2423 3875 2442 3907
rect 2442 3875 2457 3907
rect 2496 3875 2510 3907
rect 2510 3875 2530 3907
rect 2569 3875 2578 3907
rect 2578 3875 2603 3907
rect 2642 3875 2646 3907
rect 2646 3875 2676 3907
rect 2715 3875 2748 3907
rect 2748 3875 2749 3907
rect 2788 3875 2816 3907
rect 2816 3875 2822 3907
rect 2861 3875 2884 3907
rect 2884 3875 2895 3907
rect 2934 3875 2952 3907
rect 2952 3875 2968 3907
rect 3007 3875 3020 3907
rect 3020 3875 3041 3907
rect 3080 3875 3088 3907
rect 3088 3875 3114 3907
rect 3153 3875 3156 3907
rect 3156 3875 3187 3907
rect 3226 3875 3258 3907
rect 3258 3875 3260 3907
rect 3299 3875 3326 3907
rect 3326 3875 3333 3907
rect 3372 3875 3394 3907
rect 3394 3875 3406 3907
rect 3444 3875 3462 3907
rect 3462 3875 3478 3907
rect 3516 3875 3530 3907
rect 3530 3875 3550 3907
rect 3588 3875 3598 3907
rect 3598 3875 3622 3907
rect 3660 3875 3666 3907
rect 3666 3875 3694 3907
rect 3732 3875 3734 3907
rect 3734 3875 3766 3907
rect 3804 3875 3836 3907
rect 3836 3875 3838 3907
rect 3876 3875 3904 3907
rect 3904 3875 3910 3907
rect 3948 3875 3972 3907
rect 3972 3875 3982 3907
rect 4020 3875 4040 3907
rect 4040 3875 4054 3907
rect 4092 3875 4108 3907
rect 4108 3875 4126 3907
rect 4164 3875 4176 3907
rect 4176 3875 4198 3907
rect 4236 3875 4244 3907
rect 4244 3875 4270 3907
rect 4308 3875 4312 3907
rect 4312 3875 4342 3907
rect 2277 3873 2311 3875
rect 2350 3873 2384 3875
rect 2423 3873 2457 3875
rect 2496 3873 2530 3875
rect 2569 3873 2603 3875
rect 2642 3873 2676 3875
rect 2715 3873 2749 3875
rect 2788 3873 2822 3875
rect 2861 3873 2895 3875
rect 2934 3873 2968 3875
rect 3007 3873 3041 3875
rect 3080 3873 3114 3875
rect 3153 3873 3187 3875
rect 3226 3873 3260 3875
rect 3299 3873 3333 3875
rect 3372 3873 3406 3875
rect 3444 3873 3478 3875
rect 3516 3873 3550 3875
rect 3588 3873 3622 3875
rect 3660 3873 3694 3875
rect 3732 3873 3766 3875
rect 3804 3873 3838 3875
rect 3876 3873 3910 3875
rect 3948 3873 3982 3875
rect 4020 3873 4054 3875
rect 4092 3873 4126 3875
rect 4164 3873 4198 3875
rect 4236 3873 4270 3875
rect 4308 3873 4342 3875
rect 4380 3873 4414 3907
rect 4452 3875 4482 3907
rect 4482 3875 4486 3907
rect 4524 3875 4550 3907
rect 4550 3875 4558 3907
rect 4596 3875 4618 3907
rect 4618 3875 4630 3907
rect 4668 3875 4686 3907
rect 4686 3875 4702 3907
rect 4740 3875 4754 3907
rect 4754 3875 4774 3907
rect 4812 3875 4822 3907
rect 4822 3875 4846 3907
rect 4884 3875 4890 3907
rect 4890 3875 4918 3907
rect 4956 3875 4958 3907
rect 4958 3875 4990 3907
rect 5028 3875 5060 3907
rect 5060 3875 5062 3907
rect 5100 3875 5128 3907
rect 5128 3875 5134 3907
rect 5172 3875 5196 3907
rect 5196 3875 5206 3907
rect 5244 3875 5264 3907
rect 5264 3875 5278 3907
rect 5316 3875 5332 3907
rect 5332 3875 5350 3907
rect 5388 3875 5400 3907
rect 5400 3875 5422 3907
rect 5460 3875 5468 3907
rect 5468 3875 5494 3907
rect 5532 3875 5536 3907
rect 5536 3875 5566 3907
rect 4452 3873 4486 3875
rect 4524 3873 4558 3875
rect 4596 3873 4630 3875
rect 4668 3873 4702 3875
rect 4740 3873 4774 3875
rect 4812 3873 4846 3875
rect 4884 3873 4918 3875
rect 4956 3873 4990 3875
rect 5028 3873 5062 3875
rect 5100 3873 5134 3875
rect 5172 3873 5206 3875
rect 5244 3873 5278 3875
rect 5316 3873 5350 3875
rect 5388 3873 5422 3875
rect 5460 3873 5494 3875
rect 5532 3873 5566 3875
rect 5604 3873 5638 3907
rect 5676 3875 5706 3907
rect 5706 3875 5710 3907
rect 5748 3875 5774 3907
rect 5774 3875 5782 3907
rect 5820 3875 5842 3907
rect 5842 3875 5854 3907
rect 5892 3875 5910 3907
rect 5910 3875 5926 3907
rect 5964 3875 5978 3907
rect 5978 3875 5998 3907
rect 6036 3875 6046 3907
rect 6046 3875 6070 3907
rect 6108 3875 6114 3907
rect 6114 3875 6142 3907
rect 6180 3875 6182 3907
rect 6182 3875 6214 3907
rect 6252 3875 6284 3907
rect 6284 3875 6286 3907
rect 6324 3875 6352 3907
rect 6352 3875 6358 3907
rect 6396 3875 6420 3907
rect 6420 3875 6430 3907
rect 6468 3875 6488 3907
rect 6488 3875 6502 3907
rect 6540 3875 6556 3907
rect 6556 3875 6574 3907
rect 6612 3875 6624 3907
rect 6624 3875 6646 3907
rect 6684 3875 6692 3907
rect 6692 3875 6718 3907
rect 6756 3875 6760 3907
rect 6760 3875 6790 3907
rect 5676 3873 5710 3875
rect 5748 3873 5782 3875
rect 5820 3873 5854 3875
rect 5892 3873 5926 3875
rect 5964 3873 5998 3875
rect 6036 3873 6070 3875
rect 6108 3873 6142 3875
rect 6180 3873 6214 3875
rect 6252 3873 6286 3875
rect 6324 3873 6358 3875
rect 6396 3873 6430 3875
rect 6468 3873 6502 3875
rect 6540 3873 6574 3875
rect 6612 3873 6646 3875
rect 6684 3873 6718 3875
rect 6756 3873 6790 3875
rect 6828 3873 6862 3907
rect 6900 3875 6930 3907
rect 6930 3875 6934 3907
rect 6972 3875 6998 3907
rect 6998 3875 7006 3907
rect 7044 3875 7066 3907
rect 7066 3875 7078 3907
rect 7116 3875 7134 3907
rect 7134 3875 7150 3907
rect 7188 3875 7202 3907
rect 7202 3875 7222 3907
rect 7260 3875 7270 3907
rect 7270 3875 7294 3907
rect 7332 3875 7338 3907
rect 7338 3875 7366 3907
rect 7404 3875 7406 3907
rect 7406 3875 7438 3907
rect 7476 3875 7508 3907
rect 7508 3875 7510 3907
rect 7548 3875 7576 3907
rect 7576 3875 7582 3907
rect 7620 3875 7644 3907
rect 7644 3875 7654 3907
rect 7692 3875 7712 3907
rect 7712 3875 7726 3907
rect 7764 3875 7780 3907
rect 7780 3875 7798 3907
rect 7836 3875 7848 3907
rect 7848 3875 7870 3907
rect 7908 3875 7916 3907
rect 7916 3875 7942 3907
rect 7980 3875 7984 3907
rect 7984 3875 8014 3907
rect 6900 3873 6934 3875
rect 6972 3873 7006 3875
rect 7044 3873 7078 3875
rect 7116 3873 7150 3875
rect 7188 3873 7222 3875
rect 7260 3873 7294 3875
rect 7332 3873 7366 3875
rect 7404 3873 7438 3875
rect 7476 3873 7510 3875
rect 7548 3873 7582 3875
rect 7620 3873 7654 3875
rect 7692 3873 7726 3875
rect 7764 3873 7798 3875
rect 7836 3873 7870 3875
rect 7908 3873 7942 3875
rect 7980 3873 8014 3875
rect 8052 3873 8086 3907
rect 8124 3875 8154 3907
rect 8154 3875 8158 3907
rect 8196 3875 8222 3907
rect 8222 3875 8230 3907
rect 8268 3875 8290 3907
rect 8290 3875 8302 3907
rect 8340 3875 8359 3907
rect 8359 3875 8374 3907
rect 8412 3875 8428 3907
rect 8428 3875 8446 3907
rect 8484 3875 8497 3907
rect 8497 3875 8518 3907
rect 8556 3875 8566 3907
rect 8566 3875 8590 3907
rect 8628 3875 8635 3907
rect 8635 3875 8662 3907
rect 8700 3875 8704 3907
rect 8704 3875 8734 3907
rect 8772 3875 8773 3907
rect 8773 3875 8806 3907
rect 8844 3875 8876 3907
rect 8876 3875 8878 3907
rect 8916 3875 8945 3907
rect 8945 3875 8950 3907
rect 8988 3875 9014 3907
rect 9014 3875 9022 3907
rect 9060 3875 9083 3907
rect 9083 3875 9094 3907
rect 9132 3875 9152 3907
rect 9152 3875 9166 3907
rect 9204 3875 9221 3907
rect 9221 3875 9238 3907
rect 9276 3875 9290 3907
rect 9290 3875 9310 3907
rect 9348 3875 9359 3907
rect 9359 3875 9382 3907
rect 9420 3875 9428 3907
rect 9428 3875 9454 3907
rect 9492 3875 9497 3907
rect 9497 3875 9526 3907
rect 9564 3875 9566 3907
rect 9566 3875 9598 3907
rect 8124 3873 8158 3875
rect 8196 3873 8230 3875
rect 8268 3873 8302 3875
rect 8340 3873 8374 3875
rect 8412 3873 8446 3875
rect 8484 3873 8518 3875
rect 8556 3873 8590 3875
rect 8628 3873 8662 3875
rect 8700 3873 8734 3875
rect 8772 3873 8806 3875
rect 8844 3873 8878 3875
rect 8916 3873 8950 3875
rect 8988 3873 9022 3875
rect 9060 3873 9094 3875
rect 9132 3873 9166 3875
rect 9204 3873 9238 3875
rect 9276 3873 9310 3875
rect 9348 3873 9382 3875
rect 9420 3873 9454 3875
rect 9492 3873 9526 3875
rect 9564 3873 9598 3875
rect 9636 3873 9670 3907
rect 9708 3875 9739 3907
rect 9739 3875 9742 3907
rect 9780 3875 9808 3907
rect 9808 3875 9814 3907
rect 9852 3875 9877 3907
rect 9877 3875 9886 3907
rect 9924 3875 9946 3907
rect 9946 3875 9958 3907
rect 9996 3875 10015 3907
rect 10015 3875 10030 3907
rect 10068 3875 10084 3907
rect 10084 3875 10102 3907
rect 10140 3875 10153 3907
rect 10153 3875 10174 3907
rect 10212 3875 10222 3907
rect 10222 3875 10246 3907
rect 10284 3875 10291 3907
rect 10291 3875 10318 3907
rect 10356 3875 10360 3907
rect 10360 3875 10390 3907
rect 10428 3875 10429 3907
rect 10429 3875 10462 3907
rect 10500 3875 10532 3907
rect 10532 3875 10534 3907
rect 10572 3875 10601 3907
rect 10601 3875 10606 3907
rect 10644 3875 10670 3907
rect 10670 3875 10678 3907
rect 10716 3875 10739 3907
rect 10739 3875 10750 3907
rect 10788 3875 10808 3907
rect 10808 3875 10822 3907
rect 10860 3875 10877 3907
rect 10877 3875 10894 3907
rect 9708 3873 9742 3875
rect 9780 3873 9814 3875
rect 9852 3873 9886 3875
rect 9924 3873 9958 3875
rect 9996 3873 10030 3875
rect 10068 3873 10102 3875
rect 10140 3873 10174 3875
rect 10212 3873 10246 3875
rect 10284 3873 10318 3875
rect 10356 3873 10390 3875
rect 10428 3873 10462 3875
rect 10500 3873 10534 3875
rect 10572 3873 10606 3875
rect 10644 3873 10678 3875
rect 10716 3873 10750 3875
rect 10788 3873 10822 3875
rect 10860 3873 10894 3875
rect 360 3764 394 3790
rect 360 3756 394 3764
rect 552 3769 586 3803
rect 632 3769 656 3803
rect 656 3769 666 3803
rect 711 3769 724 3803
rect 724 3769 745 3803
rect 790 3769 792 3803
rect 792 3769 824 3803
rect 869 3769 894 3803
rect 894 3769 903 3803
rect 948 3769 962 3803
rect 962 3769 982 3803
rect 1027 3769 1030 3803
rect 1030 3769 1061 3803
rect 1106 3769 1132 3803
rect 1132 3769 1140 3803
rect 1185 3769 1200 3803
rect 1200 3769 1219 3803
rect 1264 3769 1268 3803
rect 1268 3769 1298 3803
rect 1408 3769 1442 3803
rect 1488 3769 1512 3803
rect 1512 3769 1522 3803
rect 1567 3769 1580 3803
rect 1580 3769 1601 3803
rect 1646 3769 1648 3803
rect 1648 3769 1680 3803
rect 1725 3769 1750 3803
rect 1750 3769 1759 3803
rect 1804 3769 1818 3803
rect 1818 3769 1838 3803
rect 1883 3769 1886 3803
rect 1886 3769 1917 3803
rect 1962 3769 1988 3803
rect 1988 3769 1996 3803
rect 2041 3769 2056 3803
rect 2056 3769 2075 3803
rect 2120 3769 2124 3803
rect 2124 3769 2154 3803
rect 2264 3769 2298 3803
rect 2344 3769 2368 3803
rect 2368 3769 2378 3803
rect 2423 3769 2436 3803
rect 2436 3769 2457 3803
rect 2502 3769 2504 3803
rect 2504 3769 2536 3803
rect 2581 3769 2606 3803
rect 2606 3769 2615 3803
rect 2660 3769 2674 3803
rect 2674 3769 2694 3803
rect 2739 3769 2742 3803
rect 2742 3769 2773 3803
rect 2818 3769 2844 3803
rect 2844 3769 2852 3803
rect 2897 3769 2912 3803
rect 2912 3769 2931 3803
rect 2976 3769 2980 3803
rect 2980 3769 3010 3803
rect 3120 3769 3154 3803
rect 3200 3769 3224 3803
rect 3224 3769 3234 3803
rect 3279 3769 3292 3803
rect 3292 3769 3313 3803
rect 3358 3769 3360 3803
rect 3360 3769 3392 3803
rect 3437 3769 3462 3803
rect 3462 3769 3471 3803
rect 3516 3769 3530 3803
rect 3530 3769 3550 3803
rect 3595 3769 3598 3803
rect 3598 3769 3629 3803
rect 3674 3769 3700 3803
rect 3700 3769 3708 3803
rect 3753 3769 3768 3803
rect 3768 3769 3787 3803
rect 3832 3769 3836 3803
rect 3836 3769 3866 3803
rect 3976 3769 4010 3803
rect 4056 3769 4080 3803
rect 4080 3769 4090 3803
rect 4135 3769 4148 3803
rect 4148 3769 4169 3803
rect 4214 3769 4216 3803
rect 4216 3769 4248 3803
rect 4293 3769 4318 3803
rect 4318 3769 4327 3803
rect 4372 3769 4386 3803
rect 4386 3769 4406 3803
rect 4451 3769 4454 3803
rect 4454 3769 4485 3803
rect 4530 3769 4556 3803
rect 4556 3769 4564 3803
rect 4609 3769 4624 3803
rect 4624 3769 4643 3803
rect 4688 3769 4692 3803
rect 4692 3769 4722 3803
rect 4832 3769 4866 3803
rect 4912 3769 4936 3803
rect 4936 3769 4946 3803
rect 4991 3769 5004 3803
rect 5004 3769 5025 3803
rect 5070 3769 5072 3803
rect 5072 3769 5104 3803
rect 5149 3769 5174 3803
rect 5174 3769 5183 3803
rect 5228 3769 5242 3803
rect 5242 3769 5262 3803
rect 5307 3769 5310 3803
rect 5310 3769 5341 3803
rect 5386 3769 5412 3803
rect 5412 3769 5420 3803
rect 5465 3769 5480 3803
rect 5480 3769 5499 3803
rect 5544 3769 5548 3803
rect 5548 3769 5578 3803
rect 5688 3769 5722 3803
rect 5768 3769 5792 3803
rect 5792 3769 5802 3803
rect 5847 3769 5860 3803
rect 5860 3769 5881 3803
rect 5926 3769 5928 3803
rect 5928 3769 5960 3803
rect 6005 3769 6030 3803
rect 6030 3769 6039 3803
rect 6084 3769 6098 3803
rect 6098 3769 6118 3803
rect 6163 3769 6166 3803
rect 6166 3769 6197 3803
rect 6242 3769 6268 3803
rect 6268 3769 6276 3803
rect 6321 3769 6336 3803
rect 6336 3769 6355 3803
rect 6400 3769 6404 3803
rect 6404 3769 6434 3803
rect 6544 3769 6578 3803
rect 6624 3769 6648 3803
rect 6648 3769 6658 3803
rect 6703 3769 6716 3803
rect 6716 3769 6737 3803
rect 6782 3769 6784 3803
rect 6784 3769 6816 3803
rect 6861 3769 6886 3803
rect 6886 3769 6895 3803
rect 6940 3769 6954 3803
rect 6954 3769 6974 3803
rect 7019 3769 7022 3803
rect 7022 3769 7053 3803
rect 7098 3769 7124 3803
rect 7124 3769 7132 3803
rect 7177 3769 7192 3803
rect 7192 3769 7211 3803
rect 7256 3769 7260 3803
rect 7260 3769 7290 3803
rect 7400 3769 7434 3803
rect 7480 3769 7504 3803
rect 7504 3769 7514 3803
rect 7559 3769 7572 3803
rect 7572 3769 7593 3803
rect 7638 3769 7640 3803
rect 7640 3769 7672 3803
rect 7717 3769 7742 3803
rect 7742 3769 7751 3803
rect 7796 3769 7810 3803
rect 7810 3769 7830 3803
rect 7875 3769 7878 3803
rect 7878 3769 7909 3803
rect 7954 3769 7980 3803
rect 7980 3769 7988 3803
rect 8033 3769 8048 3803
rect 8048 3769 8067 3803
rect 8112 3769 8116 3803
rect 8116 3769 8146 3803
rect 8256 3769 8290 3803
rect 8336 3769 8360 3803
rect 8360 3769 8370 3803
rect 8415 3769 8428 3803
rect 8428 3769 8449 3803
rect 8494 3769 8496 3803
rect 8496 3769 8528 3803
rect 8573 3769 8598 3803
rect 8598 3769 8607 3803
rect 8652 3769 8666 3803
rect 8666 3769 8686 3803
rect 8731 3769 8734 3803
rect 8734 3769 8765 3803
rect 8810 3769 8836 3803
rect 8836 3769 8844 3803
rect 8889 3769 8904 3803
rect 8904 3769 8923 3803
rect 8968 3769 8972 3803
rect 8972 3769 9002 3803
rect 9112 3769 9146 3803
rect 9192 3769 9216 3803
rect 9216 3769 9226 3803
rect 9271 3769 9284 3803
rect 9284 3769 9305 3803
rect 9350 3769 9352 3803
rect 9352 3769 9384 3803
rect 9429 3769 9454 3803
rect 9454 3769 9463 3803
rect 9508 3769 9522 3803
rect 9522 3769 9542 3803
rect 9587 3769 9590 3803
rect 9590 3769 9621 3803
rect 9666 3769 9692 3803
rect 9692 3769 9700 3803
rect 9745 3769 9760 3803
rect 9760 3769 9779 3803
rect 9824 3769 9828 3803
rect 9828 3769 9858 3803
rect 9968 3769 10002 3803
rect 10048 3769 10072 3803
rect 10072 3769 10082 3803
rect 10127 3769 10140 3803
rect 10140 3769 10161 3803
rect 10206 3769 10208 3803
rect 10208 3769 10240 3803
rect 10285 3769 10310 3803
rect 10310 3769 10319 3803
rect 10364 3769 10378 3803
rect 10378 3769 10398 3803
rect 10443 3769 10446 3803
rect 10446 3769 10477 3803
rect 10522 3769 10548 3803
rect 10548 3769 10556 3803
rect 10601 3769 10616 3803
rect 10616 3769 10635 3803
rect 10680 3769 10684 3803
rect 10684 3769 10714 3803
rect 360 3693 394 3718
rect 360 3684 394 3693
rect 10912 3769 10946 3790
rect 10912 3756 10946 3769
rect 360 3623 394 3646
rect 360 3612 394 3623
rect 360 3553 394 3574
rect 360 3540 394 3553
rect 360 3483 394 3502
rect 360 3468 394 3483
rect 360 3413 394 3430
rect 360 3396 394 3413
rect 360 3343 394 3358
rect 360 3324 394 3343
rect 360 3273 394 3286
rect 360 3252 394 3273
rect 360 3203 394 3214
rect 360 3180 394 3203
rect 360 3133 394 3142
rect 360 3108 394 3133
rect 360 3063 394 3070
rect 360 3036 394 3063
rect 360 2993 394 2998
rect 360 2964 394 2993
rect 360 2923 394 2926
rect 360 2892 394 2923
rect 360 2853 394 2854
rect 360 2820 394 2853
rect 360 2749 394 2782
rect 360 2748 394 2749
rect 360 2679 394 2710
rect 360 2676 394 2679
rect 360 2609 394 2638
rect 360 2604 394 2609
rect 360 2539 394 2566
rect 360 2532 394 2539
rect 360 2469 394 2494
rect 360 2460 394 2469
rect 360 2399 394 2422
rect 360 2388 394 2399
rect 360 2329 394 2350
rect 360 2316 394 2329
rect 500 3625 534 3646
rect 500 3612 534 3625
rect 500 3557 534 3574
rect 500 3540 534 3557
rect 500 3489 534 3502
rect 500 3468 534 3489
rect 500 3421 534 3430
rect 500 3396 534 3421
rect 500 3353 534 3358
rect 500 3324 534 3353
rect 500 3285 534 3286
rect 500 3252 534 3285
rect 500 3183 534 3214
rect 500 3180 534 3183
rect 500 3115 534 3142
rect 500 3108 534 3115
rect 500 3047 534 3070
rect 500 3036 534 3047
rect 500 2979 534 2998
rect 500 2964 534 2979
rect 500 2911 534 2926
rect 500 2892 534 2911
rect 500 2843 534 2854
rect 500 2820 534 2843
rect 500 2775 534 2782
rect 500 2748 534 2775
rect 1356 3659 1390 3664
rect 1356 3630 1390 3659
rect 1356 3591 1390 3592
rect 1356 3558 1390 3591
rect 1356 3489 1390 3520
rect 1356 3486 1390 3489
rect 1356 3421 1390 3448
rect 1356 3414 1390 3421
rect 1356 3353 1390 3376
rect 1356 3342 1390 3353
rect 1356 3285 1390 3304
rect 1356 3270 1390 3285
rect 1356 3217 1390 3232
rect 1356 3198 1390 3217
rect 1356 3149 1390 3160
rect 1356 3126 1390 3149
rect 1356 3081 1390 3088
rect 1356 3054 1390 3081
rect 1356 3013 1390 3016
rect 1356 2982 1390 3013
rect 1356 2911 1390 2944
rect 1356 2910 1390 2911
rect 1356 2843 1390 2872
rect 1356 2838 1390 2843
rect 1356 2775 1390 2800
rect 1356 2766 1390 2775
rect 1356 2707 1390 2728
rect 1356 2694 1390 2707
rect 1356 2639 1390 2656
rect 1356 2622 1390 2639
rect 1356 2571 1390 2584
rect 1356 2550 1390 2571
rect 1356 2503 1390 2512
rect 1356 2478 1390 2503
rect 1356 2435 1390 2440
rect 1356 2406 1390 2435
rect 1356 2367 1390 2368
rect 1356 2334 1390 2367
rect 2212 3659 2246 3664
rect 2212 3630 2246 3659
rect 2212 3591 2246 3592
rect 2212 3558 2246 3591
rect 2212 3489 2246 3520
rect 2212 3486 2246 3489
rect 2212 3421 2246 3448
rect 2212 3414 2246 3421
rect 2212 3353 2246 3376
rect 2212 3342 2246 3353
rect 2212 3285 2246 3304
rect 2212 3270 2246 3285
rect 2212 3217 2246 3232
rect 2212 3198 2246 3217
rect 2212 3149 2246 3160
rect 2212 3126 2246 3149
rect 2212 3081 2246 3088
rect 2212 3054 2246 3081
rect 2212 3013 2246 3016
rect 2212 2982 2246 3013
rect 2212 2911 2246 2944
rect 2212 2910 2246 2911
rect 2212 2843 2246 2872
rect 2212 2838 2246 2843
rect 2212 2775 2246 2800
rect 2212 2766 2246 2775
rect 2212 2707 2246 2728
rect 2212 2694 2246 2707
rect 2212 2639 2246 2656
rect 2212 2622 2246 2639
rect 2212 2571 2246 2584
rect 2212 2550 2246 2571
rect 2212 2503 2246 2512
rect 2212 2478 2246 2503
rect 2212 2435 2246 2440
rect 2212 2406 2246 2435
rect 2212 2367 2246 2368
rect 2212 2334 2246 2367
rect 3068 3659 3102 3664
rect 3068 3630 3102 3659
rect 3068 3591 3102 3592
rect 3068 3558 3102 3591
rect 3068 3489 3102 3520
rect 3068 3486 3102 3489
rect 3068 3421 3102 3448
rect 3068 3414 3102 3421
rect 3068 3353 3102 3376
rect 3068 3342 3102 3353
rect 3068 3285 3102 3304
rect 3068 3270 3102 3285
rect 3068 3217 3102 3232
rect 3068 3198 3102 3217
rect 3068 3149 3102 3160
rect 3068 3126 3102 3149
rect 3068 3081 3102 3088
rect 3068 3054 3102 3081
rect 3068 3013 3102 3016
rect 3068 2982 3102 3013
rect 3068 2911 3102 2944
rect 3068 2910 3102 2911
rect 3068 2843 3102 2872
rect 3068 2838 3102 2843
rect 3068 2775 3102 2800
rect 3068 2766 3102 2775
rect 3068 2707 3102 2728
rect 3068 2694 3102 2707
rect 3068 2639 3102 2656
rect 3068 2622 3102 2639
rect 3068 2571 3102 2584
rect 3068 2550 3102 2571
rect 3068 2503 3102 2512
rect 3068 2478 3102 2503
rect 3068 2435 3102 2440
rect 3068 2406 3102 2435
rect 3068 2367 3102 2368
rect 3068 2334 3102 2367
rect 3924 3659 3958 3664
rect 3924 3630 3958 3659
rect 3924 3591 3958 3592
rect 3924 3558 3958 3591
rect 3924 3489 3958 3520
rect 3924 3486 3958 3489
rect 3924 3421 3958 3448
rect 3924 3414 3958 3421
rect 3924 3353 3958 3376
rect 3924 3342 3958 3353
rect 3924 3285 3958 3304
rect 3924 3270 3958 3285
rect 3924 3217 3958 3232
rect 3924 3198 3958 3217
rect 3924 3149 3958 3160
rect 3924 3126 3958 3149
rect 3924 3081 3958 3088
rect 3924 3054 3958 3081
rect 3924 3013 3958 3016
rect 3924 2982 3958 3013
rect 3924 2911 3958 2944
rect 3924 2910 3958 2911
rect 3924 2843 3958 2872
rect 3924 2838 3958 2843
rect 3924 2775 3958 2800
rect 3924 2766 3958 2775
rect 3924 2707 3958 2728
rect 3924 2694 3958 2707
rect 3924 2639 3958 2656
rect 3924 2622 3958 2639
rect 3924 2571 3958 2584
rect 3924 2550 3958 2571
rect 3924 2503 3958 2512
rect 3924 2478 3958 2503
rect 3924 2435 3958 2440
rect 3924 2406 3958 2435
rect 3924 2367 3958 2368
rect 3924 2334 3958 2367
rect 4780 3659 4814 3664
rect 4780 3630 4814 3659
rect 4780 3591 4814 3592
rect 4780 3558 4814 3591
rect 4780 3489 4814 3520
rect 4780 3486 4814 3489
rect 4780 3421 4814 3448
rect 4780 3414 4814 3421
rect 4780 3353 4814 3376
rect 4780 3342 4814 3353
rect 4780 3285 4814 3304
rect 4780 3270 4814 3285
rect 4780 3217 4814 3232
rect 4780 3198 4814 3217
rect 4780 3149 4814 3160
rect 4780 3126 4814 3149
rect 4780 3081 4814 3088
rect 4780 3054 4814 3081
rect 4780 3013 4814 3016
rect 4780 2982 4814 3013
rect 4780 2911 4814 2944
rect 4780 2910 4814 2911
rect 4780 2843 4814 2872
rect 4780 2838 4814 2843
rect 4780 2775 4814 2800
rect 4780 2766 4814 2775
rect 4780 2707 4814 2728
rect 4780 2694 4814 2707
rect 4780 2639 4814 2656
rect 4780 2622 4814 2639
rect 4780 2571 4814 2584
rect 4780 2550 4814 2571
rect 4780 2503 4814 2512
rect 4780 2478 4814 2503
rect 4780 2435 4814 2440
rect 4780 2406 4814 2435
rect 4780 2367 4814 2368
rect 4780 2334 4814 2367
rect 5636 3659 5670 3664
rect 5636 3630 5670 3659
rect 5636 3591 5670 3592
rect 5636 3558 5670 3591
rect 5636 3489 5670 3520
rect 5636 3486 5670 3489
rect 5636 3421 5670 3448
rect 5636 3414 5670 3421
rect 5636 3353 5670 3376
rect 5636 3342 5670 3353
rect 5636 3285 5670 3304
rect 5636 3270 5670 3285
rect 5636 3217 5670 3232
rect 5636 3198 5670 3217
rect 5636 3149 5670 3160
rect 5636 3126 5670 3149
rect 5636 3081 5670 3088
rect 5636 3054 5670 3081
rect 5636 3013 5670 3016
rect 5636 2982 5670 3013
rect 5636 2911 5670 2944
rect 5636 2910 5670 2911
rect 5636 2843 5670 2872
rect 5636 2838 5670 2843
rect 5636 2775 5670 2800
rect 5636 2766 5670 2775
rect 5636 2707 5670 2728
rect 5636 2694 5670 2707
rect 5636 2639 5670 2656
rect 5636 2622 5670 2639
rect 5636 2571 5670 2584
rect 5636 2550 5670 2571
rect 5636 2503 5670 2512
rect 5636 2478 5670 2503
rect 5636 2435 5670 2440
rect 5636 2406 5670 2435
rect 5636 2367 5670 2368
rect 5636 2334 5670 2367
rect 6492 3659 6526 3664
rect 6492 3630 6526 3659
rect 6492 3591 6526 3592
rect 6492 3558 6526 3591
rect 6492 3489 6526 3520
rect 6492 3486 6526 3489
rect 6492 3421 6526 3448
rect 6492 3414 6526 3421
rect 6492 3353 6526 3376
rect 6492 3342 6526 3353
rect 6492 3285 6526 3304
rect 6492 3270 6526 3285
rect 6492 3217 6526 3232
rect 6492 3198 6526 3217
rect 6492 3149 6526 3160
rect 6492 3126 6526 3149
rect 6492 3081 6526 3088
rect 6492 3054 6526 3081
rect 6492 3013 6526 3016
rect 6492 2982 6526 3013
rect 6492 2911 6526 2944
rect 6492 2910 6526 2911
rect 6492 2843 6526 2872
rect 6492 2838 6526 2843
rect 6492 2775 6526 2800
rect 6492 2766 6526 2775
rect 6492 2707 6526 2728
rect 6492 2694 6526 2707
rect 6492 2639 6526 2656
rect 6492 2622 6526 2639
rect 6492 2571 6526 2584
rect 6492 2550 6526 2571
rect 6492 2503 6526 2512
rect 6492 2478 6526 2503
rect 6492 2435 6526 2440
rect 6492 2406 6526 2435
rect 6492 2367 6526 2368
rect 6492 2334 6526 2367
rect 7348 3659 7382 3664
rect 7348 3630 7382 3659
rect 7348 3591 7382 3592
rect 7348 3558 7382 3591
rect 7348 3489 7382 3520
rect 7348 3486 7382 3489
rect 7348 3421 7382 3448
rect 7348 3414 7382 3421
rect 7348 3353 7382 3376
rect 7348 3342 7382 3353
rect 7348 3285 7382 3304
rect 7348 3270 7382 3285
rect 7348 3217 7382 3232
rect 7348 3198 7382 3217
rect 7348 3149 7382 3160
rect 7348 3126 7382 3149
rect 7348 3081 7382 3088
rect 7348 3054 7382 3081
rect 7348 3013 7382 3016
rect 7348 2982 7382 3013
rect 7348 2911 7382 2944
rect 7348 2910 7382 2911
rect 7348 2843 7382 2872
rect 7348 2838 7382 2843
rect 7348 2775 7382 2800
rect 7348 2766 7382 2775
rect 7348 2707 7382 2728
rect 7348 2694 7382 2707
rect 7348 2639 7382 2656
rect 7348 2622 7382 2639
rect 7348 2571 7382 2584
rect 7348 2550 7382 2571
rect 7348 2503 7382 2512
rect 7348 2478 7382 2503
rect 7348 2435 7382 2440
rect 7348 2406 7382 2435
rect 7348 2367 7382 2368
rect 7348 2334 7382 2367
rect 8204 3659 8238 3664
rect 8204 3630 8238 3659
rect 8204 3591 8238 3592
rect 8204 3558 8238 3591
rect 8204 3489 8238 3520
rect 8204 3486 8238 3489
rect 8204 3421 8238 3448
rect 8204 3414 8238 3421
rect 8204 3353 8238 3376
rect 8204 3342 8238 3353
rect 8204 3285 8238 3304
rect 8204 3270 8238 3285
rect 8204 3217 8238 3232
rect 8204 3198 8238 3217
rect 8204 3149 8238 3160
rect 8204 3126 8238 3149
rect 8204 3081 8238 3088
rect 8204 3054 8238 3081
rect 8204 3013 8238 3016
rect 8204 2982 8238 3013
rect 8204 2911 8238 2944
rect 8204 2910 8238 2911
rect 8204 2843 8238 2872
rect 8204 2838 8238 2843
rect 8204 2775 8238 2800
rect 8204 2766 8238 2775
rect 8204 2707 8238 2728
rect 8204 2694 8238 2707
rect 8204 2639 8238 2656
rect 8204 2622 8238 2639
rect 8204 2571 8238 2584
rect 8204 2550 8238 2571
rect 8204 2503 8238 2512
rect 8204 2478 8238 2503
rect 8204 2435 8238 2440
rect 8204 2406 8238 2435
rect 8204 2367 8238 2368
rect 8204 2334 8238 2367
rect 9060 3659 9094 3664
rect 9060 3630 9094 3659
rect 9060 3591 9094 3592
rect 9060 3558 9094 3591
rect 9060 3489 9094 3520
rect 9060 3486 9094 3489
rect 9060 3421 9094 3448
rect 9060 3414 9094 3421
rect 9060 3353 9094 3376
rect 9060 3342 9094 3353
rect 9060 3285 9094 3304
rect 9060 3270 9094 3285
rect 9060 3217 9094 3232
rect 9060 3198 9094 3217
rect 9060 3149 9094 3160
rect 9060 3126 9094 3149
rect 9060 3081 9094 3088
rect 9060 3054 9094 3081
rect 9060 3013 9094 3016
rect 9060 2982 9094 3013
rect 9060 2911 9094 2944
rect 9060 2910 9094 2911
rect 9060 2843 9094 2872
rect 9060 2838 9094 2843
rect 9060 2775 9094 2800
rect 9060 2766 9094 2775
rect 9060 2707 9094 2728
rect 9060 2694 9094 2707
rect 9060 2639 9094 2656
rect 9060 2622 9094 2639
rect 9060 2571 9094 2584
rect 9060 2550 9094 2571
rect 9060 2503 9094 2512
rect 9060 2478 9094 2503
rect 9060 2435 9094 2440
rect 9060 2406 9094 2435
rect 9060 2367 9094 2368
rect 9060 2334 9094 2367
rect 9916 3659 9950 3664
rect 9916 3630 9950 3659
rect 9916 3591 9950 3592
rect 9916 3558 9950 3591
rect 9916 3489 9950 3520
rect 9916 3486 9950 3489
rect 9916 3421 9950 3448
rect 9916 3414 9950 3421
rect 9916 3353 9950 3376
rect 9916 3342 9950 3353
rect 9916 3285 9950 3304
rect 9916 3270 9950 3285
rect 9916 3217 9950 3232
rect 9916 3198 9950 3217
rect 9916 3149 9950 3160
rect 9916 3126 9950 3149
rect 9916 3081 9950 3088
rect 9916 3054 9950 3081
rect 9916 3013 9950 3016
rect 9916 2982 9950 3013
rect 9916 2911 9950 2944
rect 9916 2910 9950 2911
rect 9916 2843 9950 2872
rect 9916 2838 9950 2843
rect 9916 2775 9950 2800
rect 9916 2766 9950 2775
rect 9916 2707 9950 2728
rect 9916 2694 9950 2707
rect 9916 2639 9950 2656
rect 9916 2622 9950 2639
rect 9916 2571 9950 2584
rect 9916 2550 9950 2571
rect 9916 2503 9950 2512
rect 9916 2478 9950 2503
rect 9916 2435 9950 2440
rect 9916 2406 9950 2435
rect 9916 2367 9950 2368
rect 9916 2334 9950 2367
rect 10772 3659 10806 3664
rect 10772 3630 10806 3659
rect 10772 3591 10806 3592
rect 10772 3558 10806 3591
rect 10772 3489 10806 3520
rect 10772 3486 10806 3489
rect 10772 3421 10806 3448
rect 10772 3414 10806 3421
rect 10772 3353 10806 3376
rect 10772 3342 10806 3353
rect 10772 3285 10806 3304
rect 10772 3270 10806 3285
rect 10772 3217 10806 3232
rect 10772 3198 10806 3217
rect 10772 3149 10806 3160
rect 10772 3126 10806 3149
rect 10772 3081 10806 3088
rect 10772 3054 10806 3081
rect 10772 3013 10806 3016
rect 10772 2982 10806 3013
rect 10772 2911 10806 2944
rect 10772 2910 10806 2911
rect 10772 2843 10806 2872
rect 10772 2838 10806 2843
rect 10772 2775 10806 2800
rect 10772 2766 10806 2775
rect 10772 2707 10806 2728
rect 10772 2694 10806 2707
rect 10772 2639 10806 2656
rect 10772 2622 10806 2639
rect 10772 2571 10806 2584
rect 10772 2550 10806 2571
rect 10772 2503 10806 2512
rect 10772 2478 10806 2503
rect 10772 2435 10806 2440
rect 10772 2406 10806 2435
rect 10772 2367 10806 2368
rect 10772 2334 10806 2367
rect 10912 3699 10946 3718
rect 10912 3684 10946 3699
rect 10912 3629 10946 3646
rect 10912 3612 10946 3629
rect 10912 3559 10946 3574
rect 10912 3540 10946 3559
rect 10912 3489 10946 3502
rect 10912 3468 10946 3489
rect 10912 3419 10946 3430
rect 10912 3396 10946 3419
rect 10912 3349 10946 3358
rect 10912 3324 10946 3349
rect 10912 3279 10946 3286
rect 10912 3252 10946 3279
rect 10912 3209 10946 3214
rect 10912 3180 10946 3209
rect 10912 3139 10946 3142
rect 10912 3108 10946 3139
rect 10912 3069 10946 3070
rect 10912 3036 10946 3069
rect 10912 2965 10946 2998
rect 10912 2964 10946 2965
rect 10912 2895 10946 2926
rect 10912 2892 10946 2895
rect 10912 2825 10946 2854
rect 10912 2820 10946 2825
rect 10912 2755 10946 2782
rect 10912 2748 10946 2755
rect 10912 2685 10946 2710
rect 10912 2676 10946 2685
rect 10912 2615 10946 2638
rect 10912 2604 10946 2615
rect 10912 2544 10946 2566
rect 10912 2532 10946 2544
rect 10912 2473 10946 2494
rect 10912 2460 10946 2473
rect 10912 2402 10946 2422
rect 10912 2388 10946 2402
rect 360 2259 394 2278
rect 360 2244 394 2259
rect 10912 2331 10946 2350
rect 10912 2316 10946 2331
rect 456 2189 463 2223
rect 463 2189 490 2223
rect 528 2189 532 2223
rect 532 2189 562 2223
rect 600 2189 601 2223
rect 601 2189 634 2223
rect 1069 2189 1084 2223
rect 1084 2189 1103 2223
rect 1141 2189 1153 2223
rect 1153 2189 1175 2223
rect 1213 2189 1222 2223
rect 1222 2189 1247 2223
rect 1458 2189 1460 2223
rect 1460 2189 1492 2223
rect 1530 2189 1562 2223
rect 1562 2189 1564 2223
rect 1602 2189 1630 2223
rect 1630 2189 1636 2223
rect 1912 2189 1936 2223
rect 1936 2189 1946 2223
rect 1984 2189 2004 2223
rect 2004 2189 2018 2223
rect 2056 2189 2072 2223
rect 2072 2189 2090 2223
rect 2317 2189 2344 2223
rect 2344 2189 2351 2223
rect 2389 2189 2412 2223
rect 2412 2189 2423 2223
rect 2461 2189 2480 2223
rect 2480 2189 2495 2223
rect 2781 2189 2786 2223
rect 2786 2189 2815 2223
rect 2853 2189 2854 2223
rect 2854 2189 2887 2223
rect 2925 2189 2956 2223
rect 2956 2189 2959 2223
rect 3219 2189 3228 2223
rect 3228 2189 3253 2223
rect 3291 2189 3296 2223
rect 3296 2189 3325 2223
rect 3363 2189 3364 2223
rect 3364 2189 3397 2223
rect 3435 2189 3466 2223
rect 3466 2189 3469 2223
rect 3507 2189 3534 2223
rect 3534 2189 3541 2223
rect 3579 2189 3602 2223
rect 3602 2189 3613 2223
rect 3993 2189 4010 2223
rect 4010 2189 4027 2223
rect 4065 2189 4078 2223
rect 4078 2189 4099 2223
rect 4137 2189 4146 2223
rect 4146 2189 4171 2223
rect 4488 2189 4520 2223
rect 4520 2189 4522 2223
rect 4560 2189 4588 2223
rect 4588 2189 4594 2223
rect 4632 2189 4656 2223
rect 4656 2189 4666 2223
rect 4882 2189 4894 2223
rect 4894 2189 4916 2223
rect 4954 2189 4962 2223
rect 4962 2189 4988 2223
rect 5026 2189 5030 2223
rect 5030 2189 5060 2223
rect 5347 2189 5370 2223
rect 5370 2189 5381 2223
rect 5419 2189 5438 2223
rect 5438 2189 5453 2223
rect 5491 2189 5506 2223
rect 5506 2189 5525 2223
rect 5741 2189 5744 2223
rect 5744 2189 5775 2223
rect 5813 2189 5846 2223
rect 5846 2189 5847 2223
rect 5885 2189 5914 2223
rect 5914 2189 5919 2223
rect 6211 2189 6220 2223
rect 6220 2189 6245 2223
rect 6283 2189 6288 2223
rect 6288 2189 6317 2223
rect 6355 2189 6356 2223
rect 6356 2189 6389 2223
rect 6629 2189 6662 2223
rect 6662 2189 6663 2223
rect 6701 2189 6730 2223
rect 6730 2189 6735 2223
rect 6773 2189 6798 2223
rect 6798 2189 6807 2223
rect 6845 2189 6866 2223
rect 6866 2189 6879 2223
rect 6917 2189 6934 2223
rect 6934 2189 6951 2223
rect 6989 2189 7002 2223
rect 7002 2189 7023 2223
rect 7061 2189 7070 2223
rect 7070 2189 7095 2223
rect 7133 2189 7138 2223
rect 7138 2189 7167 2223
rect 7205 2189 7206 2223
rect 7206 2189 7239 2223
rect 7277 2189 7308 2223
rect 7308 2189 7311 2223
rect 7349 2189 7376 2223
rect 7376 2189 7383 2223
rect 7421 2189 7444 2223
rect 7444 2189 7455 2223
rect 7493 2189 7512 2223
rect 7512 2189 7527 2223
rect 7565 2189 7580 2223
rect 7580 2189 7599 2223
rect 7637 2189 7648 2223
rect 7648 2189 7671 2223
rect 7709 2189 7716 2223
rect 7716 2189 7743 2223
rect 7781 2189 7784 2223
rect 7784 2189 7815 2223
rect 7853 2189 7886 2223
rect 7886 2189 7887 2223
rect 7925 2189 7954 2223
rect 7954 2189 7959 2223
rect 7997 2189 8022 2223
rect 8022 2189 8031 2223
rect 8069 2189 8090 2223
rect 8090 2189 8103 2223
rect 8141 2189 8158 2223
rect 8158 2189 8175 2223
rect 8213 2189 8226 2223
rect 8226 2189 8247 2223
rect 8285 2189 8294 2223
rect 8294 2189 8319 2223
rect 8357 2189 8362 2223
rect 8362 2189 8391 2223
rect 8429 2189 8430 2223
rect 8430 2189 8463 2223
rect 8501 2189 8532 2223
rect 8532 2189 8535 2223
rect 8573 2189 8600 2223
rect 8600 2189 8607 2223
rect 8645 2189 8668 2223
rect 8668 2189 8679 2223
rect 8717 2189 8736 2223
rect 8736 2189 8751 2223
rect 8789 2189 8804 2223
rect 8804 2189 8823 2223
rect 8861 2189 8872 2223
rect 8872 2189 8895 2223
rect 8933 2189 8940 2223
rect 8940 2189 8967 2223
rect 9005 2189 9008 2223
rect 9008 2189 9039 2223
rect 9077 2189 9110 2223
rect 9110 2189 9111 2223
rect 9149 2189 9178 2223
rect 9178 2189 9183 2223
rect 9221 2189 9246 2223
rect 9246 2189 9255 2223
rect 9293 2189 9314 2223
rect 9314 2189 9327 2223
rect 9365 2189 9382 2223
rect 9382 2189 9399 2223
rect 9437 2189 9450 2223
rect 9450 2189 9471 2223
rect 9509 2189 9518 2223
rect 9518 2189 9543 2223
rect 9581 2189 9586 2223
rect 9586 2189 9615 2223
rect 9653 2189 9654 2223
rect 9654 2189 9687 2223
rect 9725 2189 9756 2223
rect 9756 2189 9759 2223
rect 9797 2189 9824 2223
rect 9824 2189 9831 2223
rect 9869 2189 9892 2223
rect 9892 2189 9903 2223
rect 9941 2189 9960 2223
rect 9960 2189 9975 2223
rect 10013 2189 10028 2223
rect 10028 2189 10047 2223
rect 10085 2189 10096 2223
rect 10096 2189 10119 2223
rect 10157 2189 10164 2223
rect 10164 2189 10191 2223
rect 10229 2189 10232 2223
rect 10232 2189 10263 2223
rect 10301 2189 10334 2223
rect 10334 2189 10335 2223
rect 10373 2189 10402 2223
rect 10402 2189 10407 2223
rect 10445 2189 10470 2223
rect 10470 2189 10479 2223
rect 10517 2189 10538 2223
rect 10538 2189 10551 2223
rect 10589 2189 10606 2223
rect 10606 2189 10623 2223
rect 10661 2189 10674 2223
rect 10674 2189 10695 2223
rect 10733 2189 10742 2223
rect 10742 2189 10767 2223
rect 10805 2189 10810 2223
rect 10810 2189 10839 2223
rect 10877 2189 10878 2223
rect 10878 2189 10911 2223
rect 11506 3916 11540 3950
rect 15405 4000 15438 4016
rect 15438 4000 15439 4016
rect 15484 4000 15508 4012
rect 15508 4000 15518 4012
rect 15560 4000 15578 4012
rect 15578 4000 15594 4012
rect 15636 4000 15648 4012
rect 15648 4000 15670 4012
rect 15733 4016 15754 4034
rect 15754 4016 15767 4034
rect 15819 4016 15824 4034
rect 15824 4016 15853 4034
rect 15905 4016 15928 4034
rect 15928 4016 15939 4034
rect 15991 4016 15998 4034
rect 15998 4016 16025 4034
rect 15405 3982 15439 4000
rect 15484 3978 15518 4000
rect 15560 3978 15594 4000
rect 15636 3978 15670 4000
rect 15733 3966 15767 3978
rect 15819 3966 15853 3978
rect 15905 3966 15939 3978
rect 15991 3966 16025 3978
rect 15733 3944 15754 3966
rect 15754 3944 15767 3966
rect 15819 3944 15824 3966
rect 15824 3944 15853 3966
rect 15905 3944 15928 3966
rect 15928 3944 15939 3966
rect 15991 3944 15998 3966
rect 15998 3944 16025 3966
rect 11506 3847 11540 3878
rect 11506 3844 11540 3847
rect 11624 3874 11626 3908
rect 11626 3874 11658 3908
rect 11696 3874 11728 3908
rect 11728 3874 11730 3908
rect 14526 3874 14528 3908
rect 14528 3874 14560 3908
rect 14598 3874 14630 3908
rect 14630 3874 14632 3908
rect 15484 3898 15518 3932
rect 15560 3898 15594 3932
rect 15636 3898 15670 3932
rect 15733 3898 15767 3906
rect 15819 3898 15853 3906
rect 15905 3898 15939 3906
rect 15991 3898 16025 3906
rect 15733 3872 15754 3898
rect 15754 3872 15767 3898
rect 15819 3872 15824 3898
rect 15824 3872 15853 3898
rect 15905 3872 15928 3898
rect 15928 3872 15939 3898
rect 15991 3872 15998 3898
rect 15998 3872 16025 3898
rect 11506 3778 11540 3806
rect 11506 3772 11540 3778
rect 15554 3830 15588 3859
rect 15626 3830 15660 3859
rect 15733 3830 15767 3834
rect 15819 3830 15853 3834
rect 15905 3830 15939 3834
rect 15991 3830 16025 3834
rect 15554 3825 15578 3830
rect 15578 3825 15588 3830
rect 15626 3825 15648 3830
rect 15648 3825 15660 3830
rect 15733 3800 15754 3830
rect 15754 3800 15767 3830
rect 15819 3800 15824 3830
rect 15824 3800 15853 3830
rect 15905 3800 15928 3830
rect 15928 3800 15939 3830
rect 15991 3800 15998 3830
rect 15998 3800 16025 3830
rect 11506 3709 11540 3734
rect 11506 3700 11540 3709
rect 11624 3720 11626 3754
rect 11626 3720 11658 3754
rect 11696 3720 11728 3754
rect 11728 3720 11730 3754
rect 14526 3720 14528 3754
rect 14528 3720 14560 3754
rect 14598 3720 14630 3754
rect 14630 3720 14632 3754
rect 15733 3728 15754 3762
rect 15754 3728 15767 3762
rect 15819 3728 15824 3762
rect 15824 3728 15853 3762
rect 15905 3728 15928 3762
rect 15928 3728 15939 3762
rect 15991 3728 15998 3762
rect 15998 3728 16025 3762
rect 11506 3640 11540 3662
rect 11506 3628 11540 3640
rect 15733 3660 15754 3690
rect 15754 3660 15767 3690
rect 15819 3660 15824 3690
rect 15824 3660 15853 3690
rect 15905 3660 15928 3690
rect 15928 3660 15939 3690
rect 15991 3660 15998 3690
rect 15998 3660 16025 3690
rect 15733 3656 15767 3660
rect 15819 3656 15853 3660
rect 15905 3656 15939 3660
rect 15991 3656 16025 3660
rect 11506 3571 11540 3590
rect 11506 3556 11540 3571
rect 11624 3566 11626 3600
rect 11626 3566 11658 3600
rect 11696 3566 11728 3600
rect 11728 3566 11730 3600
rect 14526 3566 14528 3600
rect 14528 3566 14560 3600
rect 14598 3566 14630 3600
rect 14630 3566 14632 3600
rect 15733 3592 15754 3618
rect 15754 3592 15767 3618
rect 15819 3592 15824 3618
rect 15824 3592 15853 3618
rect 15905 3592 15928 3618
rect 15928 3592 15939 3618
rect 15991 3592 15998 3618
rect 15998 3592 16025 3618
rect 15733 3584 15767 3592
rect 15819 3584 15853 3592
rect 15905 3584 15939 3592
rect 15991 3584 16025 3592
rect 11506 3502 11540 3518
rect 11506 3484 11540 3502
rect 11506 3433 11540 3446
rect 11506 3412 11540 3433
rect 15733 3524 15754 3546
rect 15754 3524 15767 3546
rect 15819 3524 15824 3546
rect 15824 3524 15853 3546
rect 15905 3524 15928 3546
rect 15928 3524 15939 3546
rect 15991 3524 15998 3546
rect 15998 3524 16025 3546
rect 15733 3512 15767 3524
rect 15819 3512 15853 3524
rect 15905 3512 15939 3524
rect 15991 3512 16025 3524
rect 15733 3456 15754 3474
rect 15754 3456 15767 3474
rect 15819 3456 15824 3474
rect 15824 3456 15853 3474
rect 15905 3456 15928 3474
rect 15928 3456 15939 3474
rect 15991 3456 15998 3474
rect 15998 3456 16025 3474
rect 11624 3412 11626 3446
rect 11626 3412 11658 3446
rect 11696 3412 11728 3446
rect 11728 3412 11730 3446
rect 14526 3412 14528 3446
rect 14528 3412 14560 3446
rect 14598 3412 14630 3446
rect 14630 3412 14632 3446
rect 15733 3440 15767 3456
rect 15819 3440 15853 3456
rect 15905 3440 15939 3456
rect 15991 3440 16025 3456
rect 11506 3364 11540 3374
rect 11506 3340 11540 3364
rect 11506 3295 11540 3302
rect 11506 3268 11540 3295
rect 15733 3388 15754 3402
rect 15754 3388 15767 3402
rect 15819 3388 15824 3402
rect 15824 3388 15853 3402
rect 15905 3388 15928 3402
rect 15928 3388 15939 3402
rect 15991 3388 15998 3402
rect 15998 3388 16025 3402
rect 15733 3368 15767 3388
rect 15819 3368 15853 3388
rect 15905 3368 15939 3388
rect 15991 3368 16025 3388
rect 15733 3320 15754 3330
rect 15754 3320 15767 3330
rect 15819 3320 15824 3330
rect 15824 3320 15853 3330
rect 15905 3320 15928 3330
rect 15928 3320 15939 3330
rect 15991 3320 15998 3330
rect 15998 3320 16025 3330
rect 15733 3296 15767 3320
rect 15819 3296 15853 3320
rect 15905 3296 15939 3320
rect 15991 3296 16025 3320
rect 11506 3226 11540 3230
rect 11506 3196 11540 3226
rect 11624 3258 11626 3292
rect 11626 3258 11658 3292
rect 11696 3258 11728 3292
rect 11728 3258 11730 3292
rect 14526 3258 14528 3292
rect 14528 3258 14560 3292
rect 14598 3258 14630 3292
rect 14630 3258 14632 3292
rect 15733 3252 15754 3258
rect 15754 3252 15767 3258
rect 15819 3252 15824 3258
rect 15824 3252 15853 3258
rect 15905 3252 15928 3258
rect 15928 3252 15939 3258
rect 15991 3252 15998 3258
rect 15998 3252 16025 3258
rect 11506 3157 11540 3158
rect 11506 3124 11540 3157
rect 15733 3224 15767 3252
rect 15819 3224 15853 3252
rect 15905 3224 15939 3252
rect 15991 3224 16025 3252
rect 15733 3184 15754 3186
rect 15754 3184 15767 3186
rect 15819 3184 15824 3186
rect 15824 3184 15853 3186
rect 15905 3184 15928 3186
rect 15928 3184 15939 3186
rect 15991 3184 15998 3186
rect 15998 3184 16025 3186
rect 15733 3152 15767 3184
rect 15819 3152 15853 3184
rect 15905 3152 15939 3184
rect 15991 3152 16025 3184
rect 11624 3104 11626 3138
rect 11626 3104 11658 3138
rect 11696 3104 11728 3138
rect 11728 3104 11730 3138
rect 14526 3104 14528 3138
rect 14528 3104 14560 3138
rect 14598 3104 14630 3138
rect 14630 3104 14632 3138
rect 11506 3053 11540 3086
rect 11506 3052 11540 3053
rect 11506 2984 11540 3014
rect 11506 2980 11540 2984
rect 15733 3082 15767 3114
rect 15819 3082 15853 3114
rect 15905 3082 15939 3114
rect 15991 3082 16025 3114
rect 15733 3080 15754 3082
rect 15754 3080 15767 3082
rect 15819 3080 15824 3082
rect 15824 3080 15853 3082
rect 15905 3080 15928 3082
rect 15928 3080 15939 3082
rect 15991 3080 15998 3082
rect 15998 3080 16025 3082
rect 15733 3014 15767 3042
rect 15819 3014 15853 3042
rect 15905 3014 15939 3042
rect 15991 3014 16025 3042
rect 11624 2950 11626 2984
rect 11626 2950 11658 2984
rect 11696 2950 11728 2984
rect 11728 2950 11730 2984
rect 14526 2950 14528 2984
rect 14528 2950 14560 2984
rect 14598 2950 14630 2984
rect 14630 2950 14632 2984
rect 15733 3008 15754 3014
rect 15754 3008 15767 3014
rect 15819 3008 15824 3014
rect 15824 3008 15853 3014
rect 15905 3008 15928 3014
rect 15928 3008 15939 3014
rect 15991 3008 15998 3014
rect 15998 3008 16025 3014
rect 11506 2915 11540 2942
rect 11506 2908 11540 2915
rect 15733 2946 15767 2970
rect 15819 2946 15853 2970
rect 15905 2946 15939 2970
rect 15991 2946 16025 2970
rect 11506 2846 11540 2870
rect 11506 2836 11540 2846
rect 15733 2936 15754 2946
rect 15754 2936 15767 2946
rect 15819 2936 15824 2946
rect 15824 2936 15853 2946
rect 15905 2936 15928 2946
rect 15928 2936 15939 2946
rect 15991 2936 15998 2946
rect 15998 2936 16025 2946
rect 15733 2878 15767 2898
rect 15819 2878 15853 2898
rect 15905 2878 15939 2898
rect 15991 2878 16025 2898
rect 15733 2864 15754 2878
rect 15754 2864 15767 2878
rect 15819 2864 15824 2878
rect 15824 2864 15853 2878
rect 15905 2864 15928 2878
rect 15928 2864 15939 2878
rect 15991 2864 15998 2878
rect 15998 2864 16025 2878
rect 11506 2777 11540 2798
rect 11506 2764 11540 2777
rect 11624 2796 11626 2830
rect 11626 2796 11658 2830
rect 11696 2796 11728 2830
rect 11728 2796 11730 2830
rect 14526 2796 14528 2830
rect 14528 2796 14560 2830
rect 14598 2796 14630 2830
rect 14630 2796 14632 2830
rect 15733 2810 15767 2826
rect 15819 2810 15853 2826
rect 15905 2810 15939 2826
rect 15991 2810 16025 2826
rect 11506 2708 11540 2726
rect 11506 2692 11540 2708
rect 15733 2792 15754 2810
rect 15754 2792 15767 2810
rect 15819 2792 15824 2810
rect 15824 2792 15853 2810
rect 15905 2792 15928 2810
rect 15928 2792 15939 2810
rect 15991 2792 15998 2810
rect 15998 2792 16025 2810
rect 15733 2742 15767 2754
rect 15819 2742 15853 2754
rect 15905 2742 15939 2754
rect 15991 2742 16025 2754
rect 15733 2720 15754 2742
rect 15754 2720 15767 2742
rect 15819 2720 15824 2742
rect 15824 2720 15853 2742
rect 15905 2720 15928 2742
rect 15928 2720 15939 2742
rect 15991 2720 15998 2742
rect 15998 2720 16025 2742
rect 11506 2639 11540 2654
rect 11506 2620 11540 2639
rect 11624 2642 11626 2676
rect 11626 2642 11658 2676
rect 11696 2642 11728 2676
rect 11728 2642 11730 2676
rect 14526 2642 14528 2676
rect 14528 2642 14560 2676
rect 14598 2642 14630 2676
rect 14630 2642 14632 2676
rect 15733 2674 15767 2681
rect 15819 2674 15853 2681
rect 15905 2674 15939 2681
rect 15991 2674 16025 2681
rect 15733 2647 15754 2674
rect 15754 2647 15767 2674
rect 15819 2647 15824 2674
rect 15824 2647 15853 2674
rect 15905 2647 15928 2674
rect 15928 2647 15939 2674
rect 15991 2647 15998 2674
rect 15998 2647 16025 2674
rect 11506 2570 11540 2582
rect 11506 2548 11540 2570
rect 15733 2606 15767 2608
rect 15819 2606 15853 2608
rect 15905 2606 15939 2608
rect 15991 2606 16025 2608
rect 15733 2574 15754 2606
rect 15754 2574 15767 2606
rect 15819 2574 15824 2606
rect 15824 2574 15853 2606
rect 15905 2574 15928 2606
rect 15928 2574 15939 2606
rect 15991 2574 15998 2606
rect 15998 2574 16025 2606
rect 11506 2501 11540 2510
rect 11506 2476 11540 2501
rect 11624 2488 11626 2522
rect 11626 2488 11658 2522
rect 11696 2488 11728 2522
rect 11728 2488 11730 2522
rect 14526 2488 14528 2522
rect 14528 2488 14560 2522
rect 14598 2488 14630 2522
rect 14630 2488 14632 2522
rect 15733 2504 15754 2535
rect 15754 2504 15767 2535
rect 15819 2504 15824 2535
rect 15824 2504 15853 2535
rect 15905 2504 15928 2535
rect 15928 2504 15939 2535
rect 15991 2504 15998 2535
rect 15998 2504 16025 2535
rect 15733 2501 15767 2504
rect 15819 2501 15853 2504
rect 15905 2501 15939 2504
rect 15991 2501 16025 2504
rect 11506 2431 11540 2438
rect 11506 2404 11540 2431
rect 15733 2436 15754 2462
rect 15754 2436 15767 2462
rect 15819 2436 15824 2462
rect 15824 2436 15853 2462
rect 15905 2436 15928 2462
rect 15928 2436 15939 2462
rect 15991 2436 15998 2462
rect 15998 2436 16025 2462
rect 15733 2428 15767 2436
rect 15819 2428 15853 2436
rect 15905 2428 15939 2436
rect 15991 2428 16025 2436
rect 15733 2368 15754 2389
rect 15754 2368 15767 2389
rect 15819 2368 15824 2389
rect 15824 2368 15853 2389
rect 15905 2368 15928 2389
rect 15928 2368 15939 2389
rect 15991 2368 15998 2389
rect 15998 2368 16025 2389
rect 11506 2361 11540 2366
rect 11506 2332 11540 2361
rect 11624 2334 11626 2368
rect 11626 2334 11658 2368
rect 11696 2334 11728 2368
rect 11728 2334 11730 2368
rect 14526 2334 14528 2368
rect 14528 2334 14560 2368
rect 14598 2334 14630 2368
rect 14630 2334 14632 2368
rect 15733 2355 15767 2368
rect 15819 2355 15853 2368
rect 15905 2355 15939 2368
rect 15991 2355 16025 2368
rect 11506 2291 11540 2294
rect 11506 2260 11540 2291
rect 15733 2300 15754 2316
rect 15754 2300 15767 2316
rect 15819 2300 15824 2316
rect 15824 2300 15853 2316
rect 15905 2300 15928 2316
rect 15928 2300 15939 2316
rect 15991 2300 15998 2316
rect 15998 2300 16025 2316
rect 15733 2282 15767 2300
rect 15819 2282 15853 2300
rect 15905 2282 15939 2300
rect 15991 2282 16025 2300
rect 15733 2232 15754 2243
rect 15754 2232 15767 2243
rect 15819 2232 15824 2243
rect 15824 2232 15853 2243
rect 15905 2232 15928 2243
rect 15928 2232 15939 2243
rect 15991 2232 15998 2243
rect 15998 2232 16025 2243
rect 11506 2221 11540 2222
rect 11506 2188 11540 2221
rect 11624 2180 11626 2214
rect 11626 2180 11658 2214
rect 11696 2180 11728 2214
rect 11728 2180 11730 2214
rect 14526 2180 14528 2214
rect 14528 2180 14560 2214
rect 14598 2180 14630 2214
rect 14630 2180 14632 2214
rect 15733 2209 15767 2232
rect 15819 2209 15853 2232
rect 15905 2209 15939 2232
rect 15991 2209 16025 2232
rect 15733 2164 15754 2170
rect 15754 2164 15767 2170
rect 15819 2164 15824 2170
rect 15824 2164 15853 2170
rect 15905 2164 15928 2170
rect 15928 2164 15939 2170
rect 15991 2164 15998 2170
rect 15998 2164 16025 2170
rect 6625 2110 6659 2144
rect 6698 2110 6732 2144
rect 6771 2110 6805 2144
rect 6844 2110 6878 2144
rect 6917 2110 6951 2144
rect 6990 2110 7024 2144
rect 7063 2110 7097 2144
rect 7136 2110 7170 2144
rect 7209 2110 7243 2144
rect 7282 2110 7316 2144
rect 7355 2110 7389 2144
rect 7428 2110 7462 2144
rect 7501 2110 7535 2144
rect 7574 2110 7608 2144
rect 7647 2110 7681 2144
rect 7720 2110 7754 2144
rect 7792 2110 7826 2144
rect 7864 2110 7898 2144
rect 7936 2110 7970 2144
rect 8008 2110 8042 2144
rect 8080 2110 8114 2144
rect 8152 2110 8186 2144
rect 8224 2110 8258 2144
rect 8296 2110 8330 2144
rect 8368 2110 8402 2144
rect 8440 2110 8474 2144
rect 8512 2110 8546 2144
rect 8584 2110 8618 2144
rect 8656 2110 8690 2144
rect 8728 2110 8762 2144
rect 8800 2110 8834 2144
rect 8872 2110 8906 2144
rect 8944 2110 8978 2144
rect 9016 2110 9050 2144
rect 9088 2110 9122 2144
rect 9160 2110 9194 2144
rect 9232 2110 9266 2144
rect 9304 2110 9338 2144
rect 9376 2110 9410 2144
rect 9448 2110 9482 2144
rect 9520 2110 9554 2144
rect 9592 2110 9626 2144
rect 9664 2110 9698 2144
rect 9736 2110 9770 2144
rect 9808 2110 9842 2144
rect 9880 2110 9914 2144
rect 9952 2110 9986 2144
rect 10024 2110 10058 2144
rect 10096 2110 10130 2144
rect 10168 2110 10202 2144
rect 10240 2110 10274 2144
rect 10312 2110 10346 2144
rect 10384 2110 10418 2144
rect 10456 2110 10490 2144
rect 10528 2110 10562 2144
rect 10600 2110 10634 2144
rect 10672 2110 10706 2144
rect 10744 2110 10778 2144
rect 10816 2110 10850 2144
rect 10888 2110 10922 2144
rect 11506 2117 11540 2150
rect 11506 2116 11540 2117
rect 15733 2136 15767 2164
rect 15819 2136 15853 2164
rect 15905 2136 15939 2164
rect 15991 2136 16025 2164
rect 15733 2096 15754 2097
rect 15754 2096 15767 2097
rect 15819 2096 15824 2097
rect 15824 2096 15853 2097
rect 15905 2096 15928 2097
rect 15928 2096 15939 2097
rect 15991 2096 15998 2097
rect 15998 2096 16025 2097
rect 11506 2069 11540 2078
rect 360 2035 370 2060
rect 370 2035 394 2060
rect 449 2035 474 2069
rect 474 2035 483 2069
rect 521 2035 543 2069
rect 543 2035 555 2069
rect 593 2035 612 2069
rect 612 2035 627 2069
rect 665 2035 681 2069
rect 681 2035 699 2069
rect 1069 2035 1095 2069
rect 1095 2035 1103 2069
rect 1141 2035 1164 2069
rect 1164 2035 1175 2069
rect 1213 2035 1233 2069
rect 1233 2035 1247 2069
rect 1458 2035 1474 2069
rect 1474 2035 1492 2069
rect 1530 2035 1543 2069
rect 1543 2035 1564 2069
rect 1602 2035 1612 2069
rect 1612 2035 1636 2069
rect 1912 2035 1923 2069
rect 1923 2035 1946 2069
rect 1984 2035 1992 2069
rect 1992 2035 2018 2069
rect 2056 2035 2061 2069
rect 2061 2035 2090 2069
rect 2317 2035 2337 2069
rect 2337 2035 2351 2069
rect 2389 2035 2406 2069
rect 2406 2035 2423 2069
rect 2461 2035 2475 2069
rect 2475 2035 2495 2069
rect 2781 2035 2785 2069
rect 2785 2035 2815 2069
rect 2853 2035 2854 2069
rect 2854 2035 2887 2069
rect 2925 2035 2958 2069
rect 2958 2035 2959 2069
rect 3219 2035 3234 2069
rect 3234 2035 3253 2069
rect 3291 2035 3303 2069
rect 3303 2035 3325 2069
rect 3363 2035 3372 2069
rect 3372 2035 3397 2069
rect 3435 2035 3441 2069
rect 3441 2035 3469 2069
rect 3507 2035 3510 2069
rect 3510 2035 3541 2069
rect 3579 2035 3613 2069
rect 3993 2035 4027 2069
rect 4065 2035 4096 2069
rect 4096 2035 4099 2069
rect 4137 2035 4165 2069
rect 4165 2035 4171 2069
rect 4488 2035 4509 2069
rect 4509 2035 4522 2069
rect 4560 2035 4577 2069
rect 4577 2035 4594 2069
rect 4632 2035 4645 2069
rect 4645 2035 4666 2069
rect 4882 2035 4883 2069
rect 4883 2035 4916 2069
rect 4954 2035 4985 2069
rect 4985 2035 4988 2069
rect 5026 2035 5053 2069
rect 5053 2035 5060 2069
rect 5347 2035 5359 2069
rect 5359 2035 5381 2069
rect 5419 2035 5427 2069
rect 5427 2035 5453 2069
rect 5491 2035 5495 2069
rect 5495 2035 5525 2069
rect 5741 2035 5767 2069
rect 5767 2035 5775 2069
rect 5813 2035 5835 2069
rect 5835 2035 5847 2069
rect 5885 2035 5903 2069
rect 5903 2035 5919 2069
rect 6211 2035 6243 2069
rect 6243 2035 6245 2069
rect 6283 2035 6311 2069
rect 6311 2035 6317 2069
rect 6355 2035 6379 2069
rect 6379 2035 6389 2069
rect 6629 2035 6651 2069
rect 6651 2035 6663 2069
rect 6701 2035 6719 2069
rect 6719 2035 6735 2069
rect 6773 2035 6787 2069
rect 6787 2035 6807 2069
rect 6845 2035 6855 2069
rect 6855 2035 6879 2069
rect 6917 2035 6923 2069
rect 6923 2035 6951 2069
rect 6989 2035 6991 2069
rect 6991 2035 7023 2069
rect 7061 2035 7093 2069
rect 7093 2035 7095 2069
rect 7133 2035 7161 2069
rect 7161 2035 7167 2069
rect 7205 2035 7229 2069
rect 7229 2035 7239 2069
rect 7277 2035 7297 2069
rect 7297 2035 7311 2069
rect 7349 2035 7365 2069
rect 7365 2035 7383 2069
rect 7421 2035 7433 2069
rect 7433 2035 7455 2069
rect 7493 2035 7501 2069
rect 7501 2035 7527 2069
rect 7565 2035 7569 2069
rect 7569 2035 7599 2069
rect 7637 2035 7671 2069
rect 7709 2035 7739 2069
rect 7739 2035 7743 2069
rect 7781 2035 7807 2069
rect 7807 2035 7815 2069
rect 7853 2035 7875 2069
rect 7875 2035 7887 2069
rect 7925 2035 7943 2069
rect 7943 2035 7959 2069
rect 7997 2035 8011 2069
rect 8011 2035 8031 2069
rect 8069 2035 8079 2069
rect 8079 2035 8103 2069
rect 8141 2035 8147 2069
rect 8147 2035 8175 2069
rect 8213 2035 8215 2069
rect 8215 2035 8247 2069
rect 8285 2035 8317 2069
rect 8317 2035 8319 2069
rect 8357 2035 8385 2069
rect 8385 2035 8391 2069
rect 8429 2035 8453 2069
rect 8453 2035 8463 2069
rect 8501 2035 8521 2069
rect 8521 2035 8535 2069
rect 8573 2035 8589 2069
rect 8589 2035 8607 2069
rect 8645 2035 8657 2069
rect 8657 2035 8679 2069
rect 8717 2035 8725 2069
rect 8725 2035 8751 2069
rect 8789 2035 8793 2069
rect 8793 2035 8823 2069
rect 8861 2035 8895 2069
rect 8933 2035 8963 2069
rect 8963 2035 8967 2069
rect 9005 2035 9031 2069
rect 9031 2035 9039 2069
rect 9077 2035 9099 2069
rect 9099 2035 9111 2069
rect 9149 2035 9167 2069
rect 9167 2035 9183 2069
rect 9221 2035 9235 2069
rect 9235 2035 9255 2069
rect 9293 2035 9303 2069
rect 9303 2035 9327 2069
rect 9365 2035 9371 2069
rect 9371 2035 9399 2069
rect 9437 2035 9439 2069
rect 9439 2035 9471 2069
rect 9509 2035 9541 2069
rect 9541 2035 9543 2069
rect 9581 2035 9609 2069
rect 9609 2035 9615 2069
rect 9653 2035 9677 2069
rect 9677 2035 9687 2069
rect 9725 2035 9745 2069
rect 9745 2035 9759 2069
rect 9797 2035 9813 2069
rect 9813 2035 9831 2069
rect 9869 2035 9881 2069
rect 9881 2035 9903 2069
rect 9941 2035 9949 2069
rect 9949 2035 9975 2069
rect 10013 2035 10017 2069
rect 10017 2035 10047 2069
rect 10085 2035 10119 2069
rect 10157 2035 10187 2069
rect 10187 2035 10191 2069
rect 10229 2035 10255 2069
rect 10255 2035 10263 2069
rect 10301 2035 10323 2069
rect 10323 2035 10335 2069
rect 10373 2035 10391 2069
rect 10391 2035 10407 2069
rect 10445 2035 10459 2069
rect 10459 2035 10479 2069
rect 10517 2035 10527 2069
rect 10527 2035 10551 2069
rect 10589 2035 10595 2069
rect 10595 2035 10623 2069
rect 10661 2035 10663 2069
rect 10663 2035 10695 2069
rect 10733 2035 10765 2069
rect 10765 2035 10767 2069
rect 10805 2035 10833 2069
rect 10833 2035 10839 2069
rect 10877 2035 10901 2069
rect 10901 2035 10911 2069
rect 11506 2044 11513 2069
rect 11513 2044 11540 2069
rect 11608 2035 11615 2069
rect 11615 2035 11642 2069
rect 11680 2035 11683 2069
rect 11683 2035 11714 2069
rect 11752 2035 11785 2069
rect 11785 2035 11786 2069
rect 11824 2035 11853 2069
rect 11853 2035 11858 2069
rect 11896 2035 11921 2069
rect 11921 2035 11930 2069
rect 11968 2035 11989 2069
rect 11989 2035 12002 2069
rect 12040 2035 12057 2069
rect 12057 2035 12074 2069
rect 12112 2035 12125 2069
rect 12125 2035 12146 2069
rect 12184 2035 12193 2069
rect 12193 2035 12218 2069
rect 12256 2035 12261 2069
rect 12261 2035 12290 2069
rect 12328 2035 12329 2069
rect 12329 2035 12362 2069
rect 12400 2035 12431 2069
rect 12431 2035 12434 2069
rect 12472 2035 12499 2069
rect 12499 2035 12506 2069
rect 12544 2035 12567 2069
rect 12567 2035 12578 2069
rect 12616 2035 12635 2069
rect 12635 2035 12650 2069
rect 12688 2035 12703 2069
rect 12703 2035 12722 2069
rect 12760 2035 12771 2069
rect 12771 2035 12794 2069
rect 12832 2035 12839 2069
rect 12839 2035 12866 2069
rect 12904 2035 12907 2069
rect 12907 2035 12938 2069
rect 12976 2035 13009 2069
rect 13009 2035 13010 2069
rect 13048 2035 13077 2069
rect 13077 2035 13082 2069
rect 13120 2035 13145 2069
rect 13145 2035 13154 2069
rect 13192 2035 13213 2069
rect 13213 2035 13226 2069
rect 13264 2035 13281 2069
rect 13281 2035 13298 2069
rect 13336 2035 13349 2069
rect 13349 2035 13370 2069
rect 13408 2035 13417 2069
rect 13417 2035 13442 2069
rect 13480 2035 13485 2069
rect 13485 2035 13514 2069
rect 13552 2035 13553 2069
rect 13553 2035 13586 2069
rect 13624 2035 13655 2069
rect 13655 2035 13658 2069
rect 13696 2035 13723 2069
rect 13723 2035 13730 2069
rect 13768 2035 13791 2069
rect 13791 2035 13802 2069
rect 13840 2035 13859 2069
rect 13859 2035 13874 2069
rect 13912 2035 13927 2069
rect 13927 2035 13946 2069
rect 13984 2035 13995 2069
rect 13995 2035 14018 2069
rect 14056 2035 14063 2069
rect 14063 2035 14090 2069
rect 14128 2035 14131 2069
rect 14131 2035 14162 2069
rect 14200 2035 14233 2069
rect 14233 2035 14234 2069
rect 14272 2035 14301 2069
rect 14301 2035 14306 2069
rect 14344 2035 14369 2069
rect 14369 2035 14378 2069
rect 14416 2035 14437 2069
rect 14437 2035 14450 2069
rect 14488 2035 14505 2069
rect 14505 2035 14522 2069
rect 14560 2035 14573 2069
rect 14573 2035 14594 2069
rect 14632 2035 14641 2069
rect 14641 2035 14666 2069
rect 14704 2035 14709 2069
rect 14709 2035 14738 2069
rect 15733 2063 15767 2096
rect 15819 2063 15853 2096
rect 15905 2063 15939 2096
rect 15991 2063 16025 2096
rect 360 2026 394 2035
rect 360 1959 394 1988
rect 360 1954 394 1959
rect 15733 1994 15767 2024
rect 15819 1994 15853 2024
rect 15905 1994 15939 2024
rect 15991 1994 16025 2024
rect 15733 1990 15754 1994
rect 15754 1990 15767 1994
rect 15819 1990 15824 1994
rect 15824 1990 15853 1994
rect 15905 1990 15928 1994
rect 15928 1990 15939 1994
rect 15991 1990 15998 1994
rect 15998 1990 16025 1994
rect 360 1889 394 1916
rect 360 1882 394 1889
rect 478 1890 480 1924
rect 480 1890 512 1924
rect 550 1890 582 1924
rect 582 1890 584 1924
rect 3380 1890 3382 1924
rect 3382 1890 3414 1924
rect 3452 1890 3484 1924
rect 3484 1890 3486 1924
rect 12882 1890 12884 1924
rect 12884 1890 12916 1924
rect 12954 1890 12986 1924
rect 12986 1890 12988 1924
rect 15733 1926 15767 1951
rect 15819 1926 15853 1951
rect 15905 1926 15939 1951
rect 15991 1926 16025 1951
rect 15733 1917 15754 1926
rect 15754 1917 15767 1926
rect 15819 1917 15824 1926
rect 15824 1917 15853 1926
rect 15905 1917 15928 1926
rect 15928 1917 15939 1926
rect 15991 1917 15998 1926
rect 15998 1917 16025 1926
rect 360 1819 394 1844
rect 360 1810 394 1819
rect 13168 1827 13194 1847
rect 13194 1827 13202 1847
rect 13244 1827 13264 1847
rect 13264 1827 13278 1847
rect 13320 1827 13334 1847
rect 13334 1827 13354 1847
rect 13396 1827 13404 1847
rect 13404 1827 13430 1847
rect 13472 1827 13474 1847
rect 13474 1827 13506 1847
rect 13548 1827 13578 1847
rect 13578 1827 13582 1847
rect 13624 1827 13648 1847
rect 13648 1827 13658 1847
rect 13700 1827 13718 1847
rect 13718 1827 13734 1847
rect 13776 1827 13788 1847
rect 13788 1827 13810 1847
rect 13851 1827 13858 1847
rect 13858 1827 13885 1847
rect 13926 1827 13928 1847
rect 13928 1827 13960 1847
rect 14001 1827 14034 1847
rect 14034 1827 14035 1847
rect 14076 1827 14104 1847
rect 14104 1827 14110 1847
rect 14151 1827 14174 1847
rect 14174 1827 14185 1847
rect 14226 1827 14244 1847
rect 14244 1827 14260 1847
rect 14301 1827 14314 1847
rect 14314 1827 14335 1847
rect 14376 1827 14384 1847
rect 14384 1827 14410 1847
rect 14451 1827 14454 1847
rect 14454 1827 14485 1847
rect 14526 1827 14558 1847
rect 14558 1827 14560 1847
rect 14601 1827 14628 1847
rect 14628 1827 14635 1847
rect 15733 1858 15767 1878
rect 15819 1858 15853 1878
rect 15905 1858 15939 1878
rect 15991 1858 16025 1878
rect 13168 1813 13202 1827
rect 13244 1813 13278 1827
rect 13320 1813 13354 1827
rect 13396 1813 13430 1827
rect 13472 1813 13506 1827
rect 13548 1813 13582 1827
rect 13624 1813 13658 1827
rect 13700 1813 13734 1827
rect 13776 1813 13810 1827
rect 13851 1813 13885 1827
rect 13926 1813 13960 1827
rect 14001 1813 14035 1827
rect 14076 1813 14110 1827
rect 14151 1813 14185 1827
rect 14226 1813 14260 1827
rect 14301 1813 14335 1827
rect 14376 1813 14410 1827
rect 14451 1813 14485 1827
rect 14526 1813 14560 1827
rect 14601 1813 14635 1827
rect 15733 1844 15754 1858
rect 15754 1844 15767 1858
rect 15819 1844 15824 1858
rect 15824 1844 15853 1858
rect 15905 1844 15928 1858
rect 15928 1844 15939 1858
rect 15991 1844 15998 1858
rect 15998 1844 16025 1858
rect 360 1749 394 1772
rect 360 1738 394 1749
rect 478 1736 480 1770
rect 480 1736 512 1770
rect 550 1736 582 1770
rect 582 1736 584 1770
rect 3380 1736 3382 1770
rect 3382 1736 3414 1770
rect 3452 1736 3484 1770
rect 3484 1736 3486 1770
rect 12882 1736 12884 1770
rect 12884 1736 12916 1770
rect 12954 1736 12986 1770
rect 12986 1736 12988 1770
rect 15733 1790 15767 1805
rect 15819 1790 15853 1805
rect 15905 1790 15939 1805
rect 15991 1790 16025 1805
rect 15733 1771 15754 1790
rect 15754 1771 15767 1790
rect 15819 1771 15824 1790
rect 15824 1771 15853 1790
rect 15905 1771 15928 1790
rect 15928 1771 15939 1790
rect 15991 1771 15998 1790
rect 15998 1771 16025 1790
rect 15733 1722 15767 1732
rect 15819 1722 15853 1732
rect 15905 1722 15939 1732
rect 15991 1722 16025 1732
rect 360 1679 394 1700
rect 360 1666 394 1679
rect 15733 1698 15754 1722
rect 15754 1698 15767 1722
rect 15819 1698 15824 1722
rect 15824 1698 15853 1722
rect 15905 1698 15928 1722
rect 15928 1698 15939 1722
rect 15991 1698 15998 1722
rect 15998 1698 16025 1722
rect 15733 1654 15767 1659
rect 15819 1654 15853 1659
rect 15905 1654 15939 1659
rect 15991 1654 16025 1659
rect 360 1609 394 1628
rect 360 1594 394 1609
rect 15733 1625 15754 1654
rect 15754 1625 15767 1654
rect 15819 1625 15824 1654
rect 15824 1625 15853 1654
rect 15905 1625 15928 1654
rect 15928 1625 15939 1654
rect 15991 1625 15998 1654
rect 15998 1625 16025 1654
rect 478 1582 480 1616
rect 480 1582 512 1616
rect 550 1582 582 1616
rect 582 1582 584 1616
rect 3380 1582 3382 1616
rect 3382 1582 3414 1616
rect 3452 1582 3484 1616
rect 3484 1582 3486 1616
rect 12882 1582 12884 1616
rect 12884 1582 12916 1616
rect 12954 1582 12986 1616
rect 12986 1582 12988 1616
rect 360 1539 394 1556
rect 360 1522 394 1539
rect 360 1469 394 1484
rect 360 1450 394 1469
rect 15733 1552 15754 1586
rect 15754 1552 15767 1586
rect 15819 1552 15824 1586
rect 15824 1552 15853 1586
rect 15905 1552 15928 1586
rect 15928 1552 15939 1586
rect 15991 1552 15998 1586
rect 15998 1552 16025 1586
rect 15733 1484 15754 1513
rect 15754 1484 15767 1513
rect 15819 1484 15824 1513
rect 15824 1484 15853 1513
rect 15905 1484 15928 1513
rect 15928 1484 15939 1513
rect 15991 1484 15998 1513
rect 15998 1484 16025 1513
rect 15733 1479 15767 1484
rect 15819 1479 15853 1484
rect 15905 1479 15939 1484
rect 15991 1479 16025 1484
rect 478 1428 480 1462
rect 480 1428 512 1462
rect 550 1428 582 1462
rect 582 1428 584 1462
rect 3380 1428 3382 1462
rect 3382 1428 3414 1462
rect 3452 1428 3484 1462
rect 3484 1428 3486 1462
rect 12882 1428 12884 1462
rect 12884 1428 12916 1462
rect 12954 1428 12986 1462
rect 12986 1428 12988 1462
rect 360 1399 394 1412
rect 360 1378 394 1399
rect 360 1329 394 1340
rect 360 1306 394 1329
rect 15733 1416 15754 1440
rect 15754 1416 15767 1440
rect 15819 1416 15824 1440
rect 15824 1416 15853 1440
rect 15905 1416 15928 1440
rect 15928 1416 15939 1440
rect 15991 1416 15998 1440
rect 15998 1416 16025 1440
rect 15733 1406 15767 1416
rect 15819 1406 15853 1416
rect 15905 1406 15939 1416
rect 15991 1406 16025 1416
rect 13168 1371 13202 1385
rect 13244 1371 13278 1385
rect 13320 1371 13354 1385
rect 13396 1371 13430 1385
rect 13472 1371 13506 1385
rect 13548 1371 13582 1385
rect 13624 1371 13658 1385
rect 13700 1371 13734 1385
rect 13776 1371 13810 1385
rect 13851 1371 13885 1385
rect 13926 1371 13960 1385
rect 14001 1371 14035 1385
rect 14076 1371 14110 1385
rect 14151 1371 14185 1385
rect 14226 1371 14260 1385
rect 14301 1371 14335 1385
rect 14376 1371 14410 1385
rect 14451 1371 14485 1385
rect 14526 1371 14560 1385
rect 14601 1371 14635 1385
rect 13168 1351 13194 1371
rect 13194 1351 13202 1371
rect 13244 1351 13264 1371
rect 13264 1351 13278 1371
rect 13320 1351 13334 1371
rect 13334 1351 13354 1371
rect 13396 1351 13404 1371
rect 13404 1351 13430 1371
rect 13472 1351 13474 1371
rect 13474 1351 13506 1371
rect 13548 1351 13578 1371
rect 13578 1351 13582 1371
rect 13624 1351 13648 1371
rect 13648 1351 13658 1371
rect 13700 1351 13718 1371
rect 13718 1351 13734 1371
rect 13776 1351 13788 1371
rect 13788 1351 13810 1371
rect 13851 1351 13858 1371
rect 13858 1351 13885 1371
rect 13926 1351 13928 1371
rect 13928 1351 13960 1371
rect 14001 1351 14034 1371
rect 14034 1351 14035 1371
rect 14076 1351 14104 1371
rect 14104 1351 14110 1371
rect 14151 1351 14174 1371
rect 14174 1351 14185 1371
rect 14226 1351 14244 1371
rect 14244 1351 14260 1371
rect 14301 1351 14314 1371
rect 14314 1351 14335 1371
rect 14376 1351 14384 1371
rect 14384 1351 14410 1371
rect 14451 1351 14454 1371
rect 14454 1351 14485 1371
rect 14526 1351 14558 1371
rect 14558 1351 14560 1371
rect 14601 1351 14628 1371
rect 14628 1351 14635 1371
rect 15733 1348 15754 1367
rect 15754 1348 15767 1367
rect 15819 1348 15824 1367
rect 15824 1348 15853 1367
rect 15905 1348 15928 1367
rect 15928 1348 15939 1367
rect 15991 1348 15998 1367
rect 15998 1348 16025 1367
rect 15733 1333 15767 1348
rect 15819 1333 15853 1348
rect 15905 1333 15939 1348
rect 15991 1333 16025 1348
rect 478 1274 480 1308
rect 480 1274 512 1308
rect 550 1274 582 1308
rect 582 1274 584 1308
rect 3380 1274 3382 1308
rect 3382 1274 3414 1308
rect 3452 1274 3484 1308
rect 3484 1274 3486 1308
rect 12882 1274 12884 1308
rect 12884 1274 12916 1308
rect 12954 1274 12986 1308
rect 12986 1274 12988 1308
rect 360 1259 394 1268
rect 360 1234 394 1259
rect 15733 1280 15754 1294
rect 15754 1280 15767 1294
rect 15819 1280 15824 1294
rect 15824 1280 15853 1294
rect 15905 1280 15928 1294
rect 15928 1280 15939 1294
rect 15991 1280 15998 1294
rect 15998 1280 16025 1294
rect 15733 1260 15767 1280
rect 15819 1260 15853 1280
rect 15905 1260 15939 1280
rect 15991 1260 16025 1280
rect 360 1189 394 1196
rect 360 1162 394 1189
rect 15733 1212 15754 1221
rect 15754 1212 15767 1221
rect 15819 1212 15824 1221
rect 15824 1212 15853 1221
rect 15905 1212 15928 1221
rect 15928 1212 15939 1221
rect 15991 1212 15998 1221
rect 15998 1212 16025 1221
rect 15733 1187 15767 1212
rect 15819 1187 15853 1212
rect 15905 1187 15939 1212
rect 15991 1187 16025 1212
rect 360 1119 394 1124
rect 360 1090 394 1119
rect 478 1120 480 1154
rect 480 1120 512 1154
rect 550 1120 582 1154
rect 582 1120 584 1154
rect 3380 1120 3382 1154
rect 3382 1120 3414 1154
rect 3452 1120 3484 1154
rect 3484 1120 3486 1154
rect 12882 1120 12884 1154
rect 12884 1120 12916 1154
rect 12954 1120 12986 1154
rect 12986 1120 12988 1154
rect 15733 1144 15754 1148
rect 15754 1144 15767 1148
rect 15819 1144 15824 1148
rect 15824 1144 15853 1148
rect 15905 1144 15928 1148
rect 15928 1144 15939 1148
rect 15991 1144 15998 1148
rect 15998 1144 16025 1148
rect 15733 1114 15767 1144
rect 15819 1114 15853 1144
rect 15905 1114 15939 1144
rect 15991 1114 16025 1144
rect 360 1050 394 1052
rect 360 1018 394 1050
rect 13168 1057 13194 1077
rect 13194 1057 13202 1077
rect 13244 1057 13264 1077
rect 13264 1057 13278 1077
rect 13320 1057 13334 1077
rect 13334 1057 13354 1077
rect 13396 1057 13404 1077
rect 13404 1057 13430 1077
rect 13472 1057 13474 1077
rect 13474 1057 13506 1077
rect 13548 1057 13578 1077
rect 13578 1057 13582 1077
rect 13624 1057 13648 1077
rect 13648 1057 13658 1077
rect 13700 1057 13718 1077
rect 13718 1057 13734 1077
rect 13776 1057 13788 1077
rect 13788 1057 13810 1077
rect 13851 1057 13858 1077
rect 13858 1057 13885 1077
rect 13926 1057 13928 1077
rect 13928 1057 13960 1077
rect 14001 1057 14034 1077
rect 14034 1057 14035 1077
rect 14076 1057 14104 1077
rect 14104 1057 14110 1077
rect 14151 1057 14174 1077
rect 14174 1057 14185 1077
rect 14226 1057 14244 1077
rect 14244 1057 14260 1077
rect 14301 1057 14314 1077
rect 14314 1057 14335 1077
rect 14376 1057 14384 1077
rect 14384 1057 14410 1077
rect 14451 1057 14454 1077
rect 14454 1057 14485 1077
rect 14526 1057 14558 1077
rect 14558 1057 14560 1077
rect 14601 1057 14628 1077
rect 14628 1057 14635 1077
rect 13168 1043 13202 1057
rect 13244 1043 13278 1057
rect 13320 1043 13354 1057
rect 13396 1043 13430 1057
rect 13472 1043 13506 1057
rect 13548 1043 13582 1057
rect 13624 1043 13658 1057
rect 13700 1043 13734 1057
rect 13776 1043 13810 1057
rect 13851 1043 13885 1057
rect 13926 1043 13960 1057
rect 14001 1043 14035 1057
rect 14076 1043 14110 1057
rect 14151 1043 14185 1057
rect 14226 1043 14260 1057
rect 14301 1043 14335 1057
rect 14376 1043 14410 1057
rect 14451 1043 14485 1057
rect 14526 1043 14560 1057
rect 14601 1043 14635 1057
rect 15733 1042 15767 1075
rect 15819 1042 15853 1075
rect 15905 1042 15939 1075
rect 15991 1042 16025 1075
rect 360 947 394 980
rect 360 946 394 947
rect 478 966 480 1000
rect 480 966 512 1000
rect 550 966 582 1000
rect 582 966 584 1000
rect 3380 966 3382 1000
rect 3382 966 3414 1000
rect 3452 966 3484 1000
rect 3484 966 3486 1000
rect 12882 966 12884 1000
rect 12884 966 12916 1000
rect 12954 966 12986 1000
rect 12986 966 12988 1000
rect 15733 1041 15754 1042
rect 15754 1041 15767 1042
rect 15819 1041 15824 1042
rect 15824 1041 15853 1042
rect 15905 1041 15928 1042
rect 15928 1041 15939 1042
rect 15991 1041 15998 1042
rect 15998 1041 16025 1042
rect 15733 974 15767 1002
rect 15819 974 15853 1002
rect 15905 974 15939 1002
rect 15991 974 16025 1002
rect 360 878 394 908
rect 360 874 394 878
rect 15733 968 15754 974
rect 15754 968 15767 974
rect 15819 968 15824 974
rect 15824 968 15853 974
rect 15905 968 15928 974
rect 15928 968 15939 974
rect 15991 968 15998 974
rect 15998 968 16025 974
rect 15733 906 15767 929
rect 15819 906 15853 929
rect 15905 906 15939 929
rect 15991 906 16025 929
rect 15733 895 15754 906
rect 15754 895 15767 906
rect 15819 895 15824 906
rect 15824 895 15853 906
rect 15905 895 15928 906
rect 15928 895 15939 906
rect 15991 895 15998 906
rect 15998 895 16025 906
rect 360 809 394 836
rect 360 802 394 809
rect 478 812 480 846
rect 480 812 512 846
rect 550 812 582 846
rect 582 812 584 846
rect 3380 812 3382 846
rect 3382 812 3414 846
rect 3452 812 3484 846
rect 3484 812 3486 846
rect 12882 812 12884 846
rect 12884 812 12916 846
rect 12954 812 12986 846
rect 12986 812 12988 846
rect 15733 838 15767 856
rect 15819 838 15853 856
rect 15905 838 15939 856
rect 15991 838 16025 856
rect 360 740 394 764
rect 360 730 394 740
rect 15733 822 15754 838
rect 15754 822 15767 838
rect 15819 822 15824 838
rect 15824 822 15853 838
rect 15905 822 15928 838
rect 15928 822 15939 838
rect 15991 822 15998 838
rect 15998 822 16025 838
rect 15733 770 15767 783
rect 15819 770 15853 783
rect 15905 770 15939 783
rect 15991 770 16025 783
rect 13168 741 13202 769
rect 13244 741 13278 769
rect 13320 741 13354 769
rect 13396 741 13430 769
rect 13472 741 13506 769
rect 13548 741 13582 769
rect 13624 741 13658 769
rect 13700 741 13734 769
rect 13776 741 13810 769
rect 13851 741 13885 769
rect 13926 741 13960 769
rect 14001 741 14035 769
rect 14076 741 14110 769
rect 14151 741 14185 769
rect 14226 741 14260 769
rect 14301 741 14335 769
rect 14376 741 14410 769
rect 14451 741 14485 769
rect 14526 741 14560 769
rect 14601 741 14635 769
rect 13168 735 13194 741
rect 13194 735 13202 741
rect 13244 735 13264 741
rect 13264 735 13278 741
rect 13320 735 13334 741
rect 13334 735 13354 741
rect 13396 735 13404 741
rect 13404 735 13430 741
rect 13472 735 13474 741
rect 13474 735 13506 741
rect 360 671 394 692
rect 360 658 394 671
rect 13548 735 13578 741
rect 13578 735 13582 741
rect 13624 735 13648 741
rect 13648 735 13658 741
rect 13700 735 13718 741
rect 13718 735 13734 741
rect 13776 735 13788 741
rect 13788 735 13810 741
rect 13851 735 13858 741
rect 13858 735 13885 741
rect 13926 735 13928 741
rect 13928 735 13960 741
rect 14001 735 14034 741
rect 14034 735 14035 741
rect 14076 735 14104 741
rect 14104 735 14110 741
rect 14151 735 14174 741
rect 14174 735 14185 741
rect 14226 735 14244 741
rect 14244 735 14260 741
rect 14301 735 14314 741
rect 14314 735 14335 741
rect 14376 735 14384 741
rect 14384 735 14410 741
rect 14451 735 14454 741
rect 14454 735 14485 741
rect 14526 735 14558 741
rect 14558 735 14560 741
rect 14601 735 14628 741
rect 14628 735 14635 741
rect 15733 749 15754 770
rect 15754 749 15767 770
rect 15819 749 15824 770
rect 15824 749 15853 770
rect 15905 749 15928 770
rect 15928 749 15939 770
rect 15991 749 15998 770
rect 15998 749 16025 770
rect 15733 702 15767 710
rect 15819 702 15853 710
rect 15905 702 15939 710
rect 15991 702 16025 710
rect 478 658 480 692
rect 480 658 512 692
rect 550 658 582 692
rect 582 658 584 692
rect 3380 658 3382 692
rect 3382 658 3414 692
rect 3452 658 3484 692
rect 3484 658 3486 692
rect 12882 658 12884 692
rect 12884 658 12916 692
rect 12954 658 12986 692
rect 12986 658 12988 692
rect 360 602 394 620
rect 360 586 394 602
rect 360 533 394 548
rect 360 514 394 533
rect 15733 676 15754 702
rect 15754 676 15767 702
rect 15819 676 15824 702
rect 15824 676 15853 702
rect 15905 676 15928 702
rect 15928 676 15939 702
rect 15991 676 15998 702
rect 15998 676 16025 702
rect 15733 634 15767 637
rect 15819 634 15853 637
rect 15905 634 15939 637
rect 15991 634 16025 637
rect 15733 603 15754 634
rect 15754 603 15767 634
rect 15819 603 15824 634
rect 15824 603 15853 634
rect 15905 603 15928 634
rect 15928 603 15939 634
rect 15991 603 15998 634
rect 15998 603 16025 634
rect 478 504 480 538
rect 480 504 512 538
rect 550 504 582 538
rect 582 504 584 538
rect 3380 504 3382 538
rect 3382 504 3414 538
rect 3452 504 3484 538
rect 3484 504 3486 538
rect 12882 504 12884 538
rect 12884 504 12916 538
rect 12954 504 12986 538
rect 12986 504 12988 538
rect 15733 532 15754 564
rect 15754 532 15767 564
rect 15819 532 15824 564
rect 15824 532 15853 564
rect 15905 532 15928 564
rect 15928 532 15939 564
rect 15991 532 15998 564
rect 15998 532 16025 564
rect 360 464 394 476
rect 360 442 394 464
rect 15733 530 15767 532
rect 15819 530 15853 532
rect 15905 530 15939 532
rect 15991 530 16025 532
rect 360 395 394 404
rect 360 370 394 395
rect 15733 464 15754 491
rect 15754 464 15767 491
rect 15819 464 15824 491
rect 15824 464 15853 491
rect 15905 464 15928 491
rect 15928 464 15939 491
rect 15991 464 15998 491
rect 15998 464 16025 491
rect 13168 427 13194 461
rect 13194 427 13202 461
rect 13241 427 13264 461
rect 13264 427 13275 461
rect 13314 427 13334 461
rect 13334 427 13348 461
rect 13387 427 13404 461
rect 13404 427 13421 461
rect 13460 427 13474 461
rect 13474 427 13494 461
rect 13533 427 13544 461
rect 13544 427 13567 461
rect 13606 427 13614 461
rect 13614 427 13640 461
rect 13679 427 13684 461
rect 13684 427 13713 461
rect 13752 427 13754 461
rect 13754 427 13786 461
rect 13825 427 13858 461
rect 13858 427 13859 461
rect 13898 427 13928 461
rect 13928 427 13932 461
rect 13971 427 13998 461
rect 13998 427 14005 461
rect 14044 427 14068 461
rect 14068 427 14078 461
rect 14117 427 14138 461
rect 14138 427 14151 461
rect 14190 427 14208 461
rect 14208 427 14224 461
rect 14263 427 14278 461
rect 14278 427 14297 461
rect 14336 427 14348 461
rect 14348 427 14370 461
rect 14409 427 14418 461
rect 14418 427 14443 461
rect 14482 427 14488 461
rect 14488 427 14516 461
rect 14555 427 14558 461
rect 14558 427 14589 461
rect 14628 427 14662 461
rect 14701 427 14735 461
rect 14774 430 14808 461
rect 14847 430 14881 461
rect 14920 430 14954 461
rect 14993 430 15027 461
rect 15065 430 15099 461
rect 15137 430 15171 461
rect 15209 430 15243 461
rect 15281 430 15315 461
rect 15353 430 15387 461
rect 15425 430 15459 461
rect 15497 430 15531 461
rect 15569 430 15603 461
rect 15641 430 15675 461
rect 15733 457 15767 464
rect 15819 457 15853 464
rect 15905 457 15939 464
rect 15991 457 16025 464
rect 14774 427 14808 430
rect 14847 427 14878 430
rect 14878 427 14881 430
rect 14920 427 14948 430
rect 14948 427 14954 430
rect 14993 427 15018 430
rect 15018 427 15027 430
rect 15065 427 15088 430
rect 15088 427 15099 430
rect 15137 427 15158 430
rect 15158 427 15171 430
rect 15209 427 15228 430
rect 15228 427 15243 430
rect 15281 427 15298 430
rect 15298 427 15315 430
rect 15353 427 15368 430
rect 15368 427 15387 430
rect 15425 427 15438 430
rect 15438 427 15459 430
rect 15497 427 15508 430
rect 15508 427 15531 430
rect 15569 427 15578 430
rect 15578 427 15603 430
rect 15641 427 15648 430
rect 15648 427 15675 430
rect 15733 396 15754 418
rect 15754 396 15767 418
rect 15819 396 15824 418
rect 15824 396 15853 418
rect 15905 396 15928 418
rect 15928 396 15939 418
rect 15991 396 15998 418
rect 15998 396 16025 418
rect 360 326 394 332
rect 360 298 394 326
rect 478 350 480 384
rect 480 350 512 384
rect 550 350 582 384
rect 582 350 584 384
rect 3380 350 3382 384
rect 3382 350 3414 384
rect 3452 350 3484 384
rect 3484 350 3486 384
rect 12882 350 12884 384
rect 12884 350 12916 384
rect 12954 350 12986 384
rect 12986 350 12988 384
rect 15733 384 15767 396
rect 15819 384 15853 396
rect 15905 384 15939 396
rect 15991 384 16025 396
rect 360 257 394 260
rect 360 226 394 257
rect 15733 328 15754 345
rect 15754 328 15767 345
rect 15819 328 15824 345
rect 15824 328 15853 345
rect 15905 328 15928 345
rect 15928 328 15939 345
rect 15991 328 15998 345
rect 15998 328 16025 345
rect 15733 311 15767 328
rect 15819 311 15853 328
rect 15905 311 15939 328
rect 15991 311 16025 328
rect 15733 260 15754 272
rect 15754 260 15767 272
rect 15819 260 15824 272
rect 15824 260 15853 272
rect 15905 260 15928 272
rect 15928 260 15939 272
rect 15991 260 15998 272
rect 15998 260 16025 272
rect 360 154 394 188
rect 478 196 480 230
rect 480 196 512 230
rect 550 196 582 230
rect 582 196 584 230
rect 3380 196 3382 230
rect 3382 196 3414 230
rect 3452 196 3484 230
rect 3484 196 3486 230
rect 12882 196 12884 230
rect 12884 196 12916 230
rect 12954 196 12986 230
rect 12986 196 12988 230
rect 15733 238 15767 260
rect 15819 238 15853 260
rect 15905 238 15939 260
rect 15991 238 16025 260
rect 15733 192 15754 199
rect 15754 192 15767 199
rect 15819 192 15824 199
rect 15824 192 15853 199
rect 15905 192 15928 199
rect 15928 192 15939 199
rect 15991 192 15998 199
rect 15998 192 16025 199
rect 15733 165 15767 192
rect 15819 165 15853 192
rect 15905 165 15939 192
rect 15991 165 16025 192
rect 15733 124 15754 126
rect 15754 124 15767 126
rect 15819 124 15824 126
rect 15824 124 15853 126
rect 15905 124 15928 126
rect 15928 124 15939 126
rect 15991 124 15998 126
rect 15998 124 16025 126
rect 15733 92 15767 124
rect 15819 92 15853 124
rect 15905 92 15939 124
rect 15991 92 16025 124
rect 389 50 394 84
rect 394 50 423 84
rect 461 50 463 84
rect 463 50 495 84
rect 533 50 567 84
rect 605 50 636 84
rect 636 50 639 84
rect 677 50 705 84
rect 705 50 711 84
rect 915 50 946 84
rect 946 50 949 84
rect 987 50 1015 84
rect 1015 50 1021 84
rect 1059 50 1084 84
rect 1084 50 1093 84
rect 1131 50 1153 84
rect 1153 50 1165 84
rect 1203 50 1222 84
rect 1222 50 1237 84
rect 1275 50 1291 84
rect 1291 50 1309 84
rect 1347 50 1360 84
rect 1360 50 1381 84
rect 1419 50 1429 84
rect 1429 50 1453 84
rect 1491 50 1498 84
rect 1498 50 1525 84
rect 1563 50 1567 84
rect 1567 50 1597 84
rect 1635 50 1636 84
rect 1636 50 1669 84
rect 1707 50 1740 84
rect 1740 50 1741 84
rect 1779 50 1809 84
rect 1809 50 1813 84
rect 1851 50 1878 84
rect 1878 50 1885 84
rect 1923 50 1947 84
rect 1947 50 1957 84
rect 1995 50 2016 84
rect 2016 50 2029 84
rect 2067 50 2085 84
rect 2085 50 2101 84
rect 2139 50 2154 84
rect 2154 50 2173 84
rect 2211 50 2223 84
rect 2223 50 2245 84
rect 2283 50 2292 84
rect 2292 50 2317 84
rect 2355 50 2361 84
rect 2361 50 2389 84
rect 2427 50 2430 84
rect 2430 50 2461 84
rect 2499 50 2533 84
rect 2571 50 2602 84
rect 2602 50 2605 84
rect 2643 50 2671 84
rect 2671 50 2677 84
rect 2715 50 2740 84
rect 2740 50 2749 84
rect 2787 50 2809 84
rect 2809 50 2821 84
rect 2859 50 2878 84
rect 2878 50 2893 84
rect 2931 50 2947 84
rect 2947 50 2965 84
rect 3003 50 3016 84
rect 3016 50 3037 84
rect 3075 50 3085 84
rect 3085 50 3109 84
rect 3147 50 3154 84
rect 3154 50 3181 84
rect 3219 50 3223 84
rect 3223 50 3253 84
rect 3291 50 3292 84
rect 3292 50 3325 84
rect 3363 50 3396 84
rect 3396 50 3397 84
rect 3435 50 3465 84
rect 3465 50 3469 84
rect 3507 50 3534 84
rect 3534 50 3541 84
rect 3579 50 3603 84
rect 3603 50 3613 84
rect 3651 50 3672 84
rect 3672 50 3685 84
rect 3723 50 3741 84
rect 3741 50 3757 84
rect 3795 50 3810 84
rect 3810 50 3829 84
rect 3867 50 3879 84
rect 3879 50 3901 84
rect 3939 50 3948 84
rect 3948 50 3973 84
rect 4011 50 4017 84
rect 4017 50 4045 84
rect 4083 50 4086 84
rect 4086 50 4117 84
rect 4155 50 4189 84
rect 4227 50 4258 84
rect 4258 50 4261 84
rect 4299 50 4327 84
rect 4327 50 4333 84
rect 4371 50 4396 84
rect 4396 50 4405 84
rect 4443 50 4465 84
rect 4465 50 4477 84
rect 4515 50 4534 84
rect 4534 50 4549 84
rect 4587 50 4603 84
rect 4603 50 4621 84
rect 4659 50 4672 84
rect 4672 50 4693 84
rect 4731 50 4741 84
rect 4741 50 4765 84
rect 4803 50 4810 84
rect 4810 50 4837 84
rect 4875 50 4879 84
rect 4879 50 4909 84
rect 4947 50 4948 84
rect 4948 50 4981 84
rect 5019 50 5050 84
rect 5050 50 5053 84
rect 5091 50 5118 84
rect 5118 50 5125 84
rect 5163 50 5186 84
rect 5186 50 5197 84
rect 5235 50 5254 84
rect 5254 50 5269 84
rect 5307 50 5322 84
rect 5322 50 5341 84
rect 5379 50 5390 84
rect 5390 50 5413 84
rect 5451 50 5458 84
rect 5458 50 5485 84
rect 5523 50 5526 84
rect 5526 50 5557 84
rect 5595 50 5628 84
rect 5628 50 5629 84
rect 5667 50 5696 84
rect 5696 50 5701 84
rect 5739 50 5764 84
rect 5764 50 5773 84
rect 5811 50 5832 84
rect 5832 50 5845 84
rect 5883 50 5900 84
rect 5900 50 5917 84
rect 5955 50 5968 84
rect 5968 50 5989 84
rect 6027 50 6036 84
rect 6036 50 6061 84
rect 6099 50 6104 84
rect 6104 50 6133 84
rect 6171 50 6172 84
rect 6172 50 6205 84
rect 6243 50 6274 84
rect 6274 50 6277 84
rect 6315 50 6342 84
rect 6342 50 6349 84
rect 6387 50 6410 84
rect 6410 50 6421 84
rect 6459 50 6478 84
rect 6478 50 6493 84
rect 6531 50 6546 84
rect 6546 50 6565 84
rect 6603 50 6614 84
rect 6614 50 6637 84
rect 6675 50 6682 84
rect 6682 50 6709 84
rect 6747 50 6750 84
rect 6750 50 6781 84
rect 6819 50 6852 84
rect 6852 50 6853 84
rect 6891 50 6920 84
rect 6920 50 6925 84
rect 6963 50 6988 84
rect 6988 50 6997 84
rect 7035 50 7056 84
rect 7056 50 7069 84
rect 7107 50 7124 84
rect 7124 50 7141 84
rect 7179 50 7192 84
rect 7192 50 7213 84
rect 7251 50 7260 84
rect 7260 50 7285 84
rect 7323 50 7328 84
rect 7328 50 7357 84
rect 7395 50 7396 84
rect 7396 50 7429 84
rect 7467 50 7498 84
rect 7498 50 7501 84
rect 7539 50 7566 84
rect 7566 50 7573 84
rect 7611 50 7634 84
rect 7634 50 7645 84
rect 7683 50 7702 84
rect 7702 50 7717 84
rect 7755 50 7770 84
rect 7770 50 7789 84
rect 7827 50 7838 84
rect 7838 50 7861 84
rect 7899 50 7906 84
rect 7906 50 7933 84
rect 7971 50 7974 84
rect 7974 50 8005 84
rect 8043 50 8076 84
rect 8076 50 8077 84
rect 8115 50 8144 84
rect 8144 50 8149 84
rect 8187 50 8212 84
rect 8212 50 8221 84
rect 8259 50 8280 84
rect 8280 50 8293 84
rect 8331 50 8348 84
rect 8348 50 8365 84
rect 8403 50 8416 84
rect 8416 50 8437 84
rect 8475 50 8484 84
rect 8484 50 8509 84
rect 8547 50 8552 84
rect 8552 50 8581 84
rect 8619 50 8620 84
rect 8620 50 8653 84
rect 8691 50 8722 84
rect 8722 50 8725 84
rect 8763 50 8790 84
rect 8790 50 8797 84
rect 8835 50 8858 84
rect 8858 50 8869 84
rect 8907 50 8926 84
rect 8926 50 8941 84
rect 8979 50 8994 84
rect 8994 50 9013 84
rect 9051 50 9062 84
rect 9062 50 9085 84
rect 9123 50 9130 84
rect 9130 50 9157 84
rect 9195 50 9198 84
rect 9198 50 9229 84
rect 9267 50 9300 84
rect 9300 50 9301 84
rect 9339 50 9368 84
rect 9368 50 9373 84
rect 9411 50 9436 84
rect 9436 50 9445 84
rect 9483 50 9504 84
rect 9504 50 9517 84
rect 9555 50 9572 84
rect 9572 50 9589 84
rect 9627 50 9640 84
rect 9640 50 9661 84
rect 9699 50 9708 84
rect 9708 50 9733 84
rect 9771 50 9776 84
rect 9776 50 9805 84
rect 9843 50 9844 84
rect 9844 50 9877 84
rect 9915 50 9946 84
rect 9946 50 9949 84
rect 9987 50 10014 84
rect 10014 50 10021 84
rect 10059 50 10082 84
rect 10082 50 10093 84
rect 10131 50 10150 84
rect 10150 50 10165 84
rect 10203 50 10218 84
rect 10218 50 10237 84
rect 10275 50 10286 84
rect 10286 50 10309 84
rect 10347 50 10354 84
rect 10354 50 10381 84
rect 10419 50 10422 84
rect 10422 50 10453 84
rect 10491 50 10524 84
rect 10524 50 10525 84
rect 10563 50 10592 84
rect 10592 50 10597 84
rect 10635 50 10660 84
rect 10660 50 10669 84
rect 10707 50 10728 84
rect 10728 50 10741 84
rect 10779 50 10796 84
rect 10796 50 10813 84
rect 10851 50 10864 84
rect 10864 50 10885 84
rect 10923 50 10932 84
rect 10932 50 10957 84
rect 10995 50 11000 84
rect 11000 50 11029 84
rect 11067 50 11068 84
rect 11068 50 11101 84
rect 11139 50 11170 84
rect 11170 50 11173 84
rect 11211 50 11238 84
rect 11238 50 11245 84
rect 11283 50 11306 84
rect 11306 50 11317 84
rect 11355 50 11374 84
rect 11374 50 11389 84
rect 11427 50 11442 84
rect 11442 50 11461 84
rect 11499 50 11510 84
rect 11510 50 11533 84
rect 11571 50 11578 84
rect 11578 50 11605 84
rect 11643 50 11646 84
rect 11646 50 11677 84
rect 11715 50 11748 84
rect 11748 50 11749 84
rect 11787 50 11816 84
rect 11816 50 11821 84
rect 11859 50 11884 84
rect 11884 50 11893 84
rect 11931 50 11952 84
rect 11952 50 11965 84
rect 12003 50 12020 84
rect 12020 50 12037 84
rect 12075 50 12088 84
rect 12088 50 12109 84
rect 12147 50 12156 84
rect 12156 50 12181 84
rect 12219 50 12224 84
rect 12224 50 12253 84
rect 12291 50 12292 84
rect 12292 50 12325 84
rect 12363 50 12394 84
rect 12394 50 12397 84
rect 12435 50 12462 84
rect 12462 50 12469 84
rect 12507 50 12530 84
rect 12530 50 12541 84
rect 12579 50 12598 84
rect 12598 50 12613 84
rect 12651 50 12666 84
rect 12666 50 12685 84
rect 12723 50 12734 84
rect 12734 50 12757 84
rect 12795 50 12802 84
rect 12802 50 12829 84
rect 12867 50 12870 84
rect 12870 50 12901 84
rect 12939 50 12972 84
rect 12972 50 12973 84
rect 13011 50 13040 84
rect 13040 50 13045 84
rect 13083 50 13108 84
rect 13108 50 13117 84
rect 13155 50 13176 84
rect 13176 50 13189 84
rect 13227 50 13244 84
rect 13244 50 13261 84
rect 13299 50 13312 84
rect 13312 50 13333 84
rect 13371 50 13380 84
rect 13380 50 13405 84
rect 13443 50 13448 84
rect 13448 50 13477 84
rect 13515 50 13516 84
rect 13516 50 13549 84
rect 13587 50 13618 84
rect 13618 50 13621 84
rect 13659 50 13686 84
rect 13686 50 13693 84
rect 13731 50 13754 84
rect 13754 50 13765 84
rect 13803 50 13822 84
rect 13822 50 13837 84
rect 13875 50 13890 84
rect 13890 50 13909 84
rect 13947 50 13958 84
rect 13958 50 13981 84
rect 14019 50 14026 84
rect 14026 50 14053 84
rect 14091 50 14094 84
rect 14094 50 14125 84
rect 14163 50 14196 84
rect 14196 50 14197 84
rect 14235 50 14264 84
rect 14264 50 14269 84
rect 14307 50 14332 84
rect 14332 50 14341 84
rect 15733 50 15760 53
rect 15760 50 15767 53
rect 15819 50 15828 53
rect 15828 50 15853 53
rect 15905 50 15930 53
rect 15930 50 15939 53
rect 15991 50 15998 53
rect 15998 50 16025 53
rect 15733 19 15767 50
rect 15819 19 15853 50
rect 15905 19 15939 50
rect 15991 19 16025 50
<< metal1 >>
rect 348 7975 354 8027
rect 406 7975 418 8027
rect 470 8018 482 8027
rect 534 8018 546 8027
rect 598 8018 610 8027
rect 662 8018 674 8027
rect 726 8018 857 8027
rect 909 8018 921 8027
rect 973 8018 985 8027
rect 1037 8018 1049 8027
rect 1101 8018 1113 8027
rect 1165 8018 1177 8027
rect 1229 8018 1241 8027
rect 479 7984 482 8018
rect 726 7984 745 8018
rect 779 7984 857 8018
rect 910 7984 921 8018
rect 982 7984 985 8018
rect 1229 7984 1236 8018
rect 470 7975 482 7984
rect 534 7975 546 7984
rect 598 7975 610 7984
rect 662 7975 674 7984
rect 726 7975 857 7984
rect 909 7975 921 7984
rect 973 7975 985 7984
rect 1037 7975 1049 7984
rect 1101 7975 1113 7984
rect 1165 7975 1177 7984
rect 1229 7975 1241 7984
rect 1293 7975 1305 8027
rect 1357 7975 1369 8027
rect 1421 7975 1433 8027
rect 1485 8018 1497 8027
rect 1549 8018 1561 8027
rect 1613 8018 1625 8027
rect 1677 8018 1689 8027
rect 1741 8018 1753 8027
rect 1805 8018 1817 8027
rect 1486 7984 1497 8018
rect 1558 7984 1561 8018
rect 1805 7984 1812 8018
rect 1485 7975 1497 7984
rect 1549 7975 1561 7984
rect 1613 7975 1625 7984
rect 1677 7975 1689 7984
rect 1741 7975 1753 7984
rect 1805 7975 1817 7984
rect 1869 7975 1881 8027
rect 1933 7975 1945 8027
rect 1997 7975 2009 8027
rect 2061 8018 2073 8027
rect 2125 8018 2137 8027
rect 2189 8018 2201 8027
rect 2253 8018 2265 8027
rect 2317 8018 2329 8027
rect 2381 8018 2393 8027
rect 2062 7984 2073 8018
rect 2134 7984 2137 8018
rect 2381 7984 2388 8018
rect 2061 7975 2073 7984
rect 2125 7975 2137 7984
rect 2189 7975 2201 7984
rect 2253 7975 2265 7984
rect 2317 7975 2329 7984
rect 2381 7975 2393 7984
rect 2445 7975 2457 8027
rect 2509 7975 2521 8027
rect 2573 7975 2585 8027
rect 2637 8018 2649 8027
rect 2701 8018 2713 8027
rect 2765 8018 2777 8027
rect 2829 8018 2841 8027
rect 2893 8018 2905 8027
rect 2957 8018 2969 8027
rect 2638 7984 2649 8018
rect 2710 7984 2713 8018
rect 2957 7984 2964 8018
rect 2637 7975 2649 7984
rect 2701 7975 2713 7984
rect 2765 7975 2777 7984
rect 2829 7975 2841 7984
rect 2893 7975 2905 7984
rect 2957 7975 2969 7984
rect 3021 7975 3033 8027
rect 3085 7975 3097 8027
rect 3149 7975 3161 8027
rect 3213 8018 3225 8027
rect 3277 8018 3289 8027
rect 3341 8018 3353 8027
rect 3405 8018 3417 8027
rect 3469 8018 3481 8027
rect 3533 8018 3545 8027
rect 3214 7984 3225 8018
rect 3286 7984 3289 8018
rect 3533 7984 3540 8018
rect 3213 7975 3225 7984
rect 3277 7975 3289 7984
rect 3341 7975 3353 7984
rect 3405 7975 3417 7984
rect 3469 7975 3481 7984
rect 3533 7975 3545 7984
rect 3597 7975 3609 8027
rect 3661 7975 3673 8027
rect 3725 7975 3737 8027
rect 3789 8018 3801 8027
rect 3853 8018 3865 8027
rect 3917 8018 3929 8027
rect 3981 8018 3993 8027
rect 4045 8018 4057 8027
rect 4109 8018 4121 8027
rect 3790 7984 3801 8018
rect 3862 7984 3865 8018
rect 4109 7984 4116 8018
rect 3789 7975 3801 7984
rect 3853 7975 3865 7984
rect 3917 7975 3929 7984
rect 3981 7975 3993 7984
rect 4045 7975 4057 7984
rect 4109 7975 4121 7984
rect 4173 7975 4185 8027
rect 4237 7975 4249 8027
rect 4301 7975 4313 8027
rect 4365 8018 4377 8027
rect 4429 8018 4441 8027
rect 4493 8018 4505 8027
rect 4557 8018 4722 8027
rect 4774 8018 4786 8027
rect 4838 8018 4850 8027
rect 4902 8018 4914 8027
rect 4366 7984 4377 8018
rect 4438 7984 4441 8018
rect 4557 7984 4583 8018
rect 4617 7984 4657 8018
rect 4691 7984 4722 8018
rect 4902 7984 4910 8018
rect 4365 7975 4377 7984
rect 4429 7975 4441 7984
rect 4493 7975 4505 7984
rect 4557 7975 4722 7984
rect 4774 7975 4786 7984
rect 4838 7975 4850 7984
rect 4902 7975 4914 7984
rect 4966 7975 4978 8027
rect 5030 7975 5042 8027
rect 5094 7975 5106 8027
rect 5158 8018 5170 8027
rect 5222 8018 5234 8027
rect 5286 8018 5298 8027
rect 5350 8018 5362 8027
rect 5414 8018 5426 8027
rect 5478 8018 5490 8027
rect 5160 7984 5170 8018
rect 5232 7984 5234 8018
rect 5478 7984 5486 8018
rect 5158 7975 5170 7984
rect 5222 7975 5234 7984
rect 5286 7975 5298 7984
rect 5350 7975 5362 7984
rect 5414 7975 5426 7984
rect 5478 7975 5490 7984
rect 5542 7975 5554 8027
rect 5606 7975 5618 8027
rect 5670 7975 5682 8027
rect 5734 8018 5746 8027
rect 5798 8018 5810 8027
rect 5862 8018 5874 8027
rect 5926 8018 5938 8027
rect 5990 8018 6002 8027
rect 6054 8018 6066 8027
rect 5736 7984 5746 8018
rect 5808 7984 5810 8018
rect 6054 7984 6062 8018
rect 5734 7975 5746 7984
rect 5798 7975 5810 7984
rect 5862 7975 5874 7984
rect 5926 7975 5938 7984
rect 5990 7975 6002 7984
rect 6054 7975 6066 7984
rect 6118 7975 6130 8027
rect 6182 7975 6194 8027
rect 6246 7975 6258 8027
rect 6310 8018 6322 8027
rect 6374 8018 6386 8027
rect 6438 8018 6450 8027
rect 6502 8018 6514 8027
rect 6566 8018 6578 8027
rect 6630 8018 6810 8027
rect 6862 8018 6874 8027
rect 6926 8018 6938 8027
rect 6990 8018 7002 8027
rect 6312 7984 6322 8018
rect 6384 7984 6386 8018
rect 6630 7984 6667 8018
rect 6701 7984 6741 8018
rect 6775 7984 6810 8018
rect 6990 7984 6994 8018
rect 6310 7975 6322 7984
rect 6374 7975 6386 7984
rect 6438 7975 6450 7984
rect 6502 7975 6514 7984
rect 6566 7975 6578 7984
rect 6630 7975 6810 7984
rect 6862 7975 6874 7984
rect 6926 7975 6938 7984
rect 6990 7975 7002 7984
rect 7054 7975 7066 8027
rect 7118 7975 7130 8027
rect 7182 7975 7194 8027
rect 7246 7975 7258 8027
rect 7310 8018 7322 8027
rect 7374 8018 7386 8027
rect 7438 8018 7450 8027
rect 7502 8018 7514 8027
rect 7566 8018 7578 8027
rect 7316 7984 7322 8018
rect 7566 7984 7570 8018
rect 7310 7975 7322 7984
rect 7374 7975 7386 7984
rect 7438 7975 7450 7984
rect 7502 7975 7514 7984
rect 7566 7975 7578 7984
rect 7630 7975 7642 8027
rect 7694 7975 7706 8027
rect 7758 7975 7770 8027
rect 7822 7975 7834 8027
rect 7886 8018 7898 8027
rect 7950 8018 7962 8027
rect 8014 8018 8026 8027
rect 8078 8018 8090 8027
rect 8142 8018 8154 8027
rect 7892 7984 7898 8018
rect 8142 7984 8146 8018
rect 7886 7975 7898 7984
rect 7950 7975 7962 7984
rect 8014 7975 8026 7984
rect 8078 7975 8090 7984
rect 8142 7975 8154 7984
rect 8206 7975 8218 8027
rect 8270 7975 8282 8027
rect 8334 7975 8346 8027
rect 8398 7975 8410 8027
rect 8462 8018 8474 8027
rect 8526 8018 8538 8027
rect 8590 8018 8602 8027
rect 8654 8018 8666 8027
rect 8718 8018 8730 8027
rect 8468 7984 8474 8018
rect 8718 7984 8722 8018
rect 8462 7975 8474 7984
rect 8526 7975 8538 7984
rect 8590 7975 8602 7984
rect 8654 7975 8666 7984
rect 8718 7975 8730 7984
rect 8782 7975 8794 8027
rect 8846 7975 8858 8027
rect 8910 7975 8922 8027
rect 8974 7975 8986 8027
rect 9038 8018 9050 8027
rect 9102 8018 9114 8027
rect 9166 8018 9178 8027
rect 9230 8018 9242 8027
rect 9294 8018 9306 8027
rect 9044 7984 9050 8018
rect 9294 7984 9298 8018
rect 9038 7975 9050 7984
rect 9102 7975 9114 7984
rect 9166 7975 9178 7984
rect 9230 7975 9242 7984
rect 9294 7975 9306 7984
rect 9358 7975 9370 8027
rect 9422 7975 9434 8027
rect 9486 7975 9498 8027
rect 9550 7975 9562 8027
rect 9614 8018 9626 8027
rect 9678 8018 9690 8027
rect 9742 8018 9754 8027
rect 9806 8018 9818 8027
rect 9870 8018 9882 8027
rect 9620 7984 9626 8018
rect 9870 7984 9874 8018
rect 9614 7975 9626 7984
rect 9678 7975 9690 7984
rect 9742 7975 9754 7984
rect 9806 7975 9818 7984
rect 9870 7975 9882 7984
rect 9934 7975 9946 8027
rect 9998 7975 10010 8027
rect 10062 7975 10074 8027
rect 10126 7975 10138 8027
rect 10190 8018 10202 8027
rect 10254 8018 10266 8027
rect 10318 8018 10330 8027
rect 10382 8018 10394 8027
rect 10446 8018 10458 8027
rect 10196 7984 10202 8018
rect 10446 7984 10450 8018
rect 10190 7975 10202 7984
rect 10254 7975 10266 7984
rect 10318 7975 10330 7984
rect 10382 7975 10394 7984
rect 10446 7975 10458 7984
rect 10510 7975 10522 8027
rect 10574 7975 10586 8027
rect 10638 7975 10650 8027
rect 10702 7975 10714 8027
rect 10766 8018 10778 8027
rect 10830 8018 10842 8027
rect 10894 8018 10906 8027
rect 10958 8018 10970 8027
rect 11022 8018 11034 8027
rect 10772 7984 10778 8018
rect 11022 7984 11026 8018
rect 10766 7975 10778 7984
rect 10830 7975 10842 7984
rect 10894 7975 10906 7984
rect 10958 7975 10970 7984
rect 11022 7975 11034 7984
rect 11086 7975 11098 8027
rect 11150 7975 11162 8027
rect 11214 7975 11226 8027
rect 11278 7975 11290 8027
rect 11342 8018 11354 8027
rect 11406 8018 11418 8027
rect 11470 8018 11482 8027
rect 11534 8018 11546 8027
rect 11598 8018 11610 8027
rect 11348 7984 11354 8018
rect 11598 7984 11602 8018
rect 11342 7975 11354 7984
rect 11406 7975 11418 7984
rect 11470 7975 11482 7984
rect 11534 7975 11546 7984
rect 11598 7975 11610 7984
rect 11662 7975 11674 8027
rect 11726 7975 11738 8027
rect 11790 7975 11802 8027
rect 11854 7975 11866 8027
rect 11918 8018 11930 8027
rect 11982 8018 11994 8027
rect 12046 8018 12058 8027
rect 12110 8018 12122 8027
rect 12174 8018 12186 8027
rect 11924 7984 11930 8018
rect 12174 7984 12178 8018
rect 11918 7975 11930 7984
rect 11982 7975 11994 7984
rect 12046 7975 12058 7984
rect 12110 7975 12122 7984
rect 12174 7975 12186 7984
rect 12238 7975 12250 8027
rect 12302 7975 12314 8027
rect 12366 7975 12378 8027
rect 12430 7975 12442 8027
rect 12494 8018 12506 8027
rect 12558 8018 12570 8027
rect 12622 8018 12634 8027
rect 12686 8018 12698 8027
rect 12750 8018 12762 8027
rect 12500 7984 12506 8018
rect 12750 7984 12754 8018
rect 12494 7975 12506 7984
rect 12558 7975 12570 7984
rect 12622 7975 12634 7984
rect 12686 7975 12698 7984
rect 12750 7975 12762 7984
rect 12814 7975 12826 8027
rect 12878 7975 12890 8027
rect 12942 7975 12954 8027
rect 13006 7975 13018 8027
rect 13070 8018 13082 8027
rect 13134 8018 13146 8027
rect 13198 8018 13210 8027
rect 13262 8018 13274 8027
rect 13326 8018 13338 8027
rect 13076 7984 13082 8018
rect 13326 7984 13330 8018
rect 13070 7975 13082 7984
rect 13134 7975 13146 7984
rect 13198 7975 13210 7984
rect 13262 7975 13274 7984
rect 13326 7975 13338 7984
rect 13390 7975 13402 8027
rect 13454 7975 13466 8027
rect 13518 7975 13530 8027
rect 13582 7975 13594 8027
rect 13646 7975 13652 8027
rect 348 7966 360 7975
rect 394 7966 421 7975
rect 348 7938 421 7966
tri 421 7938 458 7975 nw
rect 348 7928 406 7938
rect 348 7894 360 7928
rect 394 7894 406 7928
tri 406 7923 421 7938 nw
tri 13678 7923 13684 7929 se
rect 13684 7923 13736 8108
rect 15725 8010 16033 8042
rect 15725 7976 15733 8010
rect 15767 7976 15819 8010
rect 15853 7976 15905 8010
rect 15939 7976 15991 8010
rect 16025 7976 16033 8010
rect 15725 7938 16033 7976
tri 13736 7923 13742 7929 sw
tri 13659 7904 13678 7923 se
rect 13678 7904 13742 7923
tri 13742 7904 13761 7923 sw
rect 15725 7904 15733 7938
rect 15767 7904 15819 7938
rect 15853 7904 15905 7938
rect 15939 7904 15991 7938
rect 16025 7904 16033 7938
rect 348 7856 406 7894
tri 13637 7882 13659 7904 se
rect 13659 7882 13761 7904
tri 13761 7882 13783 7904 sw
rect 348 7822 360 7856
rect 394 7822 406 7856
rect 348 7784 406 7822
rect 348 7750 360 7784
rect 394 7750 406 7784
rect 348 7712 406 7750
rect 348 7678 360 7712
rect 394 7678 406 7712
rect 348 7640 406 7678
rect 466 7830 473 7882
rect 525 7830 537 7882
rect 589 7830 596 7882
rect 3203 7830 3209 7882
rect 3261 7830 3273 7882
rect 3325 7830 3333 7882
rect 3334 7831 3335 7881
rect 3363 7831 3364 7881
rect 3365 7873 3498 7882
rect 3365 7839 3380 7873
rect 3414 7839 3452 7873
rect 3486 7839 3498 7873
rect 3365 7830 3498 7839
rect 12870 7873 15255 7882
rect 12870 7839 12882 7873
rect 12916 7839 12954 7873
rect 12988 7866 15255 7873
tri 15255 7866 15271 7882 sw
rect 15725 7866 16033 7904
rect 12988 7864 15271 7866
tri 15271 7864 15273 7866 sw
rect 12988 7839 15273 7864
rect 12870 7832 15273 7839
tri 15273 7832 15305 7864 sw
rect 15725 7832 15733 7866
rect 15767 7832 15819 7866
rect 15853 7832 15905 7866
rect 15939 7832 15991 7866
rect 16025 7832 16033 7866
rect 12870 7830 15305 7832
tri 15305 7830 15307 7832 sw
rect 466 7728 596 7830
tri 15233 7794 15269 7830 ne
rect 15269 7794 15307 7830
tri 15307 7794 15343 7830 sw
rect 15725 7794 16033 7832
tri 15269 7790 15273 7794 ne
rect 15273 7790 15343 7794
tri 15343 7790 15347 7794 sw
tri 15273 7760 15303 7790 ne
rect 15303 7760 15347 7790
tri 15347 7760 15377 7790 sw
rect 15725 7760 15733 7794
rect 15767 7760 15819 7794
rect 15853 7760 15905 7794
rect 15939 7760 15991 7794
rect 16025 7760 16033 7794
tri 15303 7728 15335 7760 ne
rect 15335 7728 15377 7760
tri 15377 7728 15409 7760 sw
rect 466 7676 473 7728
rect 525 7676 537 7728
rect 589 7676 596 7728
rect 3207 7676 3213 7728
rect 3265 7676 3277 7728
rect 3329 7726 3337 7728
rect 3338 7727 3364 7728
rect 3365 7726 3498 7728
rect 3329 7719 3498 7726
rect 3329 7685 3380 7719
rect 3414 7685 3452 7719
rect 3486 7685 3498 7719
rect 3329 7678 3498 7685
rect 3329 7676 3337 7678
rect 3338 7676 3364 7677
rect 3365 7676 3498 7678
rect 10278 7676 10285 7728
rect 10337 7676 10349 7728
rect 10401 7676 10408 7728
rect 12870 7724 15189 7728
tri 15189 7724 15193 7728 sw
tri 15335 7724 15339 7728 ne
rect 15339 7724 15409 7728
tri 15409 7724 15413 7728 sw
rect 12870 7722 15193 7724
tri 15193 7722 15195 7724 sw
tri 15339 7722 15341 7724 ne
rect 15341 7722 15413 7724
tri 15413 7722 15415 7724 sw
rect 15725 7722 16033 7760
rect 12870 7719 15195 7722
rect 12870 7685 12882 7719
rect 12916 7685 12954 7719
rect 12988 7688 15195 7719
tri 15195 7688 15229 7722 sw
tri 15341 7716 15347 7722 ne
rect 15347 7716 15415 7722
tri 15415 7716 15421 7722 sw
tri 15347 7688 15375 7716 ne
rect 15375 7688 15421 7716
tri 15421 7688 15449 7716 sw
rect 15725 7688 15733 7722
rect 15767 7688 15819 7722
rect 15853 7688 15905 7722
rect 15939 7688 15991 7722
rect 16025 7688 16033 7722
rect 12988 7685 15229 7688
rect 12870 7676 15229 7685
tri 15229 7676 15241 7688 sw
tri 15375 7676 15387 7688 ne
rect 15387 7676 15449 7688
tri 15449 7676 15461 7688 sw
rect 348 7606 360 7640
rect 394 7606 406 7640
rect 348 7568 406 7606
rect 348 7534 360 7568
rect 394 7534 406 7568
rect 348 7496 406 7534
rect 348 7462 360 7496
rect 394 7462 406 7496
rect 348 7424 406 7462
rect 348 7390 360 7424
rect 394 7390 406 7424
rect 348 7352 406 7390
rect 466 7522 473 7574
rect 525 7522 537 7574
rect 589 7522 596 7574
rect 3203 7522 3209 7574
rect 3261 7522 3273 7574
rect 3325 7522 3333 7574
rect 3334 7523 3335 7573
rect 3363 7523 3364 7573
rect 3365 7565 3498 7574
rect 3365 7531 3380 7565
rect 3414 7531 3452 7565
rect 3486 7531 3498 7565
rect 3365 7522 3498 7531
rect 466 7420 596 7522
rect 466 7368 473 7420
rect 525 7368 537 7420
rect 589 7368 596 7420
rect 3207 7368 3213 7420
rect 3265 7368 3277 7420
rect 3329 7418 3337 7420
rect 3338 7419 3364 7420
rect 3365 7418 3498 7420
rect 3329 7411 3498 7418
rect 3329 7377 3380 7411
rect 3414 7377 3452 7411
rect 3486 7377 3498 7411
rect 3329 7370 3498 7377
rect 3329 7368 3337 7370
rect 3338 7368 3364 7369
rect 3365 7368 3498 7370
rect 9422 7368 9429 7420
rect 9481 7368 9493 7420
rect 9545 7368 9552 7420
rect 348 7318 360 7352
rect 394 7318 406 7352
rect 348 7280 406 7318
rect 348 7246 360 7280
rect 394 7246 406 7280
rect 348 7208 406 7246
rect 348 7174 360 7208
rect 394 7174 406 7208
rect 348 7136 406 7174
rect 348 7102 360 7136
rect 394 7102 406 7136
rect 348 7064 406 7102
rect 348 7030 360 7064
rect 394 7030 406 7064
rect 466 7214 473 7266
rect 525 7214 537 7266
rect 589 7214 596 7266
rect 3203 7214 3209 7266
rect 3261 7214 3273 7266
rect 3325 7214 3333 7266
rect 3334 7215 3335 7265
rect 3363 7215 3364 7265
rect 3365 7257 3498 7266
rect 3365 7223 3380 7257
rect 3414 7223 3452 7257
rect 3486 7223 3498 7257
rect 3365 7214 3498 7223
rect 466 7112 596 7214
rect 466 7060 473 7112
rect 525 7060 537 7112
rect 589 7060 596 7112
rect 3207 7060 3213 7112
rect 3265 7060 3277 7112
rect 3329 7110 3337 7112
rect 3338 7111 3364 7112
rect 3365 7110 3498 7112
rect 3329 7103 3498 7110
rect 3329 7069 3380 7103
rect 3414 7069 3452 7103
rect 3486 7069 3498 7103
rect 3329 7062 3498 7069
rect 3329 7060 3337 7062
rect 3338 7060 3364 7061
rect 3365 7060 3498 7062
rect 8566 7060 8573 7112
rect 8625 7060 8637 7112
rect 8689 7060 8696 7112
rect 348 6992 406 7030
rect 348 6958 360 6992
rect 394 6958 406 6992
rect 348 6920 406 6958
rect 348 6886 360 6920
rect 394 6886 406 6920
rect 348 6848 406 6886
rect 348 6814 360 6848
rect 394 6814 406 6848
rect 348 6776 406 6814
rect 348 6742 360 6776
rect 394 6742 406 6776
rect 466 6906 473 6958
rect 525 6906 537 6958
rect 589 6906 596 6958
rect 3203 6906 3209 6958
rect 3261 6906 3273 6958
rect 3325 6906 3333 6958
rect 3334 6907 3335 6957
rect 3363 6907 3364 6957
rect 3365 6949 3498 6958
rect 3365 6915 3380 6949
rect 3414 6915 3452 6949
rect 3486 6915 3498 6949
rect 3365 6906 3498 6915
rect 466 6804 596 6906
rect 466 6752 473 6804
rect 525 6752 537 6804
rect 589 6752 596 6804
rect 3207 6752 3213 6804
rect 3265 6752 3277 6804
rect 3329 6802 3337 6804
rect 3338 6803 3364 6804
rect 3365 6802 3498 6804
rect 3329 6795 3498 6802
rect 3329 6761 3380 6795
rect 3414 6761 3452 6795
rect 3486 6761 3498 6795
rect 3329 6754 3498 6761
rect 3329 6752 3337 6754
rect 3338 6752 3364 6753
rect 3365 6752 3498 6754
rect 7710 6752 7717 6804
rect 7769 6752 7781 6804
rect 7833 6752 7840 6804
rect 348 6704 406 6742
rect 348 6670 360 6704
rect 394 6670 406 6704
rect 348 6632 406 6670
rect 348 6598 360 6632
rect 394 6598 406 6632
rect 348 6560 406 6598
rect 348 6526 360 6560
rect 394 6526 406 6560
rect 348 6488 406 6526
rect 348 6454 360 6488
rect 394 6454 406 6488
rect 348 6416 406 6454
rect 466 6598 473 6650
rect 525 6598 537 6650
rect 589 6598 596 6650
rect 3203 6598 3209 6650
rect 3261 6598 3273 6650
rect 3325 6598 3333 6650
rect 3334 6599 3335 6649
rect 3363 6599 3364 6649
rect 3365 6641 3498 6650
rect 3365 6607 3380 6641
rect 3414 6607 3452 6641
rect 3486 6607 3498 6641
rect 3365 6598 3498 6607
rect 466 6496 596 6598
rect 466 6444 473 6496
rect 525 6444 537 6496
rect 589 6444 596 6496
rect 3207 6444 3213 6496
rect 3265 6444 3277 6496
rect 3329 6494 3337 6496
rect 3338 6495 3364 6496
rect 3365 6494 3498 6496
rect 3329 6487 3498 6494
rect 3329 6453 3380 6487
rect 3414 6453 3452 6487
rect 3486 6453 3498 6487
rect 3329 6446 3498 6453
rect 3329 6444 3337 6446
rect 3338 6444 3364 6445
rect 3365 6444 3498 6446
rect 6854 6444 6861 6496
rect 6913 6444 6925 6496
rect 6977 6444 6984 6496
rect 348 6382 360 6416
rect 394 6382 406 6416
rect 348 6344 406 6382
rect 348 6310 360 6344
rect 394 6310 406 6344
rect 348 6272 406 6310
rect 348 6238 360 6272
rect 394 6238 406 6272
rect 348 6200 406 6238
rect 348 6166 360 6200
rect 394 6166 406 6200
rect 348 6128 406 6166
rect 466 6290 473 6342
rect 525 6290 537 6342
rect 589 6290 596 6342
rect 3203 6290 3209 6342
rect 3261 6290 3273 6342
rect 3325 6290 3333 6342
rect 3334 6291 3335 6341
rect 3363 6291 3364 6341
rect 3365 6333 3498 6342
rect 3365 6299 3380 6333
rect 3414 6299 3452 6333
rect 3486 6299 3498 6333
rect 3365 6290 3498 6299
rect 466 6188 596 6290
rect 466 6136 473 6188
rect 525 6136 537 6188
rect 589 6136 596 6188
rect 3207 6136 3213 6188
rect 3265 6136 3277 6188
rect 3329 6186 3337 6188
rect 3338 6187 3364 6188
rect 3365 6186 3498 6188
rect 3329 6179 3498 6186
rect 3329 6145 3380 6179
rect 3414 6145 3452 6179
rect 3486 6145 3498 6179
rect 3329 6138 3498 6145
rect 3329 6136 3337 6138
rect 3338 6136 3364 6137
rect 3365 6136 3498 6138
rect 5998 6136 6005 6188
rect 6057 6136 6069 6188
rect 6121 6136 6128 6188
rect 348 6094 360 6128
rect 394 6094 406 6128
rect 348 6066 406 6094
tri 406 6066 434 6094 sw
rect 348 6042 434 6066
tri 434 6042 458 6066 sw
rect 348 5990 354 6042
rect 406 6033 418 6042
rect 470 6033 482 6042
rect 534 6033 546 6042
rect 598 6033 610 6042
rect 598 5999 605 6033
rect 406 5990 418 5999
rect 470 5990 482 5999
rect 534 5990 546 5999
rect 598 5990 610 5999
rect 662 5990 674 6042
rect 726 6032 869 6042
rect 921 6033 933 6042
rect 985 6033 997 6042
rect 1049 6033 1061 6042
rect 726 5998 765 6032
rect 799 5998 837 6032
rect 985 5999 986 6033
rect 1049 5999 1058 6033
rect 726 5990 869 5998
rect 921 5990 933 5999
rect 985 5990 997 5999
rect 1049 5990 1061 5999
rect 1113 5990 1125 6042
rect 1177 5990 1189 6042
rect 1241 5990 1253 6042
rect 1305 6033 1317 6042
rect 1369 6033 1381 6042
rect 1433 6033 1445 6042
rect 1497 6033 1509 6042
rect 1561 6033 1573 6042
rect 1625 6033 1637 6042
rect 1308 5999 1317 6033
rect 1380 5999 1381 6033
rect 1561 5999 1562 6033
rect 1625 5999 1634 6033
rect 1305 5990 1317 5999
rect 1369 5990 1381 5999
rect 1433 5990 1445 5999
rect 1497 5990 1509 5999
rect 1561 5990 1573 5999
rect 1625 5990 1637 5999
rect 1689 5990 1701 6042
rect 1753 5990 1765 6042
rect 1817 5990 1829 6042
rect 1881 6033 1893 6042
rect 1945 6033 1957 6042
rect 2009 6033 2021 6042
rect 2073 6033 2085 6042
rect 2137 6033 2149 6042
rect 2201 6033 2213 6042
rect 1884 5999 1893 6033
rect 1956 5999 1957 6033
rect 2137 5999 2138 6033
rect 2201 5999 2210 6033
rect 1881 5990 1893 5999
rect 1945 5990 1957 5999
rect 2009 5990 2021 5999
rect 2073 5990 2085 5999
rect 2137 5990 2149 5999
rect 2201 5990 2213 5999
rect 2265 5990 2277 6042
rect 2329 5990 2341 6042
rect 2393 5990 2405 6042
rect 2457 6033 2469 6042
rect 2521 6033 2533 6042
rect 2585 6033 2597 6042
rect 2649 6033 2661 6042
rect 2713 6033 2725 6042
rect 2777 6033 2789 6042
rect 2460 5999 2469 6033
rect 2532 5999 2533 6033
rect 2713 5999 2714 6033
rect 2777 5999 2786 6033
rect 2457 5990 2469 5999
rect 2521 5990 2533 5999
rect 2585 5990 2597 5999
rect 2649 5990 2661 5999
rect 2713 5990 2725 5999
rect 2777 5990 2789 5999
rect 2841 5990 2853 6042
rect 2905 5990 2917 6042
rect 2969 5990 2981 6042
rect 3033 6033 3045 6042
rect 3097 6033 3109 6042
rect 3161 6033 3173 6042
rect 3225 6033 3237 6042
rect 3289 6033 3301 6042
rect 3353 6033 3365 6042
rect 3036 5999 3045 6033
rect 3108 5999 3109 6033
rect 3289 5999 3290 6033
rect 3353 5999 3362 6033
rect 3033 5990 3045 5999
rect 3097 5990 3109 5999
rect 3161 5990 3173 5999
rect 3225 5990 3237 5999
rect 3289 5990 3301 5999
rect 3353 5990 3365 5999
rect 3417 5990 3429 6042
rect 3481 5990 3493 6042
rect 3545 5990 3557 6042
rect 3609 6033 3621 6042
rect 3673 6033 3685 6042
rect 3737 6033 3749 6042
rect 3801 6033 3813 6042
rect 3865 6033 3877 6042
rect 3929 6033 3941 6042
rect 3612 5999 3621 6033
rect 3684 5999 3685 6033
rect 3865 5999 3866 6033
rect 3929 5999 3938 6033
rect 3609 5990 3621 5999
rect 3673 5990 3685 5999
rect 3737 5990 3749 5999
rect 3801 5990 3813 5999
rect 3865 5990 3877 5999
rect 3929 5990 3941 5999
rect 3993 5990 4005 6042
rect 4057 5990 4069 6042
rect 4121 5990 4133 6042
rect 4185 6033 4197 6042
rect 4249 6033 4261 6042
rect 4313 6033 4325 6042
rect 4377 6033 4389 6042
rect 4441 6033 4453 6042
rect 4505 6033 4517 6042
rect 4188 5999 4197 6033
rect 4260 5999 4261 6033
rect 4441 5999 4442 6033
rect 4505 5999 4514 6033
rect 4569 6032 4757 6042
rect 4185 5990 4197 5999
rect 4249 5990 4261 5999
rect 4313 5990 4325 5999
rect 4377 5990 4389 5999
rect 4441 5990 4453 5999
rect 4505 5990 4517 5999
rect 4569 5998 4618 6032
rect 4652 5998 4690 6032
rect 4724 5998 4757 6032
rect 4569 5990 4757 5998
rect 4809 5990 4821 6042
rect 4873 6033 4885 6042
rect 4937 6033 4949 6042
rect 5001 6033 5013 6042
rect 5065 6033 5077 6042
rect 5129 6033 5141 6042
rect 4879 5999 4885 6033
rect 5129 5999 5133 6033
rect 4873 5990 4885 5999
rect 4937 5990 4949 5999
rect 5001 5990 5013 5999
rect 5065 5990 5077 5999
rect 5129 5990 5141 5999
rect 5193 5990 5205 6042
rect 5257 5990 5269 6042
rect 5321 5990 5333 6042
rect 5385 5990 5397 6042
rect 5449 6033 5461 6042
rect 5513 6033 5525 6042
rect 5577 6033 5589 6042
rect 5641 6033 5653 6042
rect 5705 6033 5717 6042
rect 5455 5999 5461 6033
rect 5705 5999 5709 6033
rect 5449 5990 5461 5999
rect 5513 5990 5525 5999
rect 5577 5990 5589 5999
rect 5641 5990 5653 5999
rect 5705 5990 5717 5999
rect 5769 5990 5781 6042
rect 5833 5990 5845 6042
rect 5897 5990 5903 6042
rect 348 5756 354 5808
rect 406 5756 418 5808
rect 470 5756 482 5808
rect 534 5799 546 5808
rect 598 5799 610 5808
rect 662 5799 674 5808
rect 726 5799 738 5808
rect 790 5799 802 5808
rect 540 5765 546 5799
rect 790 5765 794 5799
rect 534 5756 546 5765
rect 598 5756 610 5765
rect 662 5756 674 5765
rect 726 5756 738 5765
rect 790 5756 802 5765
rect 854 5756 866 5808
rect 918 5756 930 5808
rect 982 5756 994 5808
rect 1046 5756 1058 5808
rect 1110 5799 1122 5808
rect 1174 5799 1186 5808
rect 1238 5799 1250 5808
rect 1302 5799 1314 5808
rect 1366 5799 1378 5808
rect 1116 5765 1122 5799
rect 1366 5765 1370 5799
rect 1110 5756 1122 5765
rect 1174 5756 1186 5765
rect 1238 5756 1250 5765
rect 1302 5756 1314 5765
rect 1366 5756 1378 5765
rect 1430 5756 1442 5808
rect 1494 5756 1506 5808
rect 1558 5756 1570 5808
rect 1622 5756 1634 5808
rect 1686 5799 1698 5808
rect 1750 5799 1762 5808
rect 1814 5799 1826 5808
rect 1878 5799 1890 5808
rect 1942 5799 1954 5808
rect 1692 5765 1698 5799
rect 1942 5765 1946 5799
rect 1686 5756 1698 5765
rect 1750 5756 1762 5765
rect 1814 5756 1826 5765
rect 1878 5756 1890 5765
rect 1942 5756 1954 5765
rect 2006 5756 2018 5808
rect 2070 5756 2082 5808
rect 2134 5756 2146 5808
rect 2198 5756 2210 5808
rect 2262 5799 2274 5808
rect 2326 5799 2338 5808
rect 2390 5799 2402 5808
rect 2454 5799 2466 5808
rect 2518 5799 2530 5808
rect 2268 5765 2274 5799
rect 2518 5765 2522 5799
rect 2262 5756 2274 5765
rect 2326 5756 2338 5765
rect 2390 5756 2402 5765
rect 2454 5756 2466 5765
rect 2518 5756 2530 5765
rect 2582 5756 2594 5808
rect 2646 5756 2658 5808
rect 2710 5756 2722 5808
rect 2774 5756 2786 5808
rect 2838 5799 2850 5808
rect 2902 5799 2914 5808
rect 2966 5799 2978 5808
rect 3030 5799 3042 5808
rect 3094 5799 3106 5808
rect 2844 5765 2850 5799
rect 3094 5765 3098 5799
rect 2838 5756 2850 5765
rect 2902 5756 2914 5765
rect 2966 5756 2978 5765
rect 3030 5756 3042 5765
rect 3094 5756 3106 5765
rect 3158 5756 3170 5808
rect 3222 5756 3234 5808
rect 3286 5756 3298 5808
rect 3350 5756 3362 5808
rect 3414 5799 3427 5808
rect 3479 5799 3492 5808
rect 3544 5799 3557 5808
rect 3609 5799 3622 5808
rect 3674 5799 3687 5808
rect 3739 5799 3752 5808
rect 3420 5765 3427 5799
rect 3739 5765 3746 5799
rect 3414 5756 3427 5765
rect 3479 5756 3492 5765
rect 3544 5756 3557 5765
rect 3609 5756 3622 5765
rect 3674 5756 3687 5765
rect 3739 5756 3752 5765
rect 3804 5756 3817 5808
rect 3869 5756 3882 5808
rect 3934 5756 3947 5808
rect 3999 5756 4012 5808
rect 4064 5799 4077 5808
rect 4129 5799 4142 5808
rect 4194 5799 4207 5808
rect 4259 5799 4272 5808
rect 4324 5799 4337 5808
rect 4389 5799 4402 5808
rect 4454 5799 4467 5808
rect 4068 5765 4077 5799
rect 4140 5765 4142 5799
rect 4389 5765 4394 5799
rect 4454 5765 4466 5799
rect 4064 5756 4077 5765
rect 4129 5756 4142 5765
rect 4194 5756 4207 5765
rect 4259 5756 4272 5765
rect 4324 5756 4337 5765
rect 4389 5756 4402 5765
rect 4454 5756 4467 5765
rect 4519 5756 4532 5808
rect 4584 5756 4597 5808
rect 4649 5756 4662 5808
rect 4714 5799 4727 5808
rect 4779 5799 4792 5808
rect 4844 5799 4857 5808
rect 4909 5799 4922 5808
rect 4974 5799 4987 5808
rect 5039 5799 5052 5808
rect 5104 5799 5117 5808
rect 4716 5765 4727 5799
rect 4788 5765 4792 5799
rect 5039 5765 5042 5799
rect 5104 5765 5114 5799
rect 4714 5756 4727 5765
rect 4779 5756 4792 5765
rect 4844 5756 4857 5765
rect 4909 5756 4922 5765
rect 4974 5756 4987 5765
rect 5039 5756 5052 5765
rect 5104 5756 5117 5765
rect 5169 5756 5182 5808
rect 5234 5756 5247 5808
rect 5299 5756 5312 5808
rect 5364 5756 5377 5808
rect 5429 5799 5442 5808
rect 5494 5799 5507 5808
rect 5559 5799 5572 5808
rect 5624 5799 5637 5808
rect 5689 5799 5702 5808
rect 5754 5799 5767 5808
rect 5436 5765 5442 5799
rect 5689 5765 5690 5799
rect 5754 5765 5763 5799
rect 5429 5756 5442 5765
rect 5494 5756 5507 5765
rect 5559 5756 5572 5765
rect 5624 5756 5637 5765
rect 5689 5756 5702 5765
rect 5754 5756 5767 5765
rect 5819 5756 5832 5808
rect 5884 5756 5897 5808
rect 5949 5756 5955 5808
rect 348 5731 360 5756
rect 394 5744 446 5756
tri 446 5744 458 5756 nw
rect 394 5734 436 5744
tri 436 5734 446 5744 nw
rect 394 5731 412 5734
rect 348 5710 412 5731
tri 412 5710 436 5734 nw
rect 348 5693 406 5710
tri 406 5704 412 5710 nw
rect 348 5659 360 5693
rect 394 5659 406 5693
rect 348 5621 406 5659
rect 348 5587 360 5621
rect 394 5587 406 5621
rect 348 5549 406 5587
rect 348 5515 360 5549
rect 394 5515 406 5549
rect 348 5477 406 5515
rect 348 5443 360 5477
rect 394 5443 406 5477
rect 348 5405 406 5443
rect 348 5402 360 5405
rect 394 5402 406 5405
rect 348 5350 351 5402
rect 403 5350 406 5402
rect 348 5338 406 5350
rect 348 5286 351 5338
rect 403 5286 406 5338
rect 348 5274 406 5286
rect 348 5222 351 5274
rect 403 5222 406 5274
rect 348 5210 406 5222
rect 348 5158 351 5210
rect 403 5158 406 5210
rect 348 5155 360 5158
rect 394 5155 406 5158
rect 348 5146 406 5155
rect 348 5094 351 5146
rect 403 5094 406 5146
rect 348 5083 360 5094
rect 394 5083 406 5094
rect 348 5082 406 5083
rect 348 5030 351 5082
rect 403 5030 406 5082
rect 348 5018 360 5030
rect 394 5018 406 5030
rect 348 4966 351 5018
rect 403 4966 406 5018
rect 348 4954 360 4966
rect 394 4954 406 4966
rect 348 4902 351 4954
rect 403 4902 406 4954
rect 348 4901 406 4902
rect 348 4890 360 4901
rect 394 4890 406 4901
rect 348 4838 351 4890
rect 403 4838 406 4890
rect 348 4829 406 4838
rect 348 4826 360 4829
rect 394 4826 406 4829
rect 348 4774 351 4826
rect 403 4774 406 4826
rect 348 4762 406 4774
rect 348 4710 351 4762
rect 403 4710 406 4762
rect 348 4698 406 4710
rect 348 4646 351 4698
rect 403 4646 406 4698
rect 348 4634 406 4646
rect 348 4582 351 4634
rect 403 4582 406 4634
rect 348 4579 360 4582
rect 394 4579 406 4582
rect 348 4570 406 4579
rect 348 4518 351 4570
rect 403 4518 406 4570
rect 348 4507 360 4518
rect 394 4507 406 4518
rect 468 5411 526 5417
rect 468 5402 480 5411
rect 514 5402 526 5411
rect 468 5350 471 5402
rect 523 5350 526 5402
rect 468 5339 526 5350
rect 468 5338 480 5339
rect 514 5338 526 5339
rect 468 5286 471 5338
rect 523 5286 526 5338
rect 468 5274 526 5286
rect 468 5222 471 5274
rect 523 5222 526 5274
rect 468 5210 526 5222
rect 468 5158 471 5210
rect 523 5158 526 5210
rect 468 5146 526 5158
rect 468 5094 471 5146
rect 523 5094 526 5146
rect 468 5089 480 5094
rect 514 5089 526 5094
rect 468 5082 526 5089
rect 468 5030 471 5082
rect 523 5030 526 5082
rect 468 5018 480 5030
rect 514 5018 526 5030
rect 468 4966 471 5018
rect 523 4966 526 5018
rect 468 4954 480 4966
rect 514 4954 526 4966
rect 468 4902 471 4954
rect 523 4902 526 4954
rect 468 4890 480 4902
rect 514 4890 526 4902
rect 468 4838 471 4890
rect 523 4838 526 4890
rect 468 4835 526 4838
rect 468 4826 480 4835
rect 514 4826 526 4835
rect 468 4774 471 4826
rect 523 4774 526 4826
rect 468 4763 526 4774
rect 468 4762 480 4763
rect 514 4762 526 4763
rect 468 4710 471 4762
rect 523 4710 526 4762
rect 468 4698 526 4710
rect 468 4646 471 4698
rect 523 4646 526 4698
rect 468 4634 526 4646
rect 468 4582 471 4634
rect 523 4582 526 4634
rect 468 4570 526 4582
rect 468 4518 471 4570
rect 523 4518 526 4570
rect 468 4513 480 4518
rect 514 4513 526 4518
rect 468 4507 526 4513
rect 1324 5411 1382 5417
rect 1324 5402 1336 5411
rect 1370 5402 1382 5411
rect 1324 5350 1327 5402
rect 1379 5350 1382 5402
rect 1324 5339 1382 5350
rect 1324 5338 1336 5339
rect 1370 5338 1382 5339
rect 1324 5286 1327 5338
rect 1379 5286 1382 5338
rect 1324 5274 1382 5286
rect 1324 5222 1327 5274
rect 1379 5222 1382 5274
rect 1324 5210 1382 5222
rect 1324 5158 1327 5210
rect 1379 5158 1382 5210
rect 1324 5146 1382 5158
rect 1324 5094 1327 5146
rect 1379 5094 1382 5146
rect 1324 5089 1336 5094
rect 1370 5089 1382 5094
rect 1324 5082 1382 5089
rect 1324 5030 1327 5082
rect 1379 5030 1382 5082
rect 1324 5018 1336 5030
rect 1370 5018 1382 5030
rect 1324 4966 1327 5018
rect 1379 4966 1382 5018
rect 1324 4954 1336 4966
rect 1370 4954 1382 4966
rect 1324 4902 1327 4954
rect 1379 4902 1382 4954
rect 1324 4890 1336 4902
rect 1370 4890 1382 4902
rect 1324 4838 1327 4890
rect 1379 4838 1382 4890
rect 1324 4835 1382 4838
rect 1324 4826 1336 4835
rect 1370 4826 1382 4835
rect 1324 4774 1327 4826
rect 1379 4774 1382 4826
rect 1324 4763 1382 4774
rect 1324 4762 1336 4763
rect 1370 4762 1382 4763
rect 1324 4710 1327 4762
rect 1379 4710 1382 4762
rect 1324 4698 1382 4710
rect 1324 4646 1327 4698
rect 1379 4646 1382 4698
rect 1324 4634 1382 4646
rect 1324 4582 1327 4634
rect 1379 4582 1382 4634
rect 1324 4570 1382 4582
rect 1324 4518 1327 4570
rect 1379 4518 1382 4570
rect 1324 4513 1336 4518
rect 1370 4513 1382 4518
rect 1324 4507 1382 4513
rect 2180 5411 2238 5417
rect 2180 5402 2192 5411
rect 2226 5402 2238 5411
rect 2180 5350 2183 5402
rect 2235 5350 2238 5402
rect 2180 5339 2238 5350
rect 2180 5338 2192 5339
rect 2226 5338 2238 5339
rect 2180 5286 2183 5338
rect 2235 5286 2238 5338
rect 2180 5274 2238 5286
rect 2180 5222 2183 5274
rect 2235 5222 2238 5274
rect 2180 5210 2238 5222
rect 2180 5158 2183 5210
rect 2235 5158 2238 5210
rect 2180 5146 2238 5158
rect 2180 5094 2183 5146
rect 2235 5094 2238 5146
rect 2180 5089 2192 5094
rect 2226 5089 2238 5094
rect 2180 5082 2238 5089
rect 2180 5030 2183 5082
rect 2235 5030 2238 5082
rect 2180 5018 2192 5030
rect 2226 5018 2238 5030
rect 2180 4966 2183 5018
rect 2235 4966 2238 5018
rect 2180 4954 2192 4966
rect 2226 4954 2238 4966
rect 2180 4902 2183 4954
rect 2235 4902 2238 4954
rect 2180 4890 2192 4902
rect 2226 4890 2238 4902
rect 2180 4838 2183 4890
rect 2235 4838 2238 4890
rect 2180 4835 2238 4838
rect 2180 4826 2192 4835
rect 2226 4826 2238 4835
rect 2180 4774 2183 4826
rect 2235 4774 2238 4826
rect 2180 4763 2238 4774
rect 2180 4762 2192 4763
rect 2226 4762 2238 4763
rect 2180 4710 2183 4762
rect 2235 4710 2238 4762
rect 2180 4698 2238 4710
rect 2180 4646 2183 4698
rect 2235 4646 2238 4698
rect 2180 4634 2238 4646
rect 2180 4582 2183 4634
rect 2235 4582 2238 4634
rect 2180 4570 2238 4582
rect 2180 4518 2183 4570
rect 2235 4518 2238 4570
rect 2180 4513 2192 4518
rect 2226 4513 2238 4518
rect 2180 4507 2238 4513
rect 3036 5411 3094 5417
rect 3036 5402 3048 5411
rect 3082 5402 3094 5411
rect 3036 5350 3039 5402
rect 3091 5350 3094 5402
rect 3036 5339 3094 5350
rect 3036 5338 3048 5339
rect 3082 5338 3094 5339
rect 3036 5286 3039 5338
rect 3091 5286 3094 5338
rect 3036 5274 3094 5286
rect 3036 5222 3039 5274
rect 3091 5222 3094 5274
rect 3036 5210 3094 5222
rect 3036 5158 3039 5210
rect 3091 5158 3094 5210
rect 3036 5146 3094 5158
rect 3036 5094 3039 5146
rect 3091 5094 3094 5146
rect 3036 5089 3048 5094
rect 3082 5089 3094 5094
rect 3036 5082 3094 5089
rect 3036 5030 3039 5082
rect 3091 5030 3094 5082
rect 3036 5018 3048 5030
rect 3082 5018 3094 5030
rect 3036 4966 3039 5018
rect 3091 4966 3094 5018
rect 3036 4954 3048 4966
rect 3082 4954 3094 4966
rect 3036 4902 3039 4954
rect 3091 4902 3094 4954
rect 3036 4890 3048 4902
rect 3082 4890 3094 4902
rect 3036 4838 3039 4890
rect 3091 4838 3094 4890
rect 3036 4835 3094 4838
rect 3036 4826 3048 4835
rect 3082 4826 3094 4835
rect 3036 4774 3039 4826
rect 3091 4774 3094 4826
rect 3036 4763 3094 4774
rect 3036 4762 3048 4763
rect 3082 4762 3094 4763
rect 3036 4710 3039 4762
rect 3091 4710 3094 4762
rect 3036 4698 3094 4710
rect 3036 4646 3039 4698
rect 3091 4646 3094 4698
rect 3036 4634 3094 4646
rect 3036 4582 3039 4634
rect 3091 4582 3094 4634
rect 3036 4570 3094 4582
rect 3036 4518 3039 4570
rect 3091 4518 3094 4570
rect 3036 4513 3048 4518
rect 3082 4513 3094 4518
rect 3036 4507 3094 4513
rect 3892 5411 3950 5417
rect 3892 5402 3904 5411
rect 3938 5402 3950 5411
rect 3892 5350 3895 5402
rect 3947 5350 3950 5402
rect 3892 5339 3950 5350
rect 3892 5338 3904 5339
rect 3938 5338 3950 5339
rect 3892 5286 3895 5338
rect 3947 5286 3950 5338
rect 3892 5274 3950 5286
rect 3892 5222 3895 5274
rect 3947 5222 3950 5274
rect 3892 5210 3950 5222
rect 3892 5158 3895 5210
rect 3947 5158 3950 5210
rect 3892 5146 3950 5158
rect 3892 5094 3895 5146
rect 3947 5094 3950 5146
rect 3892 5089 3904 5094
rect 3938 5089 3950 5094
rect 3892 5082 3950 5089
rect 3892 5030 3895 5082
rect 3947 5030 3950 5082
rect 3892 5018 3904 5030
rect 3938 5018 3950 5030
rect 3892 4966 3895 5018
rect 3947 4966 3950 5018
rect 3892 4954 3904 4966
rect 3938 4954 3950 4966
rect 3892 4902 3895 4954
rect 3947 4902 3950 4954
rect 3892 4890 3904 4902
rect 3938 4890 3950 4902
rect 3892 4838 3895 4890
rect 3947 4838 3950 4890
rect 3892 4835 3950 4838
rect 3892 4826 3904 4835
rect 3938 4826 3950 4835
rect 3892 4774 3895 4826
rect 3947 4774 3950 4826
rect 3892 4763 3950 4774
rect 3892 4762 3904 4763
rect 3938 4762 3950 4763
rect 3892 4710 3895 4762
rect 3947 4710 3950 4762
rect 3892 4698 3950 4710
rect 3892 4646 3895 4698
rect 3947 4646 3950 4698
rect 3892 4634 3950 4646
rect 3892 4582 3895 4634
rect 3947 4582 3950 4634
rect 3892 4570 3950 4582
rect 3892 4518 3895 4570
rect 3947 4518 3950 4570
rect 3892 4513 3904 4518
rect 3938 4513 3950 4518
rect 3892 4507 3950 4513
rect 4748 5411 4806 5417
rect 4748 5402 4760 5411
rect 4794 5402 4806 5411
rect 4748 5350 4751 5402
rect 4803 5350 4806 5402
rect 4748 5339 4806 5350
rect 4748 5338 4760 5339
rect 4794 5338 4806 5339
rect 4748 5286 4751 5338
rect 4803 5286 4806 5338
rect 4748 5274 4806 5286
rect 4748 5222 4751 5274
rect 4803 5222 4806 5274
rect 4748 5210 4806 5222
rect 4748 5158 4751 5210
rect 4803 5158 4806 5210
rect 4748 5146 4806 5158
rect 4748 5094 4751 5146
rect 4803 5094 4806 5146
rect 4748 5089 4760 5094
rect 4794 5089 4806 5094
rect 4748 5082 4806 5089
rect 4748 5030 4751 5082
rect 4803 5030 4806 5082
rect 4748 5018 4760 5030
rect 4794 5018 4806 5030
rect 4748 4966 4751 5018
rect 4803 4966 4806 5018
rect 4748 4954 4760 4966
rect 4794 4954 4806 4966
rect 4748 4902 4751 4954
rect 4803 4902 4806 4954
rect 4748 4890 4760 4902
rect 4794 4890 4806 4902
rect 4748 4838 4751 4890
rect 4803 4838 4806 4890
rect 4748 4835 4806 4838
rect 4748 4826 4760 4835
rect 4794 4826 4806 4835
rect 4748 4774 4751 4826
rect 4803 4774 4806 4826
rect 4748 4763 4806 4774
rect 4748 4762 4760 4763
rect 4794 4762 4806 4763
rect 4748 4710 4751 4762
rect 4803 4710 4806 4762
rect 4748 4698 4806 4710
rect 4748 4646 4751 4698
rect 4803 4646 4806 4698
rect 4748 4634 4806 4646
rect 4748 4582 4751 4634
rect 4803 4582 4806 4634
rect 4748 4570 4806 4582
rect 4748 4518 4751 4570
rect 4803 4518 4806 4570
rect 4748 4513 4760 4518
rect 4794 4513 4806 4518
rect 4748 4507 4806 4513
rect 5604 5411 5662 5417
rect 5604 5402 5616 5411
rect 5650 5402 5662 5411
rect 5604 5350 5607 5402
rect 5659 5350 5662 5402
rect 5604 5339 5662 5350
rect 5604 5338 5616 5339
rect 5650 5338 5662 5339
rect 5604 5286 5607 5338
rect 5659 5286 5662 5338
rect 5604 5274 5662 5286
rect 5604 5222 5607 5274
rect 5659 5222 5662 5274
rect 5604 5210 5662 5222
rect 5604 5158 5607 5210
rect 5659 5158 5662 5210
rect 5604 5146 5662 5158
rect 5604 5094 5607 5146
rect 5659 5094 5662 5146
rect 5604 5089 5616 5094
rect 5650 5089 5662 5094
rect 5604 5082 5662 5089
rect 5604 5030 5607 5082
rect 5659 5030 5662 5082
rect 5604 5018 5616 5030
rect 5650 5018 5662 5030
rect 5604 4966 5607 5018
rect 5659 4966 5662 5018
rect 5604 4954 5616 4966
rect 5650 4954 5662 4966
rect 5604 4902 5607 4954
rect 5659 4902 5662 4954
rect 5604 4890 5616 4902
rect 5650 4890 5662 4902
rect 5604 4838 5607 4890
rect 5659 4838 5662 4890
rect 5604 4835 5662 4838
rect 5604 4826 5616 4835
rect 5650 4826 5662 4835
rect 5604 4774 5607 4826
rect 5659 4774 5662 4826
rect 5604 4763 5662 4774
rect 5604 4762 5616 4763
rect 5650 4762 5662 4763
rect 5604 4710 5607 4762
rect 5659 4710 5662 4762
rect 5604 4698 5662 4710
rect 5604 4646 5607 4698
rect 5659 4646 5662 4698
rect 5604 4634 5662 4646
rect 5604 4582 5607 4634
rect 5659 4582 5662 4634
rect 5604 4570 5662 4582
rect 5604 4518 5607 4570
rect 5659 4518 5662 4570
rect 5604 4513 5616 4518
rect 5650 4513 5662 4518
rect 5604 4507 5662 4513
rect 348 4469 406 4507
rect 348 4435 360 4469
rect 394 4435 406 4469
rect 348 4397 406 4435
rect 348 4363 360 4397
rect 394 4363 406 4397
rect 348 4325 406 4363
rect 348 4291 360 4325
rect 394 4291 406 4325
tri 5972 4308 5998 4334 se
rect 5998 4308 6128 6136
rect 6183 5990 6189 6042
rect 6241 5990 6254 6042
rect 6306 5990 6319 6042
rect 6371 6033 6384 6042
rect 6436 6033 6448 6042
rect 6500 6033 6512 6042
rect 6564 6033 6576 6042
rect 6628 6033 6640 6042
rect 6376 5999 6384 6033
rect 6628 5999 6634 6033
rect 6371 5990 6384 5999
rect 6436 5990 6448 5999
rect 6500 5990 6512 5999
rect 6564 5990 6576 5999
rect 6628 5990 6640 5999
rect 6692 5990 6704 6042
rect 6756 5990 6768 6042
rect 6820 5990 6826 6042
rect 6183 5756 6189 5808
rect 6241 5756 6254 5808
rect 6306 5756 6319 5808
rect 6371 5799 6384 5808
rect 6436 5799 6448 5808
rect 6500 5799 6512 5808
rect 6564 5799 6576 5808
rect 6628 5799 6640 5808
rect 6376 5765 6384 5799
rect 6628 5765 6634 5799
rect 6371 5756 6384 5765
rect 6436 5756 6448 5765
rect 6500 5756 6512 5765
rect 6564 5756 6576 5765
rect 6628 5756 6640 5765
rect 6692 5756 6704 5808
rect 6756 5756 6768 5808
rect 6820 5756 6826 5808
rect 6460 5411 6518 5417
rect 6460 5402 6472 5411
rect 6506 5402 6518 5411
rect 6460 5350 6463 5402
rect 6515 5350 6518 5402
rect 6460 5339 6518 5350
rect 6460 5338 6472 5339
rect 6506 5338 6518 5339
rect 6460 5286 6463 5338
rect 6515 5286 6518 5338
rect 6460 5274 6518 5286
rect 6460 5222 6463 5274
rect 6515 5222 6518 5274
rect 6460 5210 6518 5222
rect 6460 5158 6463 5210
rect 6515 5158 6518 5210
rect 6460 5146 6518 5158
rect 6460 5094 6463 5146
rect 6515 5094 6518 5146
rect 6460 5089 6472 5094
rect 6506 5089 6518 5094
rect 6460 5082 6518 5089
rect 6460 5030 6463 5082
rect 6515 5030 6518 5082
rect 6460 5018 6472 5030
rect 6506 5018 6518 5030
rect 6460 4966 6463 5018
rect 6515 4966 6518 5018
rect 6460 4954 6472 4966
rect 6506 4954 6518 4966
rect 6460 4902 6463 4954
rect 6515 4902 6518 4954
rect 6460 4890 6472 4902
rect 6506 4890 6518 4902
rect 6460 4838 6463 4890
rect 6515 4838 6518 4890
rect 6460 4835 6518 4838
rect 6460 4826 6472 4835
rect 6506 4826 6518 4835
rect 6460 4774 6463 4826
rect 6515 4774 6518 4826
rect 6460 4763 6518 4774
rect 6460 4762 6472 4763
rect 6506 4762 6518 4763
rect 6460 4710 6463 4762
rect 6515 4710 6518 4762
rect 6460 4698 6518 4710
rect 6460 4646 6463 4698
rect 6515 4646 6518 4698
rect 6460 4634 6518 4646
rect 6460 4582 6463 4634
rect 6515 4582 6518 4634
rect 6460 4570 6518 4582
rect 6460 4518 6463 4570
rect 6515 4518 6518 4570
rect 6460 4513 6472 4518
rect 6506 4513 6518 4518
rect 6460 4507 6518 4513
tri 6128 4308 6154 4334 sw
tri 6828 4308 6854 4334 se
rect 6854 4308 6984 6444
rect 7054 5990 7060 6042
rect 7112 5990 7124 6042
rect 7176 5990 7188 6042
rect 7240 6033 7252 6042
rect 7304 6033 7316 6042
rect 7368 6033 7380 6042
rect 7432 6033 7444 6042
rect 7496 6033 7508 6042
rect 7247 5999 7252 6033
rect 7496 5999 7501 6033
rect 7240 5990 7252 5999
rect 7304 5990 7316 5999
rect 7368 5990 7380 5999
rect 7432 5990 7444 5999
rect 7496 5990 7508 5999
rect 7560 5990 7572 6042
rect 7624 5990 7630 6042
rect 7054 5756 7060 5808
rect 7112 5756 7124 5808
rect 7176 5756 7188 5808
rect 7240 5799 7252 5808
rect 7304 5799 7316 5808
rect 7368 5799 7380 5808
rect 7432 5799 7444 5808
rect 7496 5799 7508 5808
rect 7247 5765 7252 5799
rect 7496 5765 7501 5799
rect 7240 5756 7252 5765
rect 7304 5756 7316 5765
rect 7368 5756 7380 5765
rect 7432 5756 7444 5765
rect 7496 5756 7508 5765
rect 7560 5756 7572 5808
rect 7624 5756 7630 5808
rect 7316 5411 7374 5417
rect 7316 5402 7328 5411
rect 7362 5402 7374 5411
rect 7316 5350 7319 5402
rect 7371 5350 7374 5402
rect 7316 5339 7374 5350
rect 7316 5338 7328 5339
rect 7362 5338 7374 5339
rect 7316 5286 7319 5338
rect 7371 5286 7374 5338
rect 7316 5274 7374 5286
rect 7316 5222 7319 5274
rect 7371 5222 7374 5274
rect 7316 5210 7374 5222
rect 7316 5158 7319 5210
rect 7371 5158 7374 5210
rect 7316 5146 7374 5158
rect 7316 5094 7319 5146
rect 7371 5094 7374 5146
rect 7316 5089 7328 5094
rect 7362 5089 7374 5094
rect 7316 5082 7374 5089
rect 7316 5030 7319 5082
rect 7371 5030 7374 5082
rect 7316 5018 7328 5030
rect 7362 5018 7374 5030
rect 7316 4966 7319 5018
rect 7371 4966 7374 5018
rect 7316 4954 7328 4966
rect 7362 4954 7374 4966
rect 7316 4902 7319 4954
rect 7371 4902 7374 4954
rect 7316 4890 7328 4902
rect 7362 4890 7374 4902
rect 7316 4838 7319 4890
rect 7371 4838 7374 4890
rect 7316 4835 7374 4838
rect 7316 4826 7328 4835
rect 7362 4826 7374 4835
rect 7316 4774 7319 4826
rect 7371 4774 7374 4826
rect 7316 4763 7374 4774
rect 7316 4762 7328 4763
rect 7362 4762 7374 4763
rect 7316 4710 7319 4762
rect 7371 4710 7374 4762
rect 7316 4698 7374 4710
rect 7316 4646 7319 4698
rect 7371 4646 7374 4698
rect 7316 4634 7374 4646
rect 7316 4582 7319 4634
rect 7371 4582 7374 4634
rect 7316 4570 7374 4582
rect 7316 4518 7319 4570
rect 7371 4518 7374 4570
rect 7316 4513 7328 4518
rect 7362 4513 7374 4518
rect 7316 4507 7374 4513
tri 6984 4308 7010 4334 sw
tri 7684 4308 7710 4334 se
rect 7710 4308 7840 6752
rect 7917 5990 7923 6042
rect 7975 5990 7987 6042
rect 8039 5990 8051 6042
rect 8103 6033 8115 6042
rect 8167 6033 8179 6042
rect 8231 6033 8243 6042
rect 8295 6033 8307 6042
rect 8359 6033 8371 6042
rect 8110 5999 8115 6033
rect 8359 5999 8364 6033
rect 8103 5990 8115 5999
rect 8167 5990 8179 5999
rect 8231 5990 8243 5999
rect 8295 5990 8307 5999
rect 8359 5990 8371 5999
rect 8423 5990 8435 6042
rect 8487 5990 8493 6042
rect 7917 5756 7923 5808
rect 7975 5756 7987 5808
rect 8039 5756 8051 5808
rect 8103 5799 8115 5808
rect 8167 5799 8179 5808
rect 8231 5799 8243 5808
rect 8295 5799 8307 5808
rect 8359 5799 8371 5808
rect 8110 5765 8115 5799
rect 8359 5765 8364 5799
rect 8103 5756 8115 5765
rect 8167 5756 8179 5765
rect 8231 5756 8243 5765
rect 8295 5756 8307 5765
rect 8359 5756 8371 5765
rect 8423 5756 8435 5808
rect 8487 5756 8493 5808
rect 8172 5411 8230 5417
rect 8172 5402 8184 5411
rect 8218 5402 8230 5411
rect 8172 5350 8175 5402
rect 8227 5350 8230 5402
rect 8172 5339 8230 5350
rect 8172 5338 8184 5339
rect 8218 5338 8230 5339
rect 8172 5286 8175 5338
rect 8227 5286 8230 5338
rect 8172 5274 8230 5286
rect 8172 5222 8175 5274
rect 8227 5222 8230 5274
rect 8172 5210 8230 5222
rect 8172 5158 8175 5210
rect 8227 5158 8230 5210
rect 8172 5146 8230 5158
rect 8172 5094 8175 5146
rect 8227 5094 8230 5146
rect 8172 5089 8184 5094
rect 8218 5089 8230 5094
rect 8172 5082 8230 5089
rect 8172 5030 8175 5082
rect 8227 5030 8230 5082
rect 8172 5018 8184 5030
rect 8218 5018 8230 5030
rect 8172 4966 8175 5018
rect 8227 4966 8230 5018
rect 8172 4954 8184 4966
rect 8218 4954 8230 4966
rect 8172 4902 8175 4954
rect 8227 4902 8230 4954
rect 8172 4890 8184 4902
rect 8218 4890 8230 4902
rect 8172 4838 8175 4890
rect 8227 4838 8230 4890
rect 8172 4835 8230 4838
rect 8172 4826 8184 4835
rect 8218 4826 8230 4835
rect 8172 4774 8175 4826
rect 8227 4774 8230 4826
rect 8172 4763 8230 4774
rect 8172 4762 8184 4763
rect 8218 4762 8230 4763
rect 8172 4710 8175 4762
rect 8227 4710 8230 4762
rect 8172 4698 8230 4710
rect 8172 4646 8175 4698
rect 8227 4646 8230 4698
rect 8172 4634 8230 4646
rect 8172 4582 8175 4634
rect 8227 4582 8230 4634
rect 8172 4570 8230 4582
rect 8172 4518 8175 4570
rect 8227 4518 8230 4570
rect 8172 4513 8184 4518
rect 8218 4513 8230 4518
rect 8172 4507 8230 4513
tri 7840 4308 7866 4334 sw
tri 8540 4308 8566 4334 se
rect 8566 4308 8696 7060
rect 8775 5990 8781 6042
rect 8833 5990 8845 6042
rect 8897 5990 8909 6042
rect 8961 6033 8973 6042
rect 9025 6033 9037 6042
rect 9089 6033 9101 6042
rect 9153 6033 9165 6042
rect 9217 6033 9229 6042
rect 8968 5999 8973 6033
rect 9217 5999 9222 6033
rect 8961 5990 8973 5999
rect 9025 5990 9037 5999
rect 9089 5990 9101 5999
rect 9153 5990 9165 5999
rect 9217 5990 9229 5999
rect 9281 5990 9293 6042
rect 9345 5990 9351 6042
rect 8775 5756 8781 5808
rect 8833 5756 8845 5808
rect 8897 5756 8909 5808
rect 8961 5799 8973 5808
rect 9025 5799 9037 5808
rect 9089 5799 9101 5808
rect 9153 5799 9165 5808
rect 9217 5799 9229 5808
rect 8968 5765 8973 5799
rect 9217 5765 9222 5799
rect 8961 5756 8973 5765
rect 9025 5756 9037 5765
rect 9089 5756 9101 5765
rect 9153 5756 9165 5765
rect 9217 5756 9229 5765
rect 9281 5756 9293 5808
rect 9345 5756 9351 5808
rect 9028 5411 9086 5417
rect 9028 5402 9040 5411
rect 9074 5402 9086 5411
rect 9028 5350 9031 5402
rect 9083 5350 9086 5402
rect 9028 5339 9086 5350
rect 9028 5338 9040 5339
rect 9074 5338 9086 5339
rect 9028 5286 9031 5338
rect 9083 5286 9086 5338
rect 9028 5274 9086 5286
rect 9028 5222 9031 5274
rect 9083 5222 9086 5274
rect 9028 5210 9086 5222
rect 9028 5158 9031 5210
rect 9083 5158 9086 5210
rect 9028 5146 9086 5158
rect 9028 5094 9031 5146
rect 9083 5094 9086 5146
rect 9028 5089 9040 5094
rect 9074 5089 9086 5094
rect 9028 5082 9086 5089
rect 9028 5030 9031 5082
rect 9083 5030 9086 5082
rect 9028 5018 9040 5030
rect 9074 5018 9086 5030
rect 9028 4966 9031 5018
rect 9083 4966 9086 5018
rect 9028 4954 9040 4966
rect 9074 4954 9086 4966
rect 9028 4902 9031 4954
rect 9083 4902 9086 4954
rect 9028 4890 9040 4902
rect 9074 4890 9086 4902
rect 9028 4838 9031 4890
rect 9083 4838 9086 4890
rect 9028 4835 9086 4838
rect 9028 4826 9040 4835
rect 9074 4826 9086 4835
rect 9028 4774 9031 4826
rect 9083 4774 9086 4826
rect 9028 4763 9086 4774
rect 9028 4762 9040 4763
rect 9074 4762 9086 4763
rect 9028 4710 9031 4762
rect 9083 4710 9086 4762
rect 9028 4698 9086 4710
rect 9028 4646 9031 4698
rect 9083 4646 9086 4698
rect 9028 4634 9086 4646
rect 9028 4582 9031 4634
rect 9083 4582 9086 4634
rect 9028 4570 9086 4582
rect 9028 4518 9031 4570
rect 9083 4518 9086 4570
rect 9028 4513 9040 4518
rect 9074 4513 9086 4518
rect 9028 4507 9086 4513
tri 8696 4308 8722 4334 sw
tri 9396 4308 9422 4334 se
rect 9422 4308 9552 7368
rect 9613 5990 9619 6042
rect 9671 5990 9683 6042
rect 9735 5990 9747 6042
rect 9799 6033 9811 6042
rect 9863 6033 9875 6042
rect 9927 6033 9939 6042
rect 9991 6033 10003 6042
rect 10055 6033 10067 6042
rect 9806 5999 9811 6033
rect 10055 5999 10060 6033
rect 9799 5990 9811 5999
rect 9863 5990 9875 5999
rect 9927 5990 9939 5999
rect 9991 5990 10003 5999
rect 10055 5990 10067 5999
rect 10119 5990 10131 6042
rect 10183 5990 10189 6042
rect 9613 5756 9619 5808
rect 9671 5756 9683 5808
rect 9735 5756 9747 5808
rect 9799 5799 9811 5808
rect 9863 5799 9875 5808
rect 9927 5799 9939 5808
rect 9991 5799 10003 5808
rect 10055 5799 10067 5808
rect 9806 5765 9811 5799
rect 10055 5765 10060 5799
rect 9799 5756 9811 5765
rect 9863 5756 9875 5765
rect 9927 5756 9939 5765
rect 9991 5756 10003 5765
rect 10055 5756 10067 5765
rect 10119 5756 10131 5808
rect 10183 5756 10189 5808
rect 9884 5411 9942 5417
rect 9884 5402 9896 5411
rect 9930 5402 9942 5411
rect 9884 5350 9887 5402
rect 9939 5350 9942 5402
rect 9884 5339 9942 5350
rect 9884 5338 9896 5339
rect 9930 5338 9942 5339
rect 9884 5286 9887 5338
rect 9939 5286 9942 5338
rect 9884 5274 9942 5286
rect 9884 5222 9887 5274
rect 9939 5222 9942 5274
rect 9884 5210 9942 5222
rect 9884 5158 9887 5210
rect 9939 5158 9942 5210
rect 9884 5146 9942 5158
rect 9884 5094 9887 5146
rect 9939 5094 9942 5146
rect 9884 5089 9896 5094
rect 9930 5089 9942 5094
rect 9884 5082 9942 5089
rect 9884 5030 9887 5082
rect 9939 5030 9942 5082
rect 9884 5018 9896 5030
rect 9930 5018 9942 5030
rect 9884 4966 9887 5018
rect 9939 4966 9942 5018
rect 9884 4954 9896 4966
rect 9930 4954 9942 4966
rect 9884 4902 9887 4954
rect 9939 4902 9942 4954
rect 9884 4890 9896 4902
rect 9930 4890 9942 4902
rect 9884 4838 9887 4890
rect 9939 4838 9942 4890
rect 9884 4835 9942 4838
rect 9884 4826 9896 4835
rect 9930 4826 9942 4835
rect 9884 4774 9887 4826
rect 9939 4774 9942 4826
rect 9884 4763 9942 4774
rect 9884 4762 9896 4763
rect 9930 4762 9942 4763
rect 9884 4710 9887 4762
rect 9939 4710 9942 4762
rect 9884 4698 9942 4710
rect 9884 4646 9887 4698
rect 9939 4646 9942 4698
rect 9884 4634 9942 4646
rect 9884 4582 9887 4634
rect 9939 4582 9942 4634
rect 9884 4570 9942 4582
rect 9884 4518 9887 4570
rect 9939 4518 9942 4570
rect 9884 4513 9896 4518
rect 9930 4513 9942 4518
rect 9884 4507 9942 4513
tri 9552 4308 9578 4334 sw
tri 10252 4308 10278 4334 se
rect 10278 4308 10408 7676
tri 15167 7650 15193 7676 ne
rect 15193 7650 15241 7676
tri 15241 7650 15267 7676 sw
tri 15387 7650 15413 7676 ne
rect 15413 7650 15461 7676
tri 15461 7650 15487 7676 sw
rect 15725 7650 16033 7688
tri 15193 7616 15227 7650 ne
rect 15227 7616 15267 7650
tri 15267 7616 15301 7650 sw
tri 15413 7642 15421 7650 ne
rect 15421 7642 15487 7650
tri 15487 7642 15495 7650 sw
tri 15421 7616 15447 7642 ne
rect 15447 7616 15495 7642
tri 15495 7616 15521 7642 sw
rect 15725 7616 15733 7650
rect 15767 7616 15819 7650
rect 15853 7616 15905 7650
rect 15939 7616 15991 7650
rect 16025 7616 16033 7650
tri 15227 7578 15265 7616 ne
rect 15265 7578 15301 7616
tri 15301 7578 15339 7616 sw
tri 15447 7578 15485 7616 ne
rect 15485 7578 15521 7616
tri 15521 7578 15559 7616 sw
rect 15725 7578 16033 7616
tri 15265 7576 15267 7578 ne
rect 15267 7576 15339 7578
tri 15339 7576 15341 7578 sw
tri 15485 7576 15487 7578 ne
rect 15487 7576 15559 7578
tri 15559 7576 15561 7578 sw
tri 15267 7574 15269 7576 ne
rect 15269 7574 15341 7576
tri 15341 7574 15343 7576 sw
tri 15487 7574 15489 7576 ne
rect 15489 7574 15561 7576
tri 15561 7574 15563 7576 sw
rect 12870 7565 15141 7574
rect 12870 7531 12882 7565
rect 12916 7531 12954 7565
rect 12988 7544 15141 7565
tri 15141 7544 15171 7574 sw
tri 15269 7544 15299 7574 ne
rect 15299 7544 15343 7574
tri 15343 7544 15373 7574 sw
tri 15489 7568 15495 7574 ne
rect 15495 7568 15563 7574
tri 15563 7568 15569 7574 sw
tri 15495 7544 15519 7568 ne
rect 15519 7544 15569 7568
tri 15569 7544 15593 7568 sw
rect 15725 7544 15733 7578
rect 15767 7544 15819 7578
rect 15853 7544 15905 7578
rect 15939 7544 15991 7578
rect 16025 7544 16033 7578
rect 12988 7531 15171 7544
rect 12870 7528 15171 7531
tri 15171 7528 15187 7544 sw
tri 15299 7528 15315 7544 ne
rect 15315 7528 15373 7544
rect 12870 7522 15187 7528
tri 15187 7522 15193 7528 sw
tri 15315 7522 15321 7528 ne
rect 15321 7522 15373 7528
tri 15373 7522 15395 7544 sw
tri 15519 7522 15541 7544 ne
rect 15541 7522 15593 7544
tri 15593 7522 15615 7544 sw
tri 15119 7506 15135 7522 ne
rect 15135 7506 15193 7522
tri 15193 7506 15209 7522 sw
tri 15321 7506 15337 7522 ne
rect 15337 7506 15395 7522
tri 15395 7506 15411 7522 sw
tri 15541 7506 15557 7522 ne
rect 15557 7506 15615 7522
tri 15615 7506 15631 7522 sw
rect 15725 7506 16033 7544
tri 15135 7472 15169 7506 ne
rect 15169 7502 15209 7506
tri 15209 7502 15213 7506 sw
tri 15337 7502 15341 7506 ne
rect 15341 7502 15411 7506
tri 15411 7502 15415 7506 sw
tri 15557 7502 15561 7506 ne
rect 15561 7502 15631 7506
tri 15631 7502 15635 7506 sw
rect 15169 7472 15213 7502
tri 15213 7472 15243 7502 sw
tri 15341 7472 15371 7502 ne
rect 15371 7472 15415 7502
tri 15415 7472 15445 7502 sw
tri 15561 7494 15569 7502 ne
rect 15569 7494 15635 7502
tri 15635 7494 15643 7502 sw
tri 15569 7472 15591 7494 ne
tri 15169 7454 15187 7472 ne
rect 15187 7454 15243 7472
tri 15243 7454 15261 7472 sw
tri 15371 7454 15389 7472 ne
rect 15389 7454 15445 7472
tri 15187 7434 15207 7454 ne
rect 15207 7434 15261 7454
tri 15261 7434 15281 7454 sw
tri 15389 7434 15409 7454 ne
rect 15409 7434 15445 7454
tri 15445 7434 15483 7472 sw
tri 15207 7420 15221 7434 ne
rect 15221 7428 15281 7434
tri 15281 7428 15287 7434 sw
tri 15409 7428 15415 7434 ne
rect 15415 7428 15483 7434
tri 15483 7428 15489 7434 sw
rect 15221 7420 15287 7428
tri 15287 7420 15295 7428 sw
tri 15415 7420 15423 7428 ne
rect 15423 7420 15489 7428
tri 15489 7420 15497 7428 sw
rect 12870 7411 15075 7420
rect 12870 7377 12882 7411
rect 12916 7377 12954 7411
rect 12988 7400 15075 7411
tri 15075 7400 15095 7420 sw
tri 15221 7400 15241 7420 ne
rect 15241 7400 15295 7420
tri 15295 7400 15315 7420 sw
tri 15423 7400 15443 7420 ne
rect 15443 7400 15497 7420
tri 15497 7400 15517 7420 sw
rect 12988 7388 15095 7400
tri 15095 7388 15107 7400 sw
tri 15241 7388 15253 7400 ne
rect 15253 7388 15315 7400
tri 15315 7388 15327 7400 sw
tri 15443 7388 15455 7400 ne
rect 15455 7388 15517 7400
tri 15517 7388 15529 7400 sw
rect 12988 7377 15107 7388
rect 12870 7368 15107 7377
tri 15107 7368 15127 7388 sw
tri 15253 7380 15261 7388 ne
rect 15261 7380 15327 7388
tri 15327 7380 15335 7388 sw
tri 15455 7380 15463 7388 ne
rect 15463 7380 15529 7388
tri 15261 7368 15273 7380 ne
rect 15273 7368 15335 7380
tri 15335 7368 15347 7380 sw
tri 15463 7368 15475 7380 ne
rect 15475 7368 15529 7380
tri 15529 7368 15549 7388 sw
tri 15053 7362 15059 7368 ne
rect 15059 7362 15127 7368
tri 15127 7362 15133 7368 sw
tri 15273 7362 15279 7368 ne
rect 15279 7362 15347 7368
tri 15347 7362 15353 7368 sw
tri 15475 7362 15481 7368 ne
rect 15481 7362 15549 7368
tri 15549 7362 15555 7368 sw
tri 15059 7328 15093 7362 ne
rect 15093 7328 15133 7362
tri 15133 7328 15167 7362 sw
tri 15279 7328 15313 7362 ne
rect 15313 7354 15353 7362
tri 15353 7354 15361 7362 sw
tri 15481 7354 15489 7362 ne
rect 15489 7354 15555 7362
tri 15555 7354 15563 7362 sw
rect 15313 7332 15361 7354
tri 15361 7332 15383 7354 sw
tri 15489 7332 15511 7354 ne
rect 15313 7328 15383 7332
tri 15383 7328 15387 7332 sw
tri 15093 7314 15107 7328 ne
rect 15107 7314 15167 7328
tri 15167 7314 15181 7328 sw
tri 15313 7314 15327 7328 ne
rect 15327 7314 15387 7328
tri 15387 7314 15401 7328 sw
tri 15107 7290 15131 7314 ne
rect 15131 7290 15181 7314
tri 15181 7290 15205 7314 sw
tri 15327 7306 15335 7314 ne
rect 15335 7306 15401 7314
tri 15401 7306 15409 7314 sw
tri 15335 7290 15351 7306 ne
rect 15351 7290 15409 7306
tri 15409 7290 15425 7306 sw
tri 15131 7266 15155 7290 ne
rect 15155 7266 15205 7290
tri 15205 7266 15229 7290 sw
tri 15351 7266 15375 7290 ne
rect 15375 7266 15425 7290
tri 15425 7266 15449 7290 sw
rect 12870 7257 15009 7266
rect 12870 7223 12882 7257
rect 12916 7223 12954 7257
rect 12988 7256 15009 7257
tri 15009 7256 15019 7266 sw
tri 15155 7256 15165 7266 ne
rect 15165 7256 15229 7266
tri 15229 7256 15239 7266 sw
tri 15375 7256 15385 7266 ne
rect 15385 7256 15449 7266
tri 15449 7256 15459 7266 sw
rect 12988 7248 15019 7256
tri 15019 7248 15027 7256 sw
tri 15165 7248 15173 7256 ne
rect 15173 7248 15239 7256
rect 12988 7240 15027 7248
tri 15027 7240 15035 7248 sw
tri 15173 7240 15181 7248 ne
rect 15181 7240 15239 7248
tri 15239 7240 15255 7256 sw
tri 15385 7240 15401 7256 ne
rect 15401 7240 15459 7256
tri 15459 7240 15475 7256 sw
rect 12988 7223 15035 7240
rect 12870 7218 15035 7223
tri 15035 7218 15057 7240 sw
tri 15181 7218 15203 7240 ne
rect 15203 7218 15255 7240
tri 15255 7218 15277 7240 sw
tri 15401 7232 15409 7240 ne
rect 15409 7232 15475 7240
tri 15475 7232 15483 7240 sw
tri 15409 7218 15423 7232 ne
rect 15423 7218 15483 7232
rect 12870 7214 15057 7218
tri 15057 7214 15061 7218 sw
tri 15203 7214 15207 7218 ne
rect 15207 7214 15277 7218
tri 15277 7214 15281 7218 sw
tri 15423 7214 15427 7218 ne
rect 15427 7214 15483 7218
tri 14987 7184 15017 7214 ne
rect 15017 7184 15061 7214
tri 15061 7184 15091 7214 sw
tri 15207 7184 15237 7214 ne
rect 15237 7184 15281 7214
tri 15281 7184 15311 7214 sw
tri 15427 7210 15431 7214 ne
tri 15017 7174 15027 7184 ne
rect 15027 7174 15091 7184
tri 15091 7174 15101 7184 sw
tri 15237 7174 15247 7184 ne
rect 15247 7174 15311 7184
tri 15027 7146 15055 7174 ne
rect 15055 7166 15101 7174
tri 15101 7166 15109 7174 sw
tri 15247 7166 15255 7174 ne
rect 15255 7166 15311 7174
tri 15311 7166 15329 7184 sw
rect 15055 7146 15109 7166
tri 15109 7146 15129 7166 sw
tri 15255 7146 15275 7166 ne
rect 15275 7146 15329 7166
tri 15329 7146 15349 7166 sw
tri 15055 7112 15089 7146 ne
rect 15089 7112 15129 7146
tri 15129 7112 15163 7146 sw
tri 15275 7112 15309 7146 ne
rect 15309 7112 15349 7146
tri 15349 7112 15383 7146 sw
rect 12870 7108 14943 7112
tri 14943 7108 14947 7112 sw
tri 15089 7108 15093 7112 ne
rect 15093 7108 15163 7112
rect 12870 7103 14947 7108
rect 12870 7069 12882 7103
rect 12916 7069 12954 7103
rect 12988 7100 14947 7103
tri 14947 7100 14955 7108 sw
tri 15093 7100 15101 7108 ne
rect 15101 7100 15163 7108
tri 15163 7100 15175 7112 sw
tri 15309 7100 15321 7112 ne
rect 15321 7100 15383 7112
rect 12988 7074 14955 7100
tri 14955 7074 14981 7100 sw
tri 15101 7074 15127 7100 ne
rect 15127 7092 15175 7100
tri 15175 7092 15183 7100 sw
tri 15321 7092 15329 7100 ne
rect 15329 7092 15383 7100
tri 15383 7092 15403 7112 sw
rect 15127 7074 15183 7092
tri 15183 7074 15201 7092 sw
tri 15329 7074 15347 7092 ne
rect 15347 7074 15403 7092
rect 12988 7069 14981 7074
rect 12870 7060 14981 7069
tri 14981 7060 14995 7074 sw
tri 15127 7060 15141 7074 ne
rect 15141 7070 15201 7074
tri 15201 7070 15205 7074 sw
tri 15347 7070 15351 7074 ne
rect 15141 7060 15205 7070
tri 15205 7060 15215 7070 sw
tri 14921 7040 14941 7060 ne
rect 14941 7040 14995 7060
tri 14995 7040 15015 7060 sw
tri 15141 7040 15161 7060 ne
rect 15161 7040 15215 7060
tri 15215 7040 15235 7060 sw
tri 14941 7034 14947 7040 ne
rect 14947 7034 15015 7040
tri 15015 7034 15021 7040 sw
tri 15161 7034 15167 7040 ne
rect 15167 7034 15235 7040
tri 14947 7002 14979 7034 ne
rect 14979 7026 15021 7034
tri 15021 7026 15029 7034 sw
tri 15167 7026 15175 7034 ne
rect 15175 7026 15235 7034
tri 15235 7026 15249 7040 sw
rect 14979 7002 15029 7026
tri 15029 7002 15053 7026 sw
tri 15175 7002 15199 7026 ne
rect 15199 7002 15249 7026
tri 15249 7002 15273 7026 sw
tri 14979 6968 15013 7002 ne
rect 15013 6968 15053 7002
tri 15053 6968 15087 7002 sw
tri 15199 6968 15233 7002 ne
rect 15233 6968 15273 7002
tri 15273 6968 15307 7002 sw
tri 15013 6960 15021 6968 ne
rect 15021 6960 15087 6968
tri 15087 6960 15095 6968 sw
tri 15233 6960 15241 6968 ne
rect 15241 6960 15307 6968
tri 15021 6958 15023 6960 ne
rect 15023 6958 15095 6960
tri 15095 6958 15097 6960 sw
tri 15241 6958 15243 6960 ne
rect 15243 6958 15307 6960
tri 15307 6958 15317 6968 sw
rect 12870 6949 14877 6958
rect 12870 6915 12882 6949
rect 12916 6915 12954 6949
rect 12988 6930 14877 6949
tri 14877 6930 14905 6958 sw
tri 15023 6930 15051 6958 ne
rect 15051 6952 15097 6958
tri 15097 6952 15103 6958 sw
tri 15243 6952 15249 6958 ne
rect 15249 6952 15317 6958
tri 15317 6952 15323 6958 sw
rect 15051 6930 15103 6952
tri 15103 6930 15125 6952 sw
tri 15249 6930 15271 6952 ne
rect 12988 6915 14905 6930
rect 12870 6906 14905 6915
tri 14905 6906 14929 6930 sw
tri 15051 6906 15075 6930 ne
rect 15075 6906 15125 6930
tri 15125 6906 15149 6930 sw
tri 14855 6896 14865 6906 ne
rect 14865 6896 14929 6906
tri 14929 6896 14939 6906 sw
tri 15075 6896 15085 6906 ne
rect 15085 6896 15149 6906
tri 15149 6896 15159 6906 sw
tri 14865 6894 14867 6896 ne
rect 14867 6894 14939 6896
tri 14939 6894 14941 6896 sw
tri 15085 6894 15087 6896 ne
rect 15087 6894 15159 6896
tri 14867 6884 14877 6894 ne
rect 14877 6886 14941 6894
tri 14941 6886 14949 6894 sw
tri 15087 6886 15095 6894 ne
rect 15095 6886 15159 6894
tri 15159 6886 15169 6896 sw
rect 14877 6884 14949 6886
tri 14877 6858 14903 6884 ne
rect 14903 6858 14949 6884
tri 14949 6858 14977 6886 sw
tri 15095 6858 15123 6886 ne
rect 15123 6858 15169 6886
tri 15169 6858 15197 6886 sw
tri 14903 6824 14937 6858 ne
rect 14937 6824 14977 6858
tri 14977 6824 15011 6858 sw
tri 15123 6824 15157 6858 ne
rect 15157 6824 15197 6858
tri 15197 6824 15231 6858 sw
tri 14937 6820 14941 6824 ne
rect 14941 6820 15011 6824
tri 15011 6820 15015 6824 sw
tri 15157 6820 15161 6824 ne
rect 15161 6820 15231 6824
tri 14941 6804 14957 6820 ne
rect 14957 6812 15015 6820
tri 15015 6812 15023 6820 sw
tri 15161 6812 15169 6820 ne
rect 15169 6812 15231 6820
tri 15231 6812 15243 6824 sw
rect 14957 6804 15023 6812
tri 15023 6804 15031 6812 sw
tri 15169 6804 15177 6812 ne
rect 15177 6804 15243 6812
rect 12870 6795 14811 6804
rect 12870 6761 12882 6795
rect 12916 6761 12954 6795
rect 12988 6786 14811 6795
tri 14811 6786 14829 6804 sw
tri 14957 6786 14975 6804 ne
rect 14975 6790 15031 6804
tri 15031 6790 15045 6804 sw
tri 15177 6790 15191 6804 ne
rect 14975 6786 15045 6790
tri 15045 6786 15049 6790 sw
rect 12988 6761 14829 6786
rect 12870 6754 14829 6761
tri 14829 6754 14861 6786 sw
tri 14975 6754 15007 6786 ne
rect 15007 6754 15049 6786
rect 12870 6752 14861 6754
tri 14861 6752 14863 6754 sw
tri 15007 6752 15009 6754 ne
rect 15009 6752 15049 6754
tri 15049 6752 15083 6786 sw
tri 14789 6714 14827 6752 ne
rect 14827 6746 14863 6752
tri 14863 6746 14869 6752 sw
tri 15009 6746 15015 6752 ne
rect 15015 6746 15083 6752
tri 15083 6746 15089 6752 sw
rect 14827 6714 14869 6746
tri 14869 6714 14901 6746 sw
tri 15015 6714 15047 6746 ne
rect 15047 6714 15089 6746
tri 15089 6714 15121 6746 sw
tri 14827 6680 14861 6714 ne
rect 14861 6680 14901 6714
tri 14901 6680 14935 6714 sw
tri 15047 6680 15081 6714 ne
rect 15081 6680 15121 6714
tri 15121 6680 15155 6714 sw
tri 14861 6650 14891 6680 ne
rect 14891 6672 14935 6680
tri 14935 6672 14943 6680 sw
tri 15081 6672 15089 6680 ne
rect 15089 6672 15155 6680
tri 15155 6672 15163 6680 sw
rect 14891 6650 14943 6672
tri 14943 6650 14965 6672 sw
tri 15089 6650 15111 6672 ne
rect 12870 6642 14745 6650
tri 14745 6642 14753 6650 sw
tri 14891 6642 14899 6650 ne
rect 14899 6642 14965 6650
tri 14965 6642 14973 6650 sw
rect 12870 6641 14753 6642
rect 12870 6607 12882 6641
rect 12916 6607 12954 6641
rect 12988 6614 14753 6641
tri 14753 6614 14781 6642 sw
tri 14899 6614 14927 6642 ne
rect 14927 6614 14973 6642
rect 12988 6608 14781 6614
tri 14781 6608 14787 6614 sw
tri 14927 6608 14933 6614 ne
rect 14933 6608 14973 6614
tri 14973 6608 15007 6642 sw
rect 12988 6607 14787 6608
rect 12870 6606 14787 6607
tri 14787 6606 14789 6608 sw
tri 14933 6606 14935 6608 ne
rect 14935 6606 15007 6608
tri 15007 6606 15009 6608 sw
rect 12870 6598 14789 6606
tri 14789 6598 14797 6606 sw
tri 14935 6598 14943 6606 ne
rect 14943 6598 15009 6606
tri 15009 6598 15017 6606 sw
tri 14723 6570 14751 6598 ne
rect 14751 6570 14797 6598
tri 14797 6570 14825 6598 sw
tri 14943 6570 14971 6598 ne
rect 14971 6570 15017 6598
tri 15017 6570 15045 6598 sw
tri 14751 6540 14781 6570 ne
rect 14781 6540 14825 6570
tri 14825 6540 14855 6570 sw
tri 14971 6540 15001 6570 ne
rect 15001 6540 15045 6570
tri 14781 6536 14785 6540 ne
rect 14785 6536 14855 6540
tri 14855 6536 14859 6540 sw
tri 15001 6536 15005 6540 ne
rect 15005 6536 15045 6540
tri 15045 6536 15079 6570 sw
tri 14785 6498 14823 6536 ne
rect 14823 6532 14859 6536
tri 14859 6532 14863 6536 sw
tri 15005 6532 15009 6536 ne
rect 15009 6532 15079 6536
tri 15079 6532 15083 6536 sw
rect 14823 6510 14863 6532
tri 14863 6510 14885 6532 sw
tri 15009 6510 15031 6532 ne
rect 14823 6498 14885 6510
tri 14885 6498 14897 6510 sw
tri 14823 6496 14825 6498 ne
rect 14825 6496 14897 6498
tri 14897 6496 14899 6498 sw
rect 12870 6487 14780 6496
rect 12870 6453 12882 6487
rect 12916 6453 12954 6487
rect 12988 6472 14780 6487
tri 14780 6472 14804 6496 sw
tri 14825 6472 14849 6496 ne
rect 14849 6472 14899 6496
rect 12988 6466 14804 6472
tri 14804 6466 14810 6472 sw
tri 14849 6466 14855 6472 ne
rect 14855 6466 14899 6472
tri 14899 6466 14929 6496 sw
rect 12988 6464 14810 6466
tri 14810 6464 14812 6466 sw
tri 14855 6464 14857 6466 ne
rect 14857 6464 14929 6466
tri 14929 6464 14931 6466 sw
rect 12988 6453 14812 6464
rect 12870 6444 14812 6453
tri 14812 6444 14832 6464 sw
tri 14857 6444 14877 6464 ne
rect 14877 6444 14931 6464
tri 14931 6444 14951 6464 sw
tri 14758 6427 14775 6444 ne
rect 14775 6427 14832 6444
tri 14832 6427 14849 6444 sw
tri 14877 6427 14894 6444 ne
rect 14894 6427 14951 6444
tri 14775 6426 14776 6427 ne
rect 14776 6426 14849 6427
tri 14849 6426 14850 6427 sw
tri 14894 6426 14895 6427 ne
rect 14895 6426 14951 6427
tri 14951 6426 14969 6444 sw
tri 14776 6422 14780 6426 ne
rect 14780 6422 14850 6426
tri 14780 6392 14810 6422 ne
rect 14810 6398 14850 6422
tri 14850 6398 14878 6426 sw
tri 14895 6398 14923 6426 ne
rect 14923 6398 14969 6426
rect 14810 6392 14878 6398
tri 14878 6392 14884 6398 sw
tri 14923 6392 14929 6398 ne
rect 14929 6392 14969 6398
tri 14969 6392 15003 6426 sw
tri 14810 6354 14848 6392 ne
rect 14848 6370 14884 6392
tri 14884 6370 14906 6392 sw
tri 14929 6370 14951 6392 ne
rect 14848 6354 14906 6370
tri 14906 6354 14922 6370 sw
tri 14848 6353 14849 6354 ne
rect 14849 6353 14922 6354
tri 14922 6353 14923 6354 sw
tri 14849 6342 14860 6353 ne
rect 14860 6342 14923 6353
rect 12870 6333 14812 6342
rect 12870 6299 12882 6333
rect 12916 6299 12954 6333
rect 12988 6331 14812 6333
tri 14812 6331 14823 6342 sw
tri 14860 6331 14871 6342 ne
rect 12988 6320 14823 6331
tri 14823 6320 14834 6331 sw
rect 12988 6311 14834 6320
tri 14834 6311 14843 6320 sw
rect 12988 6299 14843 6311
rect 12870 6290 14843 6299
tri 14757 6282 14765 6290 ne
rect 14765 6282 14843 6290
tri 14765 6256 14791 6282 ne
rect 12870 6179 14698 6188
rect 12870 6145 12882 6179
rect 12916 6145 12954 6179
rect 12988 6176 14698 6179
tri 14698 6176 14710 6188 sw
rect 12988 6145 14710 6176
rect 12870 6144 14710 6145
tri 14710 6144 14742 6176 sw
rect 12870 6136 14742 6144
tri 14640 6104 14672 6136 ne
rect 14672 6104 14742 6136
tri 14672 6086 14690 6104 ne
rect 10459 5990 10465 6042
rect 10517 5990 10529 6042
rect 10581 5990 10593 6042
rect 10645 5990 10657 6042
rect 10709 6033 10721 6042
rect 10773 6033 10785 6042
rect 10837 6033 10849 6042
rect 10901 6033 10913 6042
rect 10965 6033 10977 6042
rect 10716 5999 10721 6033
rect 10965 5999 10970 6033
rect 10709 5990 10721 5999
rect 10773 5990 10785 5999
rect 10837 5990 10849 5999
rect 10901 5990 10913 5999
rect 10965 5990 10977 5999
rect 11029 5990 11041 6042
rect 11093 5990 11105 6042
rect 11157 5990 11169 6042
rect 11221 5990 11233 6042
rect 11285 6033 11297 6042
rect 11349 6033 11361 6042
rect 11413 6033 11425 6042
rect 11477 6033 11489 6042
rect 11541 6033 11553 6042
rect 11292 5999 11297 6033
rect 11541 5999 11546 6033
rect 11285 5990 11297 5999
rect 11349 5990 11361 5999
rect 11413 5990 11425 5999
rect 11477 5990 11489 5999
rect 11541 5990 11553 5999
rect 11605 5990 11617 6042
rect 11669 5990 11681 6042
rect 11733 5990 11745 6042
rect 11797 5990 11809 6042
rect 11861 6033 11873 6042
rect 11925 6033 11937 6042
rect 11989 6033 12001 6042
rect 12053 6033 12065 6042
rect 12117 6033 12129 6042
rect 11868 5999 11873 6033
rect 12117 5999 12122 6033
rect 11861 5990 11873 5999
rect 11925 5990 11937 5999
rect 11989 5990 12001 5999
rect 12053 5990 12065 5999
rect 12117 5990 12129 5999
rect 12181 5990 12193 6042
rect 12245 5990 12257 6042
rect 12309 5990 12321 6042
rect 12373 5990 12385 6042
rect 12437 6033 12449 6042
rect 12501 6033 12513 6042
rect 12565 6033 12577 6042
rect 12629 6033 12641 6042
rect 12693 6033 12705 6042
rect 12444 5999 12449 6033
rect 12693 5999 12698 6033
rect 12437 5990 12449 5999
rect 12501 5990 12513 5999
rect 12565 5990 12577 5999
rect 12629 5990 12641 5999
rect 12693 5990 12705 5999
rect 12757 5990 12769 6042
rect 12821 5990 12833 6042
rect 12885 5990 12897 6042
rect 12949 5990 12961 6042
rect 13013 6033 13025 6042
rect 13077 6033 13089 6042
rect 13020 5999 13025 6033
rect 13013 5990 13025 5999
rect 13077 5990 13089 5999
rect 13141 5990 13153 6042
rect 13205 5990 13217 6042
rect 13269 6033 13281 6042
rect 13333 6033 13345 6042
rect 13397 6033 13409 6042
rect 13461 6033 13473 6042
rect 13274 5999 13281 6033
rect 13461 5999 13465 6033
rect 13269 5990 13281 5999
rect 13333 5990 13345 5999
rect 13397 5990 13409 5999
rect 13461 5990 13473 5999
rect 13525 5990 13537 6042
rect 13589 5990 13601 6042
rect 13653 5990 13665 6042
rect 13717 6033 13729 6042
rect 13781 6033 13793 6042
rect 13845 6033 13857 6042
rect 13909 6033 13921 6042
rect 13724 5999 13729 6033
rect 13909 5999 13915 6033
rect 13717 5990 13729 5999
rect 13781 5990 13793 5999
rect 13845 5990 13857 5999
rect 13909 5990 13921 5999
rect 13973 5990 13985 6042
rect 14037 5990 14049 6042
rect 14101 5990 14114 6042
rect 14166 6033 14179 6042
rect 14231 6033 14244 6042
rect 14296 6033 14309 6042
rect 14361 6033 14374 6042
rect 14174 5999 14179 6033
rect 14361 5999 14365 6033
rect 14166 5990 14179 5999
rect 14231 5990 14244 5999
rect 14296 5990 14309 5999
rect 14361 5990 14374 5999
rect 14426 5990 14439 6042
rect 14491 5990 14504 6042
rect 14556 5990 14562 6042
rect 10986 5910 10992 5962
rect 11044 5910 11056 5962
rect 11108 5910 11114 5962
rect 11384 5910 11390 5962
rect 11442 5910 11454 5962
rect 11506 5960 12075 5962
tri 12075 5960 12077 5962 sw
rect 11506 5922 12077 5960
tri 12077 5922 12115 5960 sw
tri 14670 5922 14690 5942 se
rect 14690 5922 14742 6104
rect 11506 5910 12115 5922
rect 10470 5756 10476 5808
rect 10528 5756 10540 5808
rect 10592 5799 10604 5808
rect 10656 5799 10668 5808
rect 10720 5799 10732 5808
rect 10784 5799 10796 5808
rect 10848 5799 10860 5808
rect 10593 5765 10604 5799
rect 10665 5765 10668 5799
rect 10592 5756 10604 5765
rect 10656 5756 10668 5765
rect 10720 5756 10732 5765
rect 10784 5756 10796 5765
rect 10848 5756 10860 5765
rect 10912 5756 10918 5808
tri 10808 5744 10820 5756 ne
rect 10820 5744 10918 5756
tri 10820 5734 10830 5744 ne
rect 10830 5734 10918 5744
tri 10830 5710 10854 5734 ne
rect 10854 5710 10918 5734
tri 10854 5704 10860 5710 ne
rect 10860 5676 10872 5710
rect 10906 5676 10918 5710
rect 10860 5638 10918 5676
rect 10860 5604 10872 5638
rect 10906 5604 10918 5638
rect 10860 5566 10918 5604
rect 10860 5532 10872 5566
rect 10906 5532 10918 5566
rect 10860 5494 10918 5532
rect 10860 5460 10872 5494
rect 10906 5460 10918 5494
rect 10860 5422 10918 5460
rect 10740 5411 10798 5417
rect 10740 5402 10752 5411
rect 10786 5402 10798 5411
rect 10740 5350 10743 5402
rect 10795 5350 10798 5402
rect 10740 5339 10798 5350
rect 10740 5338 10752 5339
rect 10786 5338 10798 5339
rect 10740 5286 10743 5338
rect 10795 5286 10798 5338
rect 10740 5274 10798 5286
rect 10740 5222 10743 5274
rect 10795 5222 10798 5274
rect 10740 5210 10798 5222
rect 10740 5158 10743 5210
rect 10795 5158 10798 5210
rect 10740 5146 10798 5158
rect 10740 5094 10743 5146
rect 10795 5094 10798 5146
rect 10740 5089 10752 5094
rect 10786 5089 10798 5094
rect 10740 5082 10798 5089
rect 10740 5030 10743 5082
rect 10795 5030 10798 5082
rect 10740 5018 10752 5030
rect 10786 5018 10798 5030
rect 10740 4966 10743 5018
rect 10795 4966 10798 5018
rect 10740 4954 10752 4966
rect 10786 4954 10798 4966
rect 10740 4902 10743 4954
rect 10795 4902 10798 4954
rect 10740 4890 10752 4902
rect 10786 4890 10798 4902
rect 10740 4838 10743 4890
rect 10795 4838 10798 4890
rect 10740 4835 10798 4838
rect 10740 4826 10752 4835
rect 10786 4826 10798 4835
rect 10740 4774 10743 4826
rect 10795 4774 10798 4826
rect 10740 4763 10798 4774
rect 10740 4762 10752 4763
rect 10786 4762 10798 4763
rect 10740 4710 10743 4762
rect 10795 4710 10798 4762
rect 10740 4698 10798 4710
rect 10740 4646 10743 4698
rect 10795 4646 10798 4698
rect 10740 4634 10798 4646
rect 10740 4582 10743 4634
rect 10795 4582 10798 4634
rect 10740 4570 10798 4582
rect 10740 4518 10743 4570
rect 10795 4518 10798 4570
rect 10740 4513 10752 4518
rect 10786 4513 10798 4518
rect 10740 4507 10798 4513
rect 10860 5402 10872 5422
rect 10906 5402 10918 5422
rect 10860 5350 10863 5402
rect 10915 5350 10918 5402
rect 10860 5338 10872 5350
rect 10906 5338 10918 5350
rect 10860 5286 10863 5338
rect 10915 5286 10918 5338
rect 10860 5278 10918 5286
rect 10860 5274 10872 5278
rect 10906 5274 10918 5278
rect 10860 5222 10863 5274
rect 10915 5222 10918 5274
rect 10860 5210 10918 5222
rect 10860 5158 10863 5210
rect 10915 5158 10918 5210
rect 10860 5146 10918 5158
rect 10860 5094 10863 5146
rect 10915 5094 10918 5146
rect 10860 5082 10918 5094
rect 10860 5030 10863 5082
rect 10915 5030 10918 5082
rect 10860 5028 10872 5030
rect 10906 5028 10918 5030
rect 10860 5018 10918 5028
rect 10860 4966 10863 5018
rect 10915 4966 10918 5018
rect 10860 4956 10872 4966
rect 10906 4956 10918 4966
rect 10860 4954 10918 4956
rect 10860 4902 10863 4954
rect 10915 4902 10918 4954
rect 10860 4890 10872 4902
rect 10906 4890 10918 4902
rect 10860 4838 10863 4890
rect 10915 4838 10918 4890
rect 10860 4826 10872 4838
rect 10906 4826 10918 4838
rect 10860 4774 10863 4826
rect 10915 4774 10918 4826
rect 10860 4762 10872 4774
rect 10906 4762 10918 4774
rect 10860 4710 10863 4762
rect 10915 4710 10918 4762
rect 10860 4702 10918 4710
rect 10860 4698 10872 4702
rect 10906 4698 10918 4702
rect 10860 4646 10863 4698
rect 10915 4646 10918 4698
rect 10860 4634 10918 4646
rect 10860 4582 10863 4634
rect 10915 4582 10918 4634
rect 10860 4570 10918 4582
rect 10860 4518 10863 4570
rect 10915 4518 10918 4570
rect 10860 4486 10918 4518
rect 10860 4452 10872 4486
rect 10906 4452 10918 4486
rect 10860 4414 10918 4452
rect 10860 4380 10872 4414
rect 10906 4380 10918 4414
rect 10860 4342 10918 4380
tri 10408 4308 10434 4334 sw
rect 10860 4308 10872 4342
rect 10906 4308 10918 4342
tri 5968 4304 5972 4308 se
rect 5972 4304 6154 4308
tri 6154 4304 6158 4308 sw
tri 6824 4304 6828 4308 se
rect 6828 4304 7010 4308
tri 7010 4304 7014 4308 sw
tri 7680 4304 7684 4308 se
rect 7684 4304 7866 4308
tri 7866 4304 7870 4308 sw
tri 8536 4304 8540 4308 se
rect 8540 4304 8722 4308
tri 8722 4304 8726 4308 sw
tri 9392 4304 9396 4308 se
rect 9396 4304 9578 4308
tri 9578 4304 9582 4308 sw
tri 10248 4304 10252 4308 se
rect 10252 4304 10434 4308
tri 10434 4304 10438 4308 sw
rect 348 4253 406 4291
tri 5939 4275 5968 4304 se
rect 5968 4275 6158 4304
tri 6158 4275 6187 4304 sw
tri 6795 4275 6824 4304 se
rect 6824 4275 7014 4304
tri 7014 4275 7043 4304 sw
tri 7651 4275 7680 4304 se
rect 7680 4275 7870 4304
tri 7870 4275 7899 4304 sw
tri 8507 4275 8536 4304 se
rect 8536 4275 8726 4304
tri 8726 4275 8755 4304 sw
tri 9363 4275 9392 4304 se
rect 9392 4275 9582 4304
tri 9582 4275 9611 4304 sw
tri 10219 4275 10248 4304 se
rect 10248 4275 10438 4304
tri 10438 4275 10467 4304 sw
tri 5934 4270 5939 4275 se
rect 5939 4270 6187 4275
tri 6187 4270 6192 4275 sw
tri 6790 4270 6795 4275 se
rect 6795 4270 7043 4275
tri 7043 4270 7048 4275 sw
tri 7646 4270 7651 4275 se
rect 7651 4270 7899 4275
tri 7899 4270 7904 4275 sw
tri 8502 4270 8507 4275 se
rect 8507 4270 8755 4275
tri 8755 4270 8760 4275 sw
tri 9358 4270 9363 4275 se
rect 9363 4270 9611 4275
tri 9611 4270 9616 4275 sw
tri 10214 4270 10219 4275 se
rect 10219 4270 10467 4275
tri 10467 4270 10472 4275 sw
rect 10860 4270 10918 4308
rect 348 4219 360 4253
rect 394 4219 406 4253
tri 5909 4245 5934 4270 se
rect 5934 4245 6192 4270
tri 6192 4245 6217 4270 sw
tri 6765 4245 6790 4270 se
rect 6790 4245 7048 4270
tri 7048 4245 7073 4270 sw
tri 7621 4245 7646 4270 se
rect 7646 4245 7904 4270
tri 7904 4245 7929 4270 sw
tri 8477 4245 8502 4270 se
rect 8502 4245 8760 4270
tri 8760 4245 8785 4270 sw
tri 9333 4245 9358 4270 se
rect 9358 4245 9616 4270
tri 9616 4245 9641 4270 sw
tri 10189 4245 10214 4270 se
rect 10214 4245 10472 4270
tri 10472 4245 10497 4270 sw
rect 348 4199 406 4219
rect 540 4239 1310 4245
rect 540 4205 552 4239
rect 586 4205 632 4239
rect 666 4205 711 4239
rect 745 4205 790 4239
rect 824 4205 869 4239
rect 903 4205 948 4239
rect 982 4205 1027 4239
rect 1061 4205 1106 4239
rect 1140 4205 1185 4239
rect 1219 4205 1264 4239
rect 1298 4205 1310 4239
tri 406 4199 408 4201 sw
rect 540 4199 1310 4205
rect 1396 4239 2166 4245
rect 1396 4205 1408 4239
rect 1442 4205 1488 4239
rect 1522 4205 1567 4239
rect 1601 4205 1646 4239
rect 1680 4205 1725 4239
rect 1759 4205 1804 4239
rect 1838 4205 1883 4239
rect 1917 4205 1962 4239
rect 1996 4205 2041 4239
rect 2075 4205 2120 4239
rect 2154 4205 2166 4239
rect 1396 4199 2166 4205
rect 2252 4239 3022 4245
rect 2252 4205 2264 4239
rect 2298 4205 2344 4239
rect 2378 4205 2423 4239
rect 2457 4205 2502 4239
rect 2536 4205 2581 4239
rect 2615 4205 2660 4239
rect 2694 4205 2739 4239
rect 2773 4205 2818 4239
rect 2852 4205 2897 4239
rect 2931 4205 2976 4239
rect 3010 4205 3022 4239
rect 2252 4199 3022 4205
rect 3108 4239 3878 4245
rect 3108 4205 3120 4239
rect 3154 4205 3200 4239
rect 3234 4205 3279 4239
rect 3313 4205 3358 4239
rect 3392 4205 3437 4239
rect 3471 4205 3516 4239
rect 3550 4205 3595 4239
rect 3629 4205 3674 4239
rect 3708 4205 3753 4239
rect 3787 4205 3832 4239
rect 3866 4205 3878 4239
rect 3108 4199 3878 4205
rect 3964 4239 4734 4245
rect 3964 4205 3976 4239
rect 4010 4205 4056 4239
rect 4090 4205 4135 4239
rect 4169 4205 4214 4239
rect 4248 4205 4293 4239
rect 4327 4205 4372 4239
rect 4406 4205 4451 4239
rect 4485 4205 4530 4239
rect 4564 4205 4609 4239
rect 4643 4205 4688 4239
rect 4722 4205 4734 4239
rect 3964 4199 4734 4205
rect 4820 4239 5590 4245
rect 4820 4205 4832 4239
rect 4866 4205 4912 4239
rect 4946 4205 4991 4239
rect 5025 4205 5070 4239
rect 5104 4205 5149 4239
rect 5183 4205 5228 4239
rect 5262 4205 5307 4239
rect 5341 4205 5386 4239
rect 5420 4205 5465 4239
rect 5499 4205 5544 4239
rect 5578 4205 5590 4239
rect 4820 4199 5590 4205
rect 5676 4239 6446 4245
rect 5676 4205 5688 4239
rect 5722 4205 5768 4239
rect 5802 4205 5847 4239
rect 5881 4205 5926 4239
rect 5960 4205 6005 4239
rect 6039 4205 6084 4239
rect 6118 4205 6163 4239
rect 6197 4205 6242 4239
rect 6276 4205 6321 4239
rect 6355 4205 6400 4239
rect 6434 4205 6446 4239
rect 5676 4199 6446 4205
rect 6532 4239 7302 4245
rect 6532 4205 6544 4239
rect 6578 4205 6624 4239
rect 6658 4205 6703 4239
rect 6737 4205 6782 4239
rect 6816 4205 6861 4239
rect 6895 4205 6940 4239
rect 6974 4205 7019 4239
rect 7053 4205 7098 4239
rect 7132 4205 7177 4239
rect 7211 4205 7256 4239
rect 7290 4205 7302 4239
rect 6532 4199 7302 4205
rect 7388 4239 8158 4245
rect 7388 4205 7400 4239
rect 7434 4205 7480 4239
rect 7514 4205 7559 4239
rect 7593 4205 7638 4239
rect 7672 4205 7717 4239
rect 7751 4205 7796 4239
rect 7830 4205 7875 4239
rect 7909 4205 7954 4239
rect 7988 4205 8033 4239
rect 8067 4205 8112 4239
rect 8146 4205 8158 4239
rect 7388 4199 8158 4205
rect 8244 4239 9014 4245
rect 8244 4205 8256 4239
rect 8290 4205 8336 4239
rect 8370 4205 8415 4239
rect 8449 4205 8494 4239
rect 8528 4205 8573 4239
rect 8607 4205 8652 4239
rect 8686 4205 8731 4239
rect 8765 4205 8810 4239
rect 8844 4205 8889 4239
rect 8923 4205 8968 4239
rect 9002 4205 9014 4239
rect 8244 4199 9014 4205
rect 9100 4239 9870 4245
rect 9100 4205 9112 4239
rect 9146 4205 9192 4239
rect 9226 4205 9271 4239
rect 9305 4205 9350 4239
rect 9384 4205 9429 4239
rect 9463 4205 9508 4239
rect 9542 4205 9587 4239
rect 9621 4205 9666 4239
rect 9700 4205 9745 4239
rect 9779 4205 9824 4239
rect 9858 4205 9870 4239
rect 9100 4199 9870 4205
rect 9956 4239 10726 4245
rect 9956 4205 9968 4239
rect 10002 4205 10048 4239
rect 10082 4205 10127 4239
rect 10161 4205 10206 4239
rect 10240 4205 10285 4239
rect 10319 4205 10364 4239
rect 10398 4205 10443 4239
rect 10477 4205 10522 4239
rect 10556 4205 10601 4239
rect 10635 4205 10680 4239
rect 10714 4205 10726 4239
rect 9956 4199 10726 4205
rect 10860 4236 10872 4270
rect 10906 4236 10918 4270
rect 348 4174 408 4199
tri 408 4174 433 4199 sw
rect 348 4168 433 4174
tri 433 4168 439 4174 sw
tri 10854 4168 10860 4174 se
rect 10860 4168 10918 4236
rect 348 4160 439 4168
tri 439 4160 447 4168 sw
tri 10846 4160 10854 4168 se
rect 10854 4160 10918 4168
rect 348 4149 447 4160
tri 447 4149 458 4160 sw
tri 10835 4149 10846 4160 se
rect 10846 4149 10918 4160
rect 348 4139 10918 4149
rect 348 4105 379 4139
rect 413 4105 452 4139
rect 486 4105 525 4139
rect 559 4105 598 4139
rect 632 4105 671 4139
rect 705 4105 744 4139
rect 778 4105 817 4139
rect 851 4105 890 4139
rect 924 4105 963 4139
rect 997 4105 1036 4139
rect 1070 4105 1109 4139
rect 1143 4105 1182 4139
rect 1216 4105 1255 4139
rect 1289 4105 1328 4139
rect 1362 4105 1401 4139
rect 1435 4105 1474 4139
rect 1508 4105 1547 4139
rect 1581 4105 1620 4139
rect 1654 4105 1693 4139
rect 1727 4105 1766 4139
rect 1800 4105 1839 4139
rect 1873 4105 1912 4139
rect 1946 4105 1985 4139
rect 2019 4105 2058 4139
rect 2092 4105 2131 4139
rect 2165 4105 2204 4139
rect 2238 4105 2277 4139
rect 2311 4105 2350 4139
rect 2384 4105 2423 4139
rect 2457 4105 2496 4139
rect 2530 4105 2569 4139
rect 2603 4105 2642 4139
rect 2676 4105 2715 4139
rect 2749 4105 2788 4139
rect 2822 4105 2861 4139
rect 2895 4105 2934 4139
rect 2968 4105 3007 4139
rect 3041 4105 3080 4139
rect 3114 4105 3153 4139
rect 3187 4105 3226 4139
rect 3260 4105 3299 4139
rect 3333 4105 3372 4139
rect 3406 4105 3444 4139
rect 3478 4105 3516 4139
rect 3550 4105 3588 4139
rect 3622 4105 3660 4139
rect 3694 4105 3732 4139
rect 3766 4105 3804 4139
rect 3838 4105 3876 4139
rect 3910 4105 3948 4139
rect 3982 4105 4020 4139
rect 4054 4105 4092 4139
rect 4126 4105 4164 4139
rect 4198 4105 4236 4139
rect 4270 4105 4308 4139
rect 4342 4105 4380 4139
rect 4414 4105 4452 4139
rect 4486 4105 4524 4139
rect 4558 4105 4596 4139
rect 4630 4105 4668 4139
rect 4702 4105 4740 4139
rect 4774 4105 4812 4139
rect 4846 4105 4884 4139
rect 4918 4105 4956 4139
rect 4990 4105 5028 4139
rect 5062 4105 5100 4139
rect 5134 4105 5172 4139
rect 5206 4105 5244 4139
rect 5278 4105 5316 4139
rect 5350 4105 5388 4139
rect 5422 4105 5460 4139
rect 5494 4105 5532 4139
rect 5566 4105 5604 4139
rect 5638 4105 5676 4139
rect 5710 4105 5748 4139
rect 5782 4105 5820 4139
rect 5854 4105 5892 4139
rect 5926 4105 5964 4139
rect 5998 4105 6036 4139
rect 6070 4105 6108 4139
rect 6142 4105 6180 4139
rect 6214 4105 6252 4139
rect 6286 4105 6324 4139
rect 6358 4105 6396 4139
rect 6430 4105 6468 4139
rect 6502 4105 6540 4139
rect 6574 4105 6612 4139
rect 6646 4105 6684 4139
rect 6718 4105 6756 4139
rect 6790 4105 6828 4139
rect 6862 4105 6900 4139
rect 6934 4105 6972 4139
rect 7006 4105 7044 4139
rect 7078 4105 7116 4139
rect 7150 4105 7188 4139
rect 7222 4105 7260 4139
rect 7294 4105 7332 4139
rect 7366 4105 7404 4139
rect 7438 4105 7476 4139
rect 7510 4105 7548 4139
rect 7582 4105 7620 4139
rect 7654 4105 7692 4139
rect 7726 4105 7764 4139
rect 7798 4105 7836 4139
rect 7870 4105 7908 4139
rect 7942 4105 7980 4139
rect 8014 4105 8052 4139
rect 8086 4105 8124 4139
rect 8158 4105 8196 4139
rect 8230 4105 8268 4139
rect 8302 4105 8340 4139
rect 8374 4105 8412 4139
rect 8446 4105 8484 4139
rect 8518 4105 8556 4139
rect 8590 4105 8628 4139
rect 8662 4105 8700 4139
rect 8734 4105 8772 4139
rect 8806 4105 8844 4139
rect 8878 4105 8916 4139
rect 8950 4105 8988 4139
rect 9022 4105 9060 4139
rect 9094 4105 9132 4139
rect 9166 4105 9204 4139
rect 9238 4105 9276 4139
rect 9310 4105 9348 4139
rect 9382 4105 9420 4139
rect 9454 4105 9492 4139
rect 9526 4105 9564 4139
rect 9598 4105 9636 4139
rect 9670 4105 9708 4139
rect 9742 4105 9780 4139
rect 9814 4105 9852 4139
rect 9886 4105 9924 4139
rect 9958 4105 9996 4139
rect 10030 4105 10068 4139
rect 10102 4105 10140 4139
rect 10174 4105 10212 4139
rect 10246 4105 10284 4139
rect 10318 4105 10356 4139
rect 10390 4105 10428 4139
rect 10462 4105 10500 4139
rect 10534 4105 10572 4139
rect 10606 4105 10644 4139
rect 10678 4105 10716 4139
rect 10750 4105 10788 4139
rect 10822 4105 10860 4139
rect 10894 4105 10918 4139
rect 348 4097 10918 4105
rect 348 3907 10958 3915
rect 348 3873 379 3907
rect 413 3873 452 3907
rect 486 3873 525 3907
rect 559 3873 598 3907
rect 632 3873 671 3907
rect 705 3873 744 3907
rect 778 3873 817 3907
rect 851 3873 890 3907
rect 924 3873 963 3907
rect 997 3873 1036 3907
rect 1070 3873 1109 3907
rect 1143 3873 1182 3907
rect 1216 3873 1255 3907
rect 1289 3873 1328 3907
rect 1362 3873 1401 3907
rect 1435 3873 1474 3907
rect 1508 3873 1547 3907
rect 1581 3873 1620 3907
rect 1654 3873 1693 3907
rect 1727 3873 1766 3907
rect 1800 3873 1839 3907
rect 1873 3873 1912 3907
rect 1946 3873 1985 3907
rect 2019 3873 2058 3907
rect 2092 3873 2131 3907
rect 2165 3873 2204 3907
rect 2238 3873 2277 3907
rect 2311 3873 2350 3907
rect 2384 3873 2423 3907
rect 2457 3873 2496 3907
rect 2530 3873 2569 3907
rect 2603 3873 2642 3907
rect 2676 3873 2715 3907
rect 2749 3873 2788 3907
rect 2822 3873 2861 3907
rect 2895 3873 2934 3907
rect 2968 3873 3007 3907
rect 3041 3873 3080 3907
rect 3114 3873 3153 3907
rect 3187 3873 3226 3907
rect 3260 3873 3299 3907
rect 3333 3873 3372 3907
rect 3406 3873 3444 3907
rect 3478 3873 3516 3907
rect 3550 3873 3588 3907
rect 3622 3873 3660 3907
rect 3694 3873 3732 3907
rect 3766 3873 3804 3907
rect 3838 3873 3876 3907
rect 3910 3873 3948 3907
rect 3982 3873 4020 3907
rect 4054 3873 4092 3907
rect 4126 3873 4164 3907
rect 4198 3873 4236 3907
rect 4270 3873 4308 3907
rect 4342 3873 4380 3907
rect 4414 3873 4452 3907
rect 4486 3873 4524 3907
rect 4558 3873 4596 3907
rect 4630 3873 4668 3907
rect 4702 3873 4740 3907
rect 4774 3873 4812 3907
rect 4846 3873 4884 3907
rect 4918 3873 4956 3907
rect 4990 3873 5028 3907
rect 5062 3873 5100 3907
rect 5134 3873 5172 3907
rect 5206 3873 5244 3907
rect 5278 3873 5316 3907
rect 5350 3873 5388 3907
rect 5422 3873 5460 3907
rect 5494 3873 5532 3907
rect 5566 3873 5604 3907
rect 5638 3873 5676 3907
rect 5710 3873 5748 3907
rect 5782 3873 5820 3907
rect 5854 3873 5892 3907
rect 5926 3873 5964 3907
rect 5998 3873 6036 3907
rect 6070 3873 6108 3907
rect 6142 3873 6180 3907
rect 6214 3873 6252 3907
rect 6286 3873 6324 3907
rect 6358 3873 6396 3907
rect 6430 3873 6468 3907
rect 6502 3873 6540 3907
rect 6574 3873 6612 3907
rect 6646 3873 6684 3907
rect 6718 3873 6756 3907
rect 6790 3873 6828 3907
rect 6862 3873 6900 3907
rect 6934 3873 6972 3907
rect 7006 3873 7044 3907
rect 7078 3873 7116 3907
rect 7150 3873 7188 3907
rect 7222 3873 7260 3907
rect 7294 3873 7332 3907
rect 7366 3873 7404 3907
rect 7438 3873 7476 3907
rect 7510 3873 7548 3907
rect 7582 3873 7620 3907
rect 7654 3873 7692 3907
rect 7726 3873 7764 3907
rect 7798 3873 7836 3907
rect 7870 3873 7908 3907
rect 7942 3873 7980 3907
rect 8014 3873 8052 3907
rect 8086 3873 8124 3907
rect 8158 3873 8196 3907
rect 8230 3873 8268 3907
rect 8302 3873 8340 3907
rect 8374 3873 8412 3907
rect 8446 3873 8484 3907
rect 8518 3873 8556 3907
rect 8590 3873 8628 3907
rect 8662 3873 8700 3907
rect 8734 3873 8772 3907
rect 8806 3873 8844 3907
rect 8878 3873 8916 3907
rect 8950 3873 8988 3907
rect 9022 3873 9060 3907
rect 9094 3873 9132 3907
rect 9166 3873 9204 3907
rect 9238 3873 9276 3907
rect 9310 3873 9348 3907
rect 9382 3873 9420 3907
rect 9454 3873 9492 3907
rect 9526 3873 9564 3907
rect 9598 3873 9636 3907
rect 9670 3873 9708 3907
rect 9742 3873 9780 3907
rect 9814 3873 9852 3907
rect 9886 3873 9924 3907
rect 9958 3873 9996 3907
rect 10030 3873 10068 3907
rect 10102 3873 10140 3907
rect 10174 3873 10212 3907
rect 10246 3873 10284 3907
rect 10318 3873 10356 3907
rect 10390 3873 10428 3907
rect 10462 3873 10500 3907
rect 10534 3873 10572 3907
rect 10606 3873 10644 3907
rect 10678 3873 10716 3907
rect 10750 3873 10788 3907
rect 10822 3873 10860 3907
rect 10894 3873 10958 3907
rect 348 3863 10958 3873
rect 348 3844 439 3863
tri 439 3844 458 3863 nw
tri 10848 3844 10867 3863 ne
rect 10867 3844 10958 3863
rect 348 3825 420 3844
tri 420 3825 439 3844 nw
tri 10867 3825 10886 3844 ne
rect 10886 3825 10958 3844
rect 348 3790 406 3825
tri 406 3811 420 3825 nw
tri 10886 3811 10900 3825 ne
rect 348 3756 360 3790
rect 394 3756 406 3790
rect 540 3803 1310 3809
rect 540 3769 552 3803
rect 586 3769 632 3803
rect 666 3769 711 3803
rect 745 3769 790 3803
rect 824 3769 869 3803
rect 903 3769 948 3803
rect 982 3769 1027 3803
rect 1061 3769 1106 3803
rect 1140 3769 1185 3803
rect 1219 3769 1264 3803
rect 1298 3769 1310 3803
rect 540 3763 1310 3769
rect 1396 3803 2166 3809
rect 1396 3769 1408 3803
rect 1442 3769 1488 3803
rect 1522 3769 1567 3803
rect 1601 3769 1646 3803
rect 1680 3769 1725 3803
rect 1759 3769 1804 3803
rect 1838 3769 1883 3803
rect 1917 3769 1962 3803
rect 1996 3769 2041 3803
rect 2075 3769 2120 3803
rect 2154 3769 2166 3803
rect 1396 3763 2166 3769
rect 2252 3803 3022 3809
rect 2252 3769 2264 3803
rect 2298 3769 2344 3803
rect 2378 3769 2423 3803
rect 2457 3769 2502 3803
rect 2536 3769 2581 3803
rect 2615 3769 2660 3803
rect 2694 3769 2739 3803
rect 2773 3769 2818 3803
rect 2852 3769 2897 3803
rect 2931 3769 2976 3803
rect 3010 3769 3022 3803
rect 2252 3763 3022 3769
rect 3108 3803 3878 3809
rect 3108 3769 3120 3803
rect 3154 3769 3200 3803
rect 3234 3769 3279 3803
rect 3313 3769 3358 3803
rect 3392 3769 3437 3803
rect 3471 3769 3516 3803
rect 3550 3769 3595 3803
rect 3629 3769 3674 3803
rect 3708 3769 3753 3803
rect 3787 3769 3832 3803
rect 3866 3769 3878 3803
rect 3108 3763 3878 3769
rect 3964 3803 4734 3809
rect 3964 3769 3976 3803
rect 4010 3769 4056 3803
rect 4090 3769 4135 3803
rect 4169 3769 4214 3803
rect 4248 3769 4293 3803
rect 4327 3769 4372 3803
rect 4406 3769 4451 3803
rect 4485 3769 4530 3803
rect 4564 3769 4609 3803
rect 4643 3769 4688 3803
rect 4722 3769 4734 3803
rect 3964 3763 4734 3769
rect 4820 3803 5590 3809
rect 4820 3769 4832 3803
rect 4866 3769 4912 3803
rect 4946 3769 4991 3803
rect 5025 3769 5070 3803
rect 5104 3769 5149 3803
rect 5183 3769 5228 3803
rect 5262 3769 5307 3803
rect 5341 3769 5386 3803
rect 5420 3769 5465 3803
rect 5499 3769 5544 3803
rect 5578 3769 5590 3803
rect 4820 3763 5590 3769
rect 5676 3803 6446 3809
rect 5676 3769 5688 3803
rect 5722 3769 5768 3803
rect 5802 3769 5847 3803
rect 5881 3769 5926 3803
rect 5960 3769 6005 3803
rect 6039 3769 6084 3803
rect 6118 3769 6163 3803
rect 6197 3769 6242 3803
rect 6276 3769 6321 3803
rect 6355 3769 6400 3803
rect 6434 3769 6446 3803
rect 5676 3763 6446 3769
rect 6532 3803 7302 3809
rect 6532 3769 6544 3803
rect 6578 3769 6624 3803
rect 6658 3769 6703 3803
rect 6737 3769 6782 3803
rect 6816 3769 6861 3803
rect 6895 3769 6940 3803
rect 6974 3769 7019 3803
rect 7053 3769 7098 3803
rect 7132 3769 7177 3803
rect 7211 3769 7256 3803
rect 7290 3769 7302 3803
rect 6532 3763 7302 3769
rect 7388 3803 8158 3809
rect 7388 3769 7400 3803
rect 7434 3769 7480 3803
rect 7514 3769 7559 3803
rect 7593 3769 7638 3803
rect 7672 3769 7717 3803
rect 7751 3769 7796 3803
rect 7830 3769 7875 3803
rect 7909 3769 7954 3803
rect 7988 3769 8033 3803
rect 8067 3769 8112 3803
rect 8146 3769 8158 3803
rect 7388 3763 8158 3769
rect 8244 3803 9014 3809
rect 8244 3769 8256 3803
rect 8290 3769 8336 3803
rect 8370 3769 8415 3803
rect 8449 3769 8494 3803
rect 8528 3769 8573 3803
rect 8607 3769 8652 3803
rect 8686 3769 8731 3803
rect 8765 3769 8810 3803
rect 8844 3769 8889 3803
rect 8923 3769 8968 3803
rect 9002 3769 9014 3803
rect 8244 3763 9014 3769
rect 9100 3803 9870 3809
rect 9100 3769 9112 3803
rect 9146 3769 9192 3803
rect 9226 3769 9271 3803
rect 9305 3769 9350 3803
rect 9384 3769 9429 3803
rect 9463 3769 9508 3803
rect 9542 3769 9587 3803
rect 9621 3769 9666 3803
rect 9700 3769 9745 3803
rect 9779 3769 9824 3803
rect 9858 3769 9870 3803
rect 9100 3763 9870 3769
rect 9956 3803 10726 3809
rect 9956 3769 9968 3803
rect 10002 3769 10048 3803
rect 10082 3769 10127 3803
rect 10161 3769 10206 3803
rect 10240 3769 10285 3803
rect 10319 3769 10364 3803
rect 10398 3769 10443 3803
rect 10477 3769 10522 3803
rect 10556 3769 10601 3803
rect 10635 3769 10680 3803
rect 10714 3769 10726 3803
rect 9956 3763 10726 3769
rect 10900 3790 10958 3825
tri 773 3756 780 3763 ne
rect 780 3756 1074 3763
tri 1074 3756 1081 3763 nw
tri 1629 3756 1636 3763 ne
rect 1636 3756 1930 3763
tri 1930 3756 1937 3763 nw
tri 2485 3756 2492 3763 ne
rect 2492 3756 2786 3763
tri 2786 3756 2793 3763 nw
tri 3341 3756 3348 3763 ne
rect 3348 3756 3642 3763
tri 3642 3756 3649 3763 nw
tri 4197 3756 4204 3763 ne
rect 4204 3756 4498 3763
tri 4498 3756 4505 3763 nw
tri 5053 3756 5060 3763 ne
rect 5060 3756 5354 3763
tri 5354 3756 5361 3763 nw
rect 5998 3759 6128 3763
tri 5860 3756 5863 3759 ne
rect 5863 3756 6263 3759
tri 6263 3756 6266 3759 nw
rect 10900 3756 10912 3790
rect 10946 3756 10958 3790
rect 348 3718 406 3756
tri 780 3754 782 3756 ne
rect 782 3754 1072 3756
tri 1072 3754 1074 3756 nw
tri 1636 3754 1638 3756 ne
rect 1638 3754 1928 3756
tri 1928 3754 1930 3756 nw
tri 2492 3754 2494 3756 ne
rect 2494 3754 2784 3756
tri 2784 3754 2786 3756 nw
tri 3348 3754 3350 3756 ne
rect 3350 3754 3640 3756
tri 3640 3754 3642 3756 nw
tri 4204 3754 4206 3756 ne
rect 4206 3754 4496 3756
tri 4496 3754 4498 3756 nw
tri 5060 3754 5062 3756 ne
rect 5062 3754 5352 3756
tri 5352 3754 5354 3756 nw
tri 5863 3754 5865 3756 ne
rect 5865 3754 6261 3756
tri 6261 3754 6263 3756 nw
tri 782 3734 802 3754 ne
rect 802 3734 1052 3754
tri 1052 3734 1072 3754 nw
tri 1638 3734 1658 3754 ne
rect 1658 3734 1908 3754
tri 1908 3734 1928 3754 nw
tri 2494 3734 2514 3754 ne
rect 2514 3734 2764 3754
tri 2764 3734 2784 3754 nw
tri 3350 3734 3370 3754 ne
rect 3370 3734 3620 3754
tri 3620 3734 3640 3754 nw
tri 4206 3734 4226 3754 ne
rect 4226 3734 4476 3754
tri 4476 3734 4496 3754 nw
tri 5062 3734 5082 3754 ne
rect 5082 3734 5332 3754
tri 5332 3734 5352 3754 nw
tri 5865 3734 5885 3754 ne
rect 5885 3734 6241 3754
tri 6241 3734 6261 3754 nw
tri 802 3718 818 3734 ne
rect 818 3718 1036 3734
tri 1036 3718 1052 3734 nw
tri 1658 3718 1674 3734 ne
rect 1674 3718 1892 3734
tri 1892 3718 1908 3734 nw
tri 2514 3718 2530 3734 ne
rect 2530 3718 2748 3734
tri 2748 3718 2764 3734 nw
tri 3370 3718 3386 3734 ne
rect 3386 3718 3604 3734
tri 3604 3718 3620 3734 nw
tri 4226 3718 4242 3734 ne
rect 4242 3718 4460 3734
tri 4460 3718 4476 3734 nw
tri 5082 3718 5098 3734 ne
rect 5098 3718 5316 3734
tri 5316 3718 5332 3734 nw
tri 5885 3718 5901 3734 ne
rect 5901 3718 6225 3734
tri 6225 3718 6241 3734 nw
rect 10900 3718 10958 3756
rect 348 3684 360 3718
rect 394 3684 406 3718
tri 818 3684 852 3718 ne
rect 852 3684 1002 3718
tri 1002 3684 1036 3718 nw
tri 1674 3684 1708 3718 ne
rect 1708 3684 1858 3718
tri 1858 3684 1892 3718 nw
tri 2530 3684 2564 3718 ne
rect 2564 3684 2714 3718
tri 2714 3684 2748 3718 nw
tri 3386 3684 3420 3718 ne
rect 3420 3684 3570 3718
tri 3570 3684 3604 3718 nw
tri 4242 3684 4276 3718 ne
rect 4276 3684 4426 3718
tri 4426 3684 4460 3718 nw
tri 5098 3684 5132 3718 ne
rect 5132 3684 5282 3718
tri 5282 3684 5316 3718 nw
tri 5901 3684 5935 3718 ne
rect 5935 3684 6191 3718
tri 6191 3684 6225 3718 nw
rect 10900 3684 10912 3718
rect 10946 3684 10958 3718
rect 348 3646 406 3684
tri 852 3674 862 3684 ne
rect 348 3612 360 3646
rect 394 3612 406 3646
rect 348 3574 406 3612
rect 348 3540 360 3574
rect 394 3540 406 3574
rect 348 3502 406 3540
rect 348 3468 360 3502
rect 394 3468 406 3502
rect 348 3430 406 3468
rect 348 3396 360 3430
rect 394 3396 406 3430
rect 348 3358 406 3396
rect 348 3324 360 3358
rect 394 3324 406 3358
rect 348 3286 406 3324
rect 348 3252 360 3286
rect 394 3252 406 3286
rect 348 3214 406 3252
rect 348 3180 360 3214
rect 394 3180 406 3214
rect 348 3142 406 3180
rect 348 3108 360 3142
rect 394 3108 406 3142
rect 348 3070 406 3108
rect 348 3036 360 3070
rect 394 3036 406 3070
rect 348 2998 406 3036
rect 348 2964 360 2998
rect 394 2964 406 2998
rect 348 2926 406 2964
rect 348 2892 360 2926
rect 394 2892 406 2926
rect 348 2854 406 2892
rect 348 2820 360 2854
rect 394 2820 406 2854
rect 348 2782 406 2820
rect 348 2748 360 2782
rect 394 2748 406 2782
rect 348 2710 406 2748
rect 488 3646 546 3652
rect 488 3637 500 3646
rect 534 3637 546 3646
rect 488 3585 491 3637
rect 543 3585 546 3637
rect 488 3574 546 3585
rect 488 3573 500 3574
rect 534 3573 546 3574
rect 488 3521 491 3573
rect 543 3521 546 3573
rect 488 3509 546 3521
rect 488 3457 491 3509
rect 543 3457 546 3509
rect 488 3445 546 3457
rect 488 3393 491 3445
rect 543 3393 546 3445
rect 488 3381 546 3393
rect 488 3329 491 3381
rect 543 3329 546 3381
rect 488 3324 500 3329
rect 534 3324 546 3329
rect 488 3317 546 3324
rect 488 3265 491 3317
rect 543 3265 546 3317
rect 488 3253 500 3265
rect 534 3253 546 3265
rect 488 3201 491 3253
rect 543 3201 546 3253
rect 488 3189 500 3201
rect 534 3189 546 3201
rect 488 3137 491 3189
rect 543 3137 546 3189
rect 488 3125 500 3137
rect 534 3125 546 3137
rect 488 3073 491 3125
rect 543 3073 546 3125
rect 488 3070 546 3073
rect 488 3061 500 3070
rect 534 3061 546 3070
rect 488 3009 491 3061
rect 543 3009 546 3061
rect 488 2998 546 3009
rect 488 2997 500 2998
rect 534 2997 546 2998
rect 488 2945 491 2997
rect 543 2945 546 2997
rect 488 2933 546 2945
rect 488 2881 491 2933
rect 543 2881 546 2933
rect 488 2869 546 2881
rect 488 2817 491 2869
rect 543 2817 546 2869
rect 488 2805 546 2817
rect 488 2753 491 2805
rect 543 2753 546 2805
rect 488 2748 500 2753
rect 534 2748 546 2753
rect 488 2742 546 2748
rect 348 2685 360 2710
rect 394 2685 406 2710
rect 348 2633 351 2685
rect 403 2633 406 2685
rect 348 2621 360 2633
rect 394 2621 406 2633
rect 348 2569 351 2621
rect 403 2569 406 2621
rect 348 2566 406 2569
rect 348 2557 360 2566
rect 394 2557 406 2566
rect 348 2505 351 2557
rect 403 2505 406 2557
rect 348 2494 406 2505
rect 348 2493 360 2494
rect 394 2493 406 2494
rect 348 2441 351 2493
rect 403 2441 406 2493
rect 348 2429 406 2441
rect 348 2377 351 2429
rect 403 2377 406 2429
rect 348 2365 406 2377
rect 348 2313 351 2365
rect 403 2313 406 2365
rect 348 2301 406 2313
rect 348 2249 351 2301
rect 403 2260 406 2301
tri 406 2260 430 2284 sw
rect 403 2249 430 2260
rect 348 2244 360 2249
rect 394 2244 430 2249
rect 348 2243 430 2244
tri 430 2243 447 2260 sw
rect 348 2232 447 2243
tri 447 2232 458 2243 sw
rect 348 2180 381 2232
rect 433 2180 445 2232
rect 497 2180 509 2232
rect 561 2223 573 2232
rect 625 2223 637 2232
rect 562 2189 573 2223
rect 634 2189 637 2223
rect 561 2180 573 2189
rect 625 2180 637 2189
rect 689 2180 695 2232
rect 348 2102 354 2154
rect 406 2102 418 2154
rect 470 2102 482 2154
rect 534 2102 546 2154
rect 598 2102 610 2154
rect 662 2102 674 2154
rect 726 2102 732 2154
rect 348 2023 354 2075
rect 406 2023 418 2075
rect 470 2069 482 2075
rect 534 2069 546 2075
rect 598 2069 610 2075
rect 662 2069 674 2075
rect 662 2035 665 2069
rect 470 2023 482 2035
rect 534 2023 546 2035
rect 598 2023 610 2035
rect 662 2023 674 2035
rect 726 2023 732 2075
rect 348 1990 425 2023
tri 425 1990 458 2023 nw
rect 348 1988 406 1990
rect 348 1954 360 1988
rect 394 1954 406 1988
tri 406 1971 425 1990 nw
rect 348 1916 406 1954
rect 348 1882 360 1916
rect 394 1882 406 1916
rect 348 1844 406 1882
rect 466 1881 473 1933
rect 525 1881 537 1933
rect 589 1881 596 1933
rect 348 1810 360 1844
rect 394 1810 406 1844
rect 348 1772 406 1810
rect 862 1779 992 3684
tri 992 3674 1002 3684 nw
tri 1708 3674 1718 3684 ne
rect 1344 3664 1402 3670
rect 1344 3637 1356 3664
rect 1390 3637 1402 3664
rect 1344 3585 1347 3637
rect 1399 3585 1402 3637
rect 1344 3573 1356 3585
rect 1390 3573 1402 3585
rect 1344 3521 1347 3573
rect 1399 3521 1402 3573
rect 1344 3520 1402 3521
rect 1344 3509 1356 3520
rect 1390 3509 1402 3520
rect 1344 3457 1347 3509
rect 1399 3457 1402 3509
rect 1344 3448 1402 3457
rect 1344 3445 1356 3448
rect 1390 3445 1402 3448
rect 1344 3393 1347 3445
rect 1399 3393 1402 3445
rect 1344 3381 1402 3393
rect 1344 3329 1347 3381
rect 1399 3329 1402 3381
rect 1344 3317 1402 3329
rect 1344 3265 1347 3317
rect 1399 3265 1402 3317
rect 1344 3253 1402 3265
rect 1344 3201 1347 3253
rect 1399 3201 1402 3253
rect 1344 3198 1356 3201
rect 1390 3198 1402 3201
rect 1344 3189 1402 3198
rect 1344 3137 1347 3189
rect 1399 3137 1402 3189
rect 1344 3126 1356 3137
rect 1390 3126 1402 3137
rect 1344 3125 1402 3126
rect 1344 3073 1347 3125
rect 1399 3073 1402 3125
rect 1344 3061 1356 3073
rect 1390 3061 1402 3073
rect 1344 3009 1347 3061
rect 1399 3009 1402 3061
rect 1344 2997 1356 3009
rect 1390 2997 1402 3009
rect 1344 2945 1347 2997
rect 1399 2945 1402 2997
rect 1344 2944 1402 2945
rect 1344 2933 1356 2944
rect 1390 2933 1402 2944
rect 1344 2881 1347 2933
rect 1399 2881 1402 2933
rect 1344 2872 1402 2881
rect 1344 2869 1356 2872
rect 1390 2869 1402 2872
rect 1344 2817 1347 2869
rect 1399 2817 1402 2869
rect 1344 2805 1402 2817
rect 1344 2753 1347 2805
rect 1399 2753 1402 2805
rect 1344 2728 1402 2753
rect 1344 2694 1356 2728
rect 1390 2694 1402 2728
rect 1344 2656 1402 2694
rect 1344 2622 1356 2656
rect 1390 2622 1402 2656
rect 1344 2584 1402 2622
rect 1344 2550 1356 2584
rect 1390 2550 1402 2584
rect 1344 2512 1402 2550
rect 1344 2478 1356 2512
rect 1390 2478 1402 2512
rect 1344 2440 1402 2478
rect 1344 2406 1356 2440
rect 1390 2406 1402 2440
rect 1344 2368 1402 2406
rect 1344 2334 1356 2368
rect 1390 2334 1402 2368
rect 1041 2177 1047 2229
rect 1099 2223 1111 2229
rect 1163 2223 1175 2229
rect 1227 2223 1239 2229
rect 1103 2189 1111 2223
rect 1099 2177 1111 2189
rect 1163 2177 1175 2189
rect 1227 2177 1239 2189
rect 1291 2177 1297 2229
rect 1041 2102 1047 2154
rect 1099 2102 1111 2154
rect 1163 2102 1175 2154
rect 1227 2102 1239 2154
rect 1291 2102 1297 2154
rect 1041 2023 1047 2075
rect 1099 2069 1111 2075
rect 1163 2069 1175 2075
rect 1227 2069 1239 2075
rect 1103 2035 1111 2069
rect 1099 2023 1111 2035
rect 1163 2023 1175 2035
rect 1227 2023 1239 2035
rect 1291 2023 1297 2075
rect 1344 1991 1402 2334
rect 1430 2177 1436 2229
rect 1488 2223 1500 2229
rect 1552 2223 1564 2229
rect 1616 2223 1628 2229
rect 1492 2189 1500 2223
rect 1488 2177 1500 2189
rect 1552 2177 1564 2189
rect 1616 2177 1628 2189
rect 1680 2177 1686 2229
rect 1430 2102 1436 2154
rect 1488 2102 1500 2154
rect 1552 2102 1564 2154
rect 1616 2102 1628 2154
rect 1680 2102 1686 2154
rect 1430 2023 1436 2075
rect 1488 2069 1500 2075
rect 1552 2069 1564 2075
rect 1616 2069 1628 2075
rect 1492 2035 1500 2069
rect 1488 2023 1500 2035
rect 1552 2023 1564 2035
rect 1616 2023 1628 2035
rect 1680 2023 1686 2075
rect 1345 1989 1401 1990
rect 1345 1960 1401 1961
tri 1336 1951 1344 1959 se
rect 1344 1951 1402 1959
tri 1402 1951 1410 1959 sw
tri 1318 1933 1336 1951 se
rect 1336 1933 1410 1951
tri 1410 1933 1428 1951 sw
rect 1309 1881 1315 1933
rect 1367 1881 1379 1933
rect 1431 1881 1437 1933
rect 348 1738 360 1772
rect 394 1738 406 1772
rect 348 1700 406 1738
rect 348 1666 360 1700
rect 394 1666 406 1700
rect 348 1628 406 1666
rect 348 1594 360 1628
rect 394 1594 406 1628
rect 348 1556 406 1594
rect 466 1727 473 1779
rect 525 1727 537 1779
rect 589 1727 596 1779
rect 862 1727 869 1779
rect 921 1727 933 1779
rect 985 1727 992 1779
rect 466 1691 596 1727
rect 466 1664 467 1690
rect 468 1663 594 1691
rect 595 1664 596 1690
rect 466 1625 596 1663
rect 466 1573 473 1625
rect 525 1573 537 1625
rect 589 1573 596 1625
rect 348 1522 360 1556
rect 394 1522 406 1556
rect 348 1484 406 1522
rect 348 1450 360 1484
rect 394 1450 406 1484
rect 1718 1471 1848 3684
tri 1848 3674 1858 3684 nw
tri 2564 3674 2574 3684 ne
rect 2200 3664 2258 3670
rect 2200 3637 2212 3664
rect 2246 3637 2258 3664
rect 2200 3585 2203 3637
rect 2255 3585 2258 3637
rect 2200 3573 2212 3585
rect 2246 3573 2258 3585
rect 2200 3521 2203 3573
rect 2255 3521 2258 3573
rect 2200 3520 2258 3521
rect 2200 3509 2212 3520
rect 2246 3509 2258 3520
rect 2200 3457 2203 3509
rect 2255 3457 2258 3509
rect 2200 3448 2258 3457
rect 2200 3445 2212 3448
rect 2246 3445 2258 3448
rect 2200 3393 2203 3445
rect 2255 3393 2258 3445
rect 2200 3381 2258 3393
rect 2200 3329 2203 3381
rect 2255 3329 2258 3381
rect 2200 3317 2258 3329
rect 2200 3265 2203 3317
rect 2255 3265 2258 3317
rect 2200 3253 2258 3265
rect 2200 3201 2203 3253
rect 2255 3201 2258 3253
rect 2200 3198 2212 3201
rect 2246 3198 2258 3201
rect 2200 3189 2258 3198
rect 2200 3137 2203 3189
rect 2255 3137 2258 3189
rect 2200 3126 2212 3137
rect 2246 3126 2258 3137
rect 2200 3125 2258 3126
rect 2200 3073 2203 3125
rect 2255 3073 2258 3125
rect 2200 3061 2212 3073
rect 2246 3061 2258 3073
rect 2200 3009 2203 3061
rect 2255 3009 2258 3061
rect 2200 2997 2212 3009
rect 2246 2997 2258 3009
rect 2200 2945 2203 2997
rect 2255 2945 2258 2997
rect 2200 2944 2258 2945
rect 2200 2933 2212 2944
rect 2246 2933 2258 2944
rect 2200 2881 2203 2933
rect 2255 2881 2258 2933
rect 2200 2872 2258 2881
rect 2200 2869 2212 2872
rect 2246 2869 2258 2872
rect 2200 2817 2203 2869
rect 2255 2817 2258 2869
rect 2200 2805 2258 2817
rect 2200 2753 2203 2805
rect 2255 2753 2258 2805
rect 2200 2728 2258 2753
rect 2200 2694 2212 2728
rect 2246 2694 2258 2728
rect 2200 2656 2258 2694
rect 2200 2622 2212 2656
rect 2246 2622 2258 2656
rect 2200 2584 2258 2622
rect 2200 2550 2212 2584
rect 2246 2550 2258 2584
rect 2200 2512 2258 2550
rect 2200 2478 2212 2512
rect 2246 2478 2258 2512
rect 2200 2440 2258 2478
rect 2200 2406 2212 2440
rect 2246 2406 2258 2440
rect 2200 2368 2258 2406
rect 2200 2334 2212 2368
rect 2246 2334 2258 2368
rect 1884 2177 1890 2229
rect 1942 2223 1954 2229
rect 2006 2223 2018 2229
rect 2070 2223 2082 2229
rect 1946 2189 1954 2223
rect 1942 2177 1954 2189
rect 2006 2177 2018 2189
rect 2070 2177 2082 2189
rect 2134 2177 2140 2229
rect 1884 2102 1890 2154
rect 1942 2102 1954 2154
rect 2006 2102 2018 2154
rect 2070 2102 2082 2154
rect 2134 2102 2140 2154
rect 1884 2023 1890 2075
rect 1942 2069 1954 2075
rect 2006 2069 2018 2075
rect 2070 2069 2082 2075
rect 1946 2035 1954 2069
rect 1942 2023 1954 2035
rect 2006 2023 2018 2035
rect 2070 2023 2082 2035
rect 2134 2023 2140 2075
rect 2200 1683 2258 2334
rect 2289 2177 2295 2229
rect 2347 2223 2359 2229
rect 2411 2223 2423 2229
rect 2475 2223 2487 2229
rect 2351 2189 2359 2223
rect 2347 2177 2359 2189
rect 2411 2177 2423 2189
rect 2475 2177 2487 2189
rect 2539 2177 2545 2229
rect 2289 2102 2295 2154
rect 2347 2102 2359 2154
rect 2411 2102 2423 2154
rect 2475 2102 2487 2154
rect 2539 2102 2545 2154
rect 2289 2023 2295 2075
rect 2347 2069 2359 2075
rect 2411 2069 2423 2075
rect 2475 2069 2487 2075
rect 2351 2035 2359 2069
rect 2347 2023 2359 2035
rect 2411 2023 2423 2035
rect 2475 2023 2487 2035
rect 2539 2023 2545 2075
rect 2201 1681 2257 1682
rect 2201 1652 2257 1653
tri 2174 1625 2200 1651 se
rect 2200 1625 2258 1651
tri 2258 1625 2284 1651 sw
rect 2165 1573 2171 1625
rect 2223 1573 2235 1625
rect 2287 1573 2293 1625
rect 348 1412 406 1450
rect 348 1378 360 1412
rect 394 1378 406 1412
rect 466 1419 473 1471
rect 525 1419 537 1471
rect 589 1419 596 1471
rect 1718 1419 1725 1471
rect 1777 1419 1789 1471
rect 1841 1419 1848 1471
rect 466 1386 596 1419
rect 467 1384 595 1385
rect 348 1340 406 1378
rect 348 1306 360 1340
rect 394 1306 406 1340
rect 348 1268 406 1306
rect 348 1234 360 1268
rect 394 1234 406 1268
rect 467 1355 595 1356
rect 466 1317 596 1354
rect 466 1265 473 1317
rect 525 1265 537 1317
rect 589 1265 596 1317
rect 348 1196 406 1234
rect 348 1162 360 1196
rect 394 1162 406 1196
rect 2574 1163 2704 3684
tri 2704 3674 2714 3684 nw
tri 3420 3674 3430 3684 ne
rect 3056 3664 3114 3670
rect 3056 3637 3068 3664
rect 3102 3637 3114 3664
rect 3056 3585 3059 3637
rect 3111 3585 3114 3637
rect 3056 3573 3068 3585
rect 3102 3573 3114 3585
rect 3056 3521 3059 3573
rect 3111 3521 3114 3573
rect 3056 3520 3114 3521
rect 3056 3509 3068 3520
rect 3102 3509 3114 3520
rect 3056 3457 3059 3509
rect 3111 3457 3114 3509
rect 3056 3448 3114 3457
rect 3056 3445 3068 3448
rect 3102 3445 3114 3448
rect 3056 3393 3059 3445
rect 3111 3393 3114 3445
rect 3056 3381 3114 3393
rect 3056 3329 3059 3381
rect 3111 3329 3114 3381
rect 3056 3317 3114 3329
rect 3056 3265 3059 3317
rect 3111 3265 3114 3317
rect 3056 3253 3114 3265
rect 3056 3201 3059 3253
rect 3111 3201 3114 3253
rect 3056 3198 3068 3201
rect 3102 3198 3114 3201
rect 3056 3189 3114 3198
rect 3056 3137 3059 3189
rect 3111 3137 3114 3189
rect 3056 3126 3068 3137
rect 3102 3126 3114 3137
rect 3056 3125 3114 3126
rect 3056 3073 3059 3125
rect 3111 3073 3114 3125
rect 3056 3061 3068 3073
rect 3102 3061 3114 3073
rect 3056 3009 3059 3061
rect 3111 3009 3114 3061
rect 3056 2997 3068 3009
rect 3102 2997 3114 3009
rect 3056 2945 3059 2997
rect 3111 2945 3114 2997
rect 3056 2944 3114 2945
rect 3056 2933 3068 2944
rect 3102 2933 3114 2944
rect 3056 2881 3059 2933
rect 3111 2881 3114 2933
rect 3056 2872 3114 2881
rect 3056 2869 3068 2872
rect 3102 2869 3114 2872
rect 3056 2817 3059 2869
rect 3111 2817 3114 2869
rect 3056 2805 3114 2817
rect 3056 2753 3059 2805
rect 3111 2753 3114 2805
rect 3056 2728 3114 2753
rect 3056 2694 3068 2728
rect 3102 2694 3114 2728
rect 3056 2656 3114 2694
rect 3056 2622 3068 2656
rect 3102 2622 3114 2656
rect 3056 2584 3114 2622
rect 3056 2550 3068 2584
rect 3102 2550 3114 2584
rect 3056 2512 3114 2550
rect 3056 2478 3068 2512
rect 3102 2478 3114 2512
rect 3430 2532 3560 3684
tri 3560 3674 3570 3684 nw
tri 4276 3674 4286 3684 ne
rect 3912 3664 3970 3670
rect 3912 3637 3924 3664
rect 3958 3637 3970 3664
rect 3912 3585 3915 3637
rect 3967 3585 3970 3637
rect 3912 3573 3924 3585
rect 3958 3573 3970 3585
rect 3912 3521 3915 3573
rect 3967 3521 3970 3573
rect 3912 3520 3970 3521
rect 3912 3509 3924 3520
rect 3958 3509 3970 3520
rect 3912 3457 3915 3509
rect 3967 3457 3970 3509
rect 3912 3448 3970 3457
rect 3912 3445 3924 3448
rect 3958 3445 3970 3448
rect 3912 3393 3915 3445
rect 3967 3393 3970 3445
rect 3912 3381 3970 3393
rect 3912 3329 3915 3381
rect 3967 3329 3970 3381
rect 3912 3317 3970 3329
rect 3912 3265 3915 3317
rect 3967 3265 3970 3317
rect 3912 3253 3970 3265
rect 3912 3201 3915 3253
rect 3967 3201 3970 3253
rect 3912 3198 3924 3201
rect 3958 3198 3970 3201
rect 3912 3189 3970 3198
rect 3912 3137 3915 3189
rect 3967 3137 3970 3189
rect 3912 3126 3924 3137
rect 3958 3126 3970 3137
rect 3912 3125 3970 3126
rect 3912 3073 3915 3125
rect 3967 3073 3970 3125
rect 3912 3061 3924 3073
rect 3958 3061 3970 3073
rect 3912 3009 3915 3061
rect 3967 3009 3970 3061
rect 3912 2997 3924 3009
rect 3958 2997 3970 3009
rect 3912 2945 3915 2997
rect 3967 2945 3970 2997
rect 3912 2944 3970 2945
rect 3912 2933 3924 2944
rect 3958 2933 3970 2944
rect 3912 2881 3915 2933
rect 3967 2881 3970 2933
rect 3912 2872 3970 2881
rect 3912 2869 3924 2872
rect 3958 2869 3970 2872
rect 3912 2817 3915 2869
rect 3967 2817 3970 2869
rect 3912 2805 3970 2817
rect 3912 2753 3915 2805
rect 3967 2753 3970 2805
rect 3912 2728 3970 2753
rect 3912 2694 3924 2728
rect 3958 2694 3970 2728
rect 3912 2656 3970 2694
rect 3912 2622 3924 2656
rect 3958 2622 3970 2656
rect 3912 2584 3970 2622
rect 3912 2550 3924 2584
rect 3958 2550 3970 2584
tri 3560 2532 3577 2549 sw
rect 3430 2522 3577 2532
tri 3577 2522 3587 2532 sw
rect 3430 2512 3587 2522
tri 3587 2512 3597 2522 sw
rect 3912 2512 3970 2550
rect 3430 2495 3597 2512
tri 3430 2478 3447 2495 ne
rect 3447 2478 3597 2495
tri 3597 2478 3631 2512 sw
rect 3912 2478 3924 2512
rect 3958 2478 3970 2512
rect 3056 2440 3114 2478
tri 3447 2460 3465 2478 ne
rect 3465 2460 3631 2478
tri 3631 2460 3649 2478 sw
tri 3465 2440 3485 2460 ne
rect 3485 2440 3649 2460
tri 3649 2440 3669 2460 sw
rect 3912 2440 3970 2478
rect 3056 2406 3068 2440
rect 3102 2406 3114 2440
tri 3485 2408 3517 2440 ne
rect 3517 2408 3669 2440
tri 3669 2408 3701 2440 sw
tri 3517 2406 3519 2408 ne
rect 3519 2406 3701 2408
tri 3701 2406 3703 2408 sw
rect 3912 2406 3924 2440
rect 3958 2406 3970 2440
rect 3056 2368 3114 2406
tri 3519 2388 3537 2406 ne
rect 3537 2388 3703 2406
tri 3703 2388 3721 2406 sw
tri 3537 2368 3557 2388 ne
rect 3557 2368 3721 2388
tri 3721 2368 3741 2388 sw
rect 3912 2368 3970 2406
rect 3056 2334 3068 2368
rect 3102 2334 3114 2368
tri 3557 2365 3560 2368 ne
rect 3560 2365 3741 2368
tri 3560 2334 3591 2365 ne
rect 3591 2334 3741 2365
tri 3741 2334 3775 2368 sw
rect 3912 2334 3924 2368
rect 3958 2334 3970 2368
rect 2753 2177 2759 2229
rect 2811 2223 2823 2229
rect 2875 2223 2887 2229
rect 2939 2223 2951 2229
rect 2815 2189 2823 2223
rect 2811 2177 2823 2189
rect 2875 2177 2887 2189
rect 2939 2177 2951 2189
rect 3003 2177 3009 2229
rect 2753 2102 2759 2154
rect 2811 2102 2823 2154
rect 2875 2102 2887 2154
rect 2939 2102 2951 2154
rect 3003 2102 3009 2154
rect 2753 2023 2759 2075
rect 2811 2069 2823 2075
rect 2875 2069 2887 2075
rect 2939 2069 2951 2075
rect 2815 2035 2823 2069
rect 2811 2023 2823 2035
rect 2875 2023 2887 2035
rect 2939 2023 2951 2035
rect 3003 2023 3009 2075
rect 3056 1377 3114 2334
tri 3591 2328 3597 2334 ne
rect 3597 2328 3775 2334
tri 3775 2328 3781 2334 sw
rect 3912 2328 3970 2334
tri 3597 2316 3609 2328 ne
rect 3609 2316 3781 2328
tri 3781 2316 3793 2328 sw
tri 3609 2294 3631 2316 ne
rect 3631 2294 3793 2316
tri 3793 2294 3815 2316 sw
tri 3631 2260 3665 2294 ne
rect 3665 2260 3815 2294
tri 3815 2260 3849 2294 sw
tri 3665 2243 3682 2260 ne
rect 3682 2243 3849 2260
tri 3849 2243 3866 2260 sw
tri 3682 2232 3693 2243 ne
rect 3693 2232 3866 2243
rect 3203 2180 3209 2232
rect 3261 2180 3273 2232
rect 3325 2180 3337 2232
rect 3389 2223 3401 2232
rect 3453 2223 3465 2232
rect 3517 2223 3529 2232
rect 3581 2223 3593 2232
rect 3397 2189 3401 2223
rect 3389 2180 3401 2189
rect 3453 2180 3465 2189
rect 3517 2180 3529 2189
rect 3581 2180 3593 2189
rect 3645 2180 3651 2232
tri 3693 2224 3701 2232 ne
rect 3701 2224 3866 2232
tri 3866 2224 3885 2243 sw
tri 3701 2223 3702 2224 ne
rect 3702 2223 3885 2224
tri 3702 2189 3736 2223 ne
rect 3736 2189 3885 2223
tri 3736 2188 3737 2189 ne
rect 3737 2188 3885 2189
tri 3737 2180 3745 2188 ne
rect 3745 2180 3885 2188
tri 3745 2170 3755 2180 ne
rect 3203 2102 3209 2154
rect 3261 2102 3273 2154
rect 3325 2102 3337 2154
rect 3389 2102 3401 2154
rect 3453 2102 3465 2154
rect 3517 2102 3529 2154
rect 3581 2102 3593 2154
rect 3645 2102 3651 2154
rect 3203 2026 3209 2078
rect 3261 2026 3273 2078
rect 3325 2026 3337 2078
rect 3389 2069 3401 2078
rect 3453 2069 3465 2078
rect 3517 2069 3529 2078
rect 3581 2069 3593 2078
rect 3397 2035 3401 2069
rect 3389 2026 3401 2035
rect 3453 2026 3465 2035
rect 3517 2026 3529 2035
rect 3581 2026 3593 2035
rect 3645 2026 3651 2078
rect 3207 1881 3213 1933
rect 3265 1881 3277 1933
rect 3329 1931 3337 1933
rect 3338 1932 3364 1933
rect 3365 1931 3498 1933
rect 3329 1924 3498 1931
rect 3329 1890 3380 1924
rect 3414 1890 3452 1924
rect 3486 1890 3498 1924
rect 3329 1883 3498 1890
rect 3329 1881 3337 1883
rect 3338 1881 3364 1882
rect 3365 1881 3498 1883
rect 3203 1727 3209 1779
rect 3261 1727 3273 1779
rect 3325 1727 3333 1779
rect 3334 1728 3335 1778
rect 3363 1728 3364 1778
rect 3365 1770 3498 1779
rect 3365 1736 3380 1770
rect 3414 1736 3452 1770
rect 3486 1736 3498 1770
rect 3365 1727 3498 1736
rect 3207 1573 3213 1625
rect 3265 1573 3277 1625
rect 3329 1623 3337 1625
rect 3338 1624 3364 1625
rect 3365 1623 3498 1625
rect 3329 1616 3498 1623
rect 3329 1582 3380 1616
rect 3414 1582 3452 1616
rect 3486 1582 3498 1616
rect 3329 1575 3498 1582
rect 3329 1573 3337 1575
rect 3338 1573 3364 1574
rect 3365 1573 3498 1575
rect 3203 1419 3209 1471
rect 3261 1419 3273 1471
rect 3325 1419 3333 1471
rect 3334 1420 3335 1470
rect 3363 1420 3364 1470
rect 3365 1462 3498 1471
rect 3365 1428 3380 1462
rect 3414 1428 3452 1462
rect 3486 1428 3498 1462
rect 3365 1419 3498 1428
rect 3056 1350 3057 1376
rect 3058 1349 3112 1377
rect 3113 1350 3114 1376
rect 3056 1333 3114 1349
tri 3114 1333 3124 1343 sw
rect 3056 1317 3124 1333
tri 3124 1317 3140 1333 sw
rect 3056 1265 3213 1317
rect 3265 1265 3277 1317
rect 3329 1315 3337 1317
rect 3338 1316 3364 1317
rect 3365 1315 3498 1317
rect 3329 1308 3498 1315
rect 3329 1274 3380 1308
rect 3414 1274 3452 1308
rect 3486 1274 3498 1308
rect 3329 1267 3498 1274
rect 3329 1265 3337 1267
rect 3338 1265 3364 1266
rect 3365 1265 3498 1267
rect 348 1124 406 1162
rect 348 1090 360 1124
rect 394 1090 406 1124
rect 348 1052 406 1090
rect 466 1111 473 1163
rect 525 1111 537 1163
rect 589 1111 596 1163
rect 2574 1111 2581 1163
rect 2633 1111 2645 1163
rect 2697 1111 2704 1163
rect 3203 1111 3209 1163
rect 3261 1111 3273 1163
rect 3325 1111 3333 1163
rect 3334 1112 3335 1162
rect 3363 1112 3364 1162
rect 3365 1154 3498 1163
rect 3365 1120 3380 1154
rect 3414 1120 3452 1154
rect 3486 1120 3498 1154
rect 3365 1111 3498 1120
rect 466 1078 596 1111
rect 467 1076 595 1077
rect 348 1018 360 1052
rect 394 1018 406 1052
rect 348 980 406 1018
rect 348 946 360 980
rect 394 946 406 980
rect 467 1047 595 1048
rect 466 1009 596 1046
rect 466 957 473 1009
rect 525 957 537 1009
rect 589 957 596 1009
rect 3207 957 3213 1009
rect 3265 957 3277 1009
rect 3329 1007 3337 1009
rect 3338 1008 3364 1009
rect 3365 1007 3498 1009
rect 3329 1000 3498 1007
rect 3329 966 3380 1000
rect 3414 966 3452 1000
rect 3486 966 3498 1000
rect 3329 959 3498 966
rect 3329 957 3337 959
rect 3338 957 3364 958
rect 3365 957 3498 959
rect 348 908 406 946
rect 348 874 360 908
rect 394 874 406 908
rect 348 836 406 874
rect 3755 855 3885 2180
rect 3965 2177 3971 2229
rect 4023 2223 4035 2229
rect 4087 2223 4099 2229
rect 4151 2223 4163 2229
rect 4027 2189 4035 2223
rect 4023 2177 4035 2189
rect 4087 2177 4099 2189
rect 4151 2177 4163 2189
rect 4215 2177 4221 2229
rect 3965 2102 3971 2154
rect 4023 2102 4035 2154
rect 4087 2102 4099 2154
rect 4151 2102 4163 2154
rect 4215 2102 4221 2154
rect 3965 2023 3971 2075
rect 4023 2069 4035 2075
rect 4087 2069 4099 2075
rect 4151 2069 4163 2075
rect 4027 2035 4035 2069
rect 4023 2023 4035 2035
rect 4087 2023 4099 2035
rect 4151 2023 4163 2035
rect 4215 2023 4221 2075
rect 348 802 360 836
rect 394 802 406 836
rect 348 764 406 802
rect 466 803 473 855
rect 525 803 537 855
rect 589 803 596 855
rect 3203 803 3209 855
rect 3261 803 3273 855
rect 3325 803 3333 855
rect 3334 804 3335 854
rect 3363 804 3364 854
rect 3365 846 3498 855
rect 3365 812 3380 846
rect 3414 812 3452 846
rect 3486 812 3498 846
rect 3365 803 3498 812
rect 3755 803 3762 855
rect 3814 803 3826 855
rect 3878 803 3885 855
rect 466 771 596 803
rect 467 769 595 770
rect 348 730 360 764
rect 394 730 406 764
rect 348 692 406 730
rect 348 658 360 692
rect 394 658 406 692
rect 348 620 406 658
rect 467 740 595 741
rect 466 701 596 739
rect 466 649 473 701
rect 525 649 537 701
rect 589 649 596 701
rect 3207 649 3213 701
rect 3265 649 3277 701
rect 3329 699 3337 701
rect 3338 700 3364 701
rect 3365 699 3498 701
rect 3329 692 3498 699
rect 3329 658 3380 692
rect 3414 658 3452 692
rect 3486 658 3498 692
rect 3329 651 3498 658
rect 3329 649 3337 651
rect 3338 649 3364 650
rect 3365 649 3498 651
rect 348 586 360 620
rect 394 586 406 620
rect 348 548 406 586
rect 348 514 360 548
rect 394 514 406 548
rect 4286 547 4416 3684
tri 4416 3674 4426 3684 nw
tri 5132 3674 5142 3684 ne
rect 4768 3664 4826 3670
rect 4768 3637 4780 3664
rect 4814 3637 4826 3664
rect 4768 3585 4771 3637
rect 4823 3585 4826 3637
rect 4768 3573 4780 3585
rect 4814 3573 4826 3585
rect 4768 3521 4771 3573
rect 4823 3521 4826 3573
rect 4768 3520 4826 3521
rect 4768 3509 4780 3520
rect 4814 3509 4826 3520
rect 4768 3457 4771 3509
rect 4823 3457 4826 3509
rect 4768 3448 4826 3457
rect 4768 3445 4780 3448
rect 4814 3445 4826 3448
rect 4768 3393 4771 3445
rect 4823 3393 4826 3445
rect 4768 3381 4826 3393
rect 4768 3329 4771 3381
rect 4823 3329 4826 3381
rect 4768 3317 4826 3329
rect 4768 3265 4771 3317
rect 4823 3265 4826 3317
rect 4768 3253 4826 3265
rect 4768 3201 4771 3253
rect 4823 3201 4826 3253
rect 4768 3198 4780 3201
rect 4814 3198 4826 3201
rect 4768 3189 4826 3198
rect 4768 3137 4771 3189
rect 4823 3137 4826 3189
rect 4768 3126 4780 3137
rect 4814 3126 4826 3137
rect 4768 3125 4826 3126
rect 4768 3073 4771 3125
rect 4823 3073 4826 3125
rect 4768 3061 4780 3073
rect 4814 3061 4826 3073
rect 4768 3009 4771 3061
rect 4823 3009 4826 3061
rect 4768 2997 4780 3009
rect 4814 2997 4826 3009
rect 4768 2945 4771 2997
rect 4823 2945 4826 2997
rect 4768 2944 4826 2945
rect 4768 2933 4780 2944
rect 4814 2933 4826 2944
rect 4768 2881 4771 2933
rect 4823 2881 4826 2933
rect 4768 2872 4826 2881
rect 4768 2869 4780 2872
rect 4814 2869 4826 2872
rect 4768 2817 4771 2869
rect 4823 2817 4826 2869
rect 4768 2805 4826 2817
rect 4768 2753 4771 2805
rect 4823 2753 4826 2805
rect 4768 2728 4826 2753
rect 4768 2694 4780 2728
rect 4814 2694 4826 2728
rect 4768 2656 4826 2694
rect 4768 2622 4780 2656
rect 4814 2622 4826 2656
rect 4768 2584 4826 2622
rect 4768 2550 4780 2584
rect 4814 2550 4826 2584
rect 4768 2512 4826 2550
rect 4768 2478 4780 2512
rect 4814 2478 4826 2512
rect 4768 2440 4826 2478
rect 4768 2406 4780 2440
rect 4814 2406 4826 2440
rect 4768 2368 4826 2406
rect 4768 2334 4780 2368
rect 4814 2334 4826 2368
rect 4460 2177 4466 2229
rect 4518 2223 4530 2229
rect 4582 2223 4594 2229
rect 4646 2223 4658 2229
rect 4522 2189 4530 2223
rect 4518 2177 4530 2189
rect 4582 2177 4594 2189
rect 4646 2177 4658 2189
rect 4710 2177 4716 2229
rect 4460 2102 4466 2154
rect 4518 2102 4530 2154
rect 4582 2102 4594 2154
rect 4646 2102 4658 2154
rect 4710 2102 4716 2154
rect 4460 2023 4466 2075
rect 4518 2069 4530 2075
rect 4582 2069 4594 2075
rect 4646 2069 4658 2075
rect 4522 2035 4530 2069
rect 4518 2023 4530 2035
rect 4582 2023 4594 2035
rect 4646 2023 4658 2035
rect 4710 2023 4716 2075
rect 4768 1069 4826 2334
rect 4854 2177 4860 2229
rect 4912 2223 4924 2229
rect 4976 2223 4988 2229
rect 5040 2223 5052 2229
rect 4916 2189 4924 2223
rect 4912 2177 4924 2189
rect 4976 2177 4988 2189
rect 5040 2177 5052 2189
rect 5104 2177 5110 2229
rect 4854 2102 4860 2154
rect 4912 2102 4924 2154
rect 4976 2102 4988 2154
rect 5040 2102 5052 2154
rect 5104 2102 5110 2154
rect 4854 2023 4860 2075
rect 4912 2069 4924 2075
rect 4976 2069 4988 2075
rect 5040 2069 5052 2075
rect 4916 2035 4924 2069
rect 4912 2023 4924 2035
rect 4976 2023 4988 2035
rect 5040 2023 5052 2035
rect 5104 2023 5110 2075
rect 4768 1042 4769 1068
rect 4770 1041 4824 1069
rect 4825 1042 4826 1068
tri 4742 1009 4768 1035 se
rect 4768 1009 4826 1041
tri 4826 1009 4852 1035 sw
rect 4733 957 4739 1009
rect 4791 957 4803 1009
rect 4855 957 4861 1009
rect 348 476 406 514
rect 348 442 360 476
rect 394 442 406 476
rect 466 495 473 547
rect 525 495 537 547
rect 589 495 596 547
rect 3203 495 3209 547
rect 3261 495 3273 547
rect 3325 495 3333 547
rect 3334 496 3335 546
rect 3363 496 3364 546
rect 3365 538 3498 547
rect 3365 504 3380 538
rect 3414 504 3452 538
rect 3486 504 3498 538
rect 3365 495 3498 504
rect 4286 495 4293 547
rect 4345 495 4357 547
rect 4409 495 4416 547
rect 466 463 596 495
rect 467 461 595 462
rect 348 404 406 442
rect 348 370 360 404
rect 394 370 406 404
rect 348 332 406 370
rect 467 432 595 433
rect 466 393 596 431
rect 466 341 473 393
rect 525 341 537 393
rect 589 341 596 393
rect 3207 341 3213 393
rect 3265 341 3277 393
rect 3329 391 3337 393
rect 3338 392 3364 393
rect 3365 391 3498 393
rect 3329 384 3498 391
rect 3329 350 3380 384
rect 3414 350 3452 384
rect 3486 350 3498 384
rect 3329 343 3498 350
rect 3329 341 3337 343
rect 3338 341 3364 342
rect 3365 341 3498 343
rect 348 298 360 332
rect 394 298 406 332
rect 348 260 406 298
rect 348 226 360 260
rect 394 226 406 260
rect 5142 239 5272 3684
tri 5272 3674 5282 3684 nw
tri 5935 3674 5945 3684 ne
rect 5945 3674 6171 3684
tri 5945 3670 5949 3674 ne
rect 5949 3670 6171 3674
rect 5624 3664 5682 3670
tri 5949 3664 5955 3670 ne
rect 5955 3664 6171 3670
tri 6171 3664 6191 3684 nw
rect 6480 3664 6538 3670
rect 5624 3637 5636 3664
rect 5670 3637 5682 3664
rect 5624 3585 5627 3637
rect 5679 3585 5682 3637
tri 5955 3630 5989 3664 ne
rect 5989 3630 6137 3664
tri 6137 3630 6171 3664 nw
rect 6480 3637 6492 3664
rect 6526 3637 6538 3664
tri 5989 3621 5998 3630 ne
rect 5624 3573 5636 3585
rect 5670 3573 5682 3585
rect 5624 3521 5627 3573
rect 5679 3521 5682 3573
rect 5624 3520 5682 3521
rect 5624 3509 5636 3520
rect 5670 3509 5682 3520
rect 5624 3457 5627 3509
rect 5679 3457 5682 3509
rect 5624 3448 5682 3457
rect 5624 3445 5636 3448
rect 5670 3445 5682 3448
rect 5624 3393 5627 3445
rect 5679 3393 5682 3445
rect 5624 3381 5682 3393
rect 5624 3329 5627 3381
rect 5679 3329 5682 3381
rect 5624 3317 5682 3329
rect 5624 3265 5627 3317
rect 5679 3265 5682 3317
rect 5624 3253 5682 3265
rect 5624 3201 5627 3253
rect 5679 3201 5682 3253
rect 5624 3198 5636 3201
rect 5670 3198 5682 3201
rect 5624 3189 5682 3198
rect 5624 3137 5627 3189
rect 5679 3137 5682 3189
rect 5624 3126 5636 3137
rect 5670 3126 5682 3137
rect 5624 3125 5682 3126
rect 5624 3073 5627 3125
rect 5679 3073 5682 3125
rect 5624 3061 5636 3073
rect 5670 3061 5682 3073
rect 5624 3009 5627 3061
rect 5679 3009 5682 3061
rect 5624 2997 5636 3009
rect 5670 2997 5682 3009
rect 5624 2945 5627 2997
rect 5679 2945 5682 2997
rect 5624 2944 5682 2945
rect 5624 2933 5636 2944
rect 5670 2933 5682 2944
rect 5624 2881 5627 2933
rect 5679 2881 5682 2933
rect 5624 2872 5682 2881
rect 5624 2869 5636 2872
rect 5670 2869 5682 2872
rect 5624 2817 5627 2869
rect 5679 2817 5682 2869
rect 5624 2805 5682 2817
rect 5624 2753 5627 2805
rect 5679 2753 5682 2805
rect 5624 2728 5682 2753
rect 5624 2694 5636 2728
rect 5670 2694 5682 2728
rect 5624 2656 5682 2694
rect 5624 2622 5636 2656
rect 5670 2622 5682 2656
rect 5624 2584 5682 2622
rect 5624 2550 5636 2584
rect 5670 2550 5682 2584
rect 5624 2512 5682 2550
rect 5624 2478 5636 2512
rect 5670 2478 5682 2512
rect 5624 2440 5682 2478
rect 5624 2406 5636 2440
rect 5670 2406 5682 2440
rect 5624 2368 5682 2406
rect 5624 2334 5636 2368
rect 5670 2334 5682 2368
rect 5319 2177 5325 2229
rect 5377 2223 5389 2229
rect 5441 2223 5453 2229
rect 5505 2223 5517 2229
rect 5381 2189 5389 2223
rect 5377 2177 5389 2189
rect 5441 2177 5453 2189
rect 5505 2177 5517 2189
rect 5569 2177 5575 2229
rect 5319 2102 5325 2154
rect 5377 2102 5389 2154
rect 5441 2102 5453 2154
rect 5505 2102 5517 2154
rect 5569 2102 5575 2154
rect 5319 2023 5325 2075
rect 5377 2069 5389 2075
rect 5441 2069 5453 2075
rect 5505 2069 5517 2075
rect 5381 2035 5389 2069
rect 5377 2023 5389 2035
rect 5441 2023 5453 2035
rect 5505 2023 5517 2035
rect 5569 2023 5575 2075
rect 5624 761 5682 2334
rect 5713 2177 5719 2229
rect 5771 2223 5783 2229
rect 5835 2223 5847 2229
rect 5899 2223 5911 2229
rect 5775 2189 5783 2223
rect 5771 2177 5783 2189
rect 5835 2177 5847 2189
rect 5899 2177 5911 2189
rect 5963 2177 5969 2229
rect 5713 2102 5719 2154
rect 5771 2102 5783 2154
rect 5835 2102 5847 2154
rect 5899 2102 5911 2154
rect 5963 2102 5969 2154
rect 5713 2023 5719 2075
rect 5771 2069 5783 2075
rect 5835 2069 5847 2075
rect 5899 2069 5911 2075
rect 5775 2035 5783 2069
rect 5771 2023 5783 2035
rect 5835 2023 5847 2035
rect 5899 2023 5911 2035
rect 5963 2023 5969 2075
tri 5986 1951 5998 1963 se
rect 5998 1951 6128 3630
tri 6128 3621 6137 3630 nw
rect 6480 3585 6483 3637
rect 6535 3585 6538 3637
rect 6480 3573 6492 3585
rect 6526 3573 6538 3585
rect 6480 3521 6483 3573
rect 6535 3521 6538 3573
rect 6480 3520 6538 3521
rect 6480 3509 6492 3520
rect 6526 3509 6538 3520
rect 6480 3457 6483 3509
rect 6535 3457 6538 3509
rect 6480 3448 6538 3457
rect 6480 3445 6492 3448
rect 6526 3445 6538 3448
rect 6480 3393 6483 3445
rect 6535 3393 6538 3445
rect 6480 3381 6538 3393
rect 6480 3329 6483 3381
rect 6535 3329 6538 3381
rect 6480 3317 6538 3329
rect 6480 3265 6483 3317
rect 6535 3265 6538 3317
rect 6480 3253 6538 3265
rect 6480 3201 6483 3253
rect 6535 3201 6538 3253
rect 6480 3198 6492 3201
rect 6526 3198 6538 3201
rect 6480 3189 6538 3198
rect 6480 3137 6483 3189
rect 6535 3137 6538 3189
rect 6480 3126 6492 3137
rect 6526 3126 6538 3137
rect 6480 3125 6538 3126
rect 6480 3073 6483 3125
rect 6535 3073 6538 3125
rect 6480 3061 6492 3073
rect 6526 3061 6538 3073
rect 6480 3009 6483 3061
rect 6535 3009 6538 3061
rect 6480 2997 6492 3009
rect 6526 2997 6538 3009
rect 6480 2945 6483 2997
rect 6535 2945 6538 2997
rect 6480 2944 6538 2945
rect 6480 2933 6492 2944
rect 6526 2933 6538 2944
rect 6480 2881 6483 2933
rect 6535 2881 6538 2933
rect 6480 2872 6538 2881
rect 6480 2869 6492 2872
rect 6526 2869 6538 2872
rect 6480 2817 6483 2869
rect 6535 2817 6538 2869
rect 6480 2805 6538 2817
rect 6480 2753 6483 2805
rect 6535 2753 6538 2805
rect 6480 2728 6538 2753
rect 6480 2694 6492 2728
rect 6526 2694 6538 2728
rect 6480 2656 6538 2694
rect 6480 2622 6492 2656
rect 6526 2622 6538 2656
rect 6480 2584 6538 2622
rect 6480 2550 6492 2584
rect 6526 2550 6538 2584
rect 6480 2512 6538 2550
rect 6480 2478 6492 2512
rect 6526 2478 6538 2512
rect 6480 2440 6538 2478
rect 6480 2406 6492 2440
rect 6526 2406 6538 2440
rect 6480 2368 6538 2406
rect 6480 2334 6492 2368
rect 6526 2334 6538 2368
rect 6183 2177 6189 2229
rect 6241 2223 6253 2229
rect 6305 2223 6317 2229
rect 6369 2223 6381 2229
rect 6245 2189 6253 2223
rect 6241 2177 6253 2189
rect 6305 2177 6317 2189
rect 6369 2177 6381 2189
rect 6433 2177 6439 2229
rect 6183 2102 6189 2154
rect 6241 2102 6253 2154
rect 6305 2102 6317 2154
rect 6369 2102 6381 2154
rect 6433 2102 6439 2154
rect 6183 2023 6189 2075
rect 6241 2069 6253 2075
rect 6305 2069 6317 2075
rect 6369 2069 6381 2075
rect 6245 2035 6253 2069
rect 6241 2023 6253 2035
rect 6305 2023 6317 2035
rect 6369 2023 6381 2035
rect 6433 2023 6439 2075
tri 5968 1933 5986 1951 se
rect 5986 1933 6128 1951
rect 5801 1881 5807 1933
rect 5859 1881 5871 1933
rect 5923 1931 5938 1933
rect 5939 1932 5965 1933
rect 5966 1931 6128 1933
rect 5923 1904 6128 1931
rect 5923 1890 6114 1904
tri 6114 1890 6128 1904 nw
rect 5923 1883 6105 1890
rect 5923 1881 5938 1883
rect 5939 1881 5965 1882
rect 5966 1881 6105 1883
tri 6105 1881 6114 1890 nw
rect 5624 734 5625 760
rect 5626 733 5680 761
rect 5681 734 5682 760
tri 5607 710 5624 727 se
rect 5624 710 5682 733
tri 5682 710 5699 727 sw
tri 5598 701 5607 710 se
rect 5607 701 5699 710
tri 5699 701 5708 710 sw
rect 5589 649 5595 701
rect 5647 649 5659 701
rect 5711 649 5717 701
rect 6480 453 6538 2334
rect 7336 3664 7394 3670
rect 7336 3637 7348 3664
rect 7382 3637 7394 3664
rect 7336 3585 7339 3637
rect 7391 3585 7394 3637
rect 7336 3573 7348 3585
rect 7382 3573 7394 3585
rect 7336 3521 7339 3573
rect 7391 3521 7394 3573
rect 7336 3520 7394 3521
rect 7336 3509 7348 3520
rect 7382 3509 7394 3520
rect 7336 3457 7339 3509
rect 7391 3457 7394 3509
rect 7336 3448 7394 3457
rect 7336 3445 7348 3448
rect 7382 3445 7394 3448
rect 7336 3393 7339 3445
rect 7391 3393 7394 3445
rect 7336 3381 7394 3393
rect 7336 3329 7339 3381
rect 7391 3329 7394 3381
rect 7336 3317 7394 3329
rect 7336 3265 7339 3317
rect 7391 3265 7394 3317
rect 7336 3253 7394 3265
rect 7336 3201 7339 3253
rect 7391 3201 7394 3253
rect 7336 3198 7348 3201
rect 7382 3198 7394 3201
rect 7336 3189 7394 3198
rect 7336 3137 7339 3189
rect 7391 3137 7394 3189
rect 7336 3126 7348 3137
rect 7382 3126 7394 3137
rect 7336 3125 7394 3126
rect 7336 3073 7339 3125
rect 7391 3073 7394 3125
rect 7336 3061 7348 3073
rect 7382 3061 7394 3073
rect 7336 3009 7339 3061
rect 7391 3009 7394 3061
rect 7336 2997 7348 3009
rect 7382 2997 7394 3009
rect 7336 2945 7339 2997
rect 7391 2945 7394 2997
rect 7336 2944 7394 2945
rect 7336 2933 7348 2944
rect 7382 2933 7394 2944
rect 7336 2881 7339 2933
rect 7391 2881 7394 2933
rect 7336 2872 7394 2881
rect 7336 2869 7348 2872
rect 7382 2869 7394 2872
rect 7336 2817 7339 2869
rect 7391 2817 7394 2869
rect 7336 2805 7394 2817
rect 7336 2753 7339 2805
rect 7391 2753 7394 2805
rect 7336 2728 7394 2753
rect 7336 2694 7348 2728
rect 7382 2694 7394 2728
rect 7336 2656 7394 2694
rect 7336 2622 7348 2656
rect 7382 2622 7394 2656
rect 7336 2584 7394 2622
rect 7336 2550 7348 2584
rect 7382 2550 7394 2584
rect 7336 2512 7394 2550
rect 7336 2478 7348 2512
rect 7382 2478 7394 2512
rect 7336 2440 7394 2478
rect 7336 2406 7348 2440
rect 7382 2406 7394 2440
rect 7336 2368 7394 2406
rect 7336 2334 7348 2368
rect 7382 2334 7394 2368
rect 7336 2328 7394 2334
rect 8192 3664 8250 3670
rect 8192 3637 8204 3664
rect 8238 3637 8250 3664
rect 8192 3585 8195 3637
rect 8247 3585 8250 3637
rect 8192 3573 8204 3585
rect 8238 3573 8250 3585
rect 8192 3521 8195 3573
rect 8247 3521 8250 3573
rect 8192 3520 8250 3521
rect 8192 3509 8204 3520
rect 8238 3509 8250 3520
rect 8192 3457 8195 3509
rect 8247 3457 8250 3509
rect 8192 3448 8250 3457
rect 8192 3445 8204 3448
rect 8238 3445 8250 3448
rect 8192 3393 8195 3445
rect 8247 3393 8250 3445
rect 8192 3381 8250 3393
rect 8192 3329 8195 3381
rect 8247 3329 8250 3381
rect 8192 3317 8250 3329
rect 8192 3265 8195 3317
rect 8247 3265 8250 3317
rect 8192 3253 8250 3265
rect 8192 3201 8195 3253
rect 8247 3201 8250 3253
rect 8192 3198 8204 3201
rect 8238 3198 8250 3201
rect 8192 3189 8250 3198
rect 8192 3137 8195 3189
rect 8247 3137 8250 3189
rect 8192 3126 8204 3137
rect 8238 3126 8250 3137
rect 8192 3125 8250 3126
rect 8192 3073 8195 3125
rect 8247 3073 8250 3125
rect 8192 3061 8204 3073
rect 8238 3061 8250 3073
rect 8192 3009 8195 3061
rect 8247 3009 8250 3061
rect 8192 2997 8204 3009
rect 8238 2997 8250 3009
rect 8192 2945 8195 2997
rect 8247 2945 8250 2997
rect 8192 2944 8250 2945
rect 8192 2933 8204 2944
rect 8238 2933 8250 2944
rect 8192 2881 8195 2933
rect 8247 2881 8250 2933
rect 8192 2872 8250 2881
rect 8192 2869 8204 2872
rect 8238 2869 8250 2872
rect 8192 2817 8195 2869
rect 8247 2817 8250 2869
rect 8192 2805 8250 2817
rect 8192 2753 8195 2805
rect 8247 2753 8250 2805
rect 8192 2728 8250 2753
rect 8192 2694 8204 2728
rect 8238 2694 8250 2728
rect 8192 2656 8250 2694
rect 8192 2622 8204 2656
rect 8238 2622 8250 2656
rect 8192 2584 8250 2622
rect 8192 2550 8204 2584
rect 8238 2550 8250 2584
rect 8192 2512 8250 2550
rect 8192 2478 8204 2512
rect 8238 2478 8250 2512
rect 8192 2440 8250 2478
rect 8192 2406 8204 2440
rect 8238 2406 8250 2440
rect 8192 2368 8250 2406
rect 8192 2334 8204 2368
rect 8238 2334 8250 2368
rect 8192 2328 8250 2334
rect 9048 3664 9106 3670
rect 9048 3637 9060 3664
rect 9094 3637 9106 3664
rect 9048 3585 9051 3637
rect 9103 3585 9106 3637
rect 9048 3573 9060 3585
rect 9094 3573 9106 3585
rect 9048 3521 9051 3573
rect 9103 3521 9106 3573
rect 9048 3520 9106 3521
rect 9048 3509 9060 3520
rect 9094 3509 9106 3520
rect 9048 3457 9051 3509
rect 9103 3457 9106 3509
rect 9048 3448 9106 3457
rect 9048 3445 9060 3448
rect 9094 3445 9106 3448
rect 9048 3393 9051 3445
rect 9103 3393 9106 3445
rect 9048 3381 9106 3393
rect 9048 3329 9051 3381
rect 9103 3329 9106 3381
rect 9048 3317 9106 3329
rect 9048 3265 9051 3317
rect 9103 3265 9106 3317
rect 9048 3253 9106 3265
rect 9048 3201 9051 3253
rect 9103 3201 9106 3253
rect 9048 3198 9060 3201
rect 9094 3198 9106 3201
rect 9048 3189 9106 3198
rect 9048 3137 9051 3189
rect 9103 3137 9106 3189
rect 9048 3126 9060 3137
rect 9094 3126 9106 3137
rect 9048 3125 9106 3126
rect 9048 3073 9051 3125
rect 9103 3073 9106 3125
rect 9048 3061 9060 3073
rect 9094 3061 9106 3073
rect 9048 3009 9051 3061
rect 9103 3009 9106 3061
rect 9048 2997 9060 3009
rect 9094 2997 9106 3009
rect 9048 2945 9051 2997
rect 9103 2945 9106 2997
rect 9048 2944 9106 2945
rect 9048 2933 9060 2944
rect 9094 2933 9106 2944
rect 9048 2881 9051 2933
rect 9103 2881 9106 2933
rect 9048 2872 9106 2881
rect 9048 2869 9060 2872
rect 9094 2869 9106 2872
rect 9048 2817 9051 2869
rect 9103 2817 9106 2869
rect 9048 2805 9106 2817
rect 9048 2753 9051 2805
rect 9103 2753 9106 2805
rect 9048 2728 9106 2753
rect 9048 2694 9060 2728
rect 9094 2694 9106 2728
rect 9048 2656 9106 2694
rect 9048 2622 9060 2656
rect 9094 2622 9106 2656
rect 9048 2584 9106 2622
rect 9048 2550 9060 2584
rect 9094 2550 9106 2584
rect 9048 2512 9106 2550
rect 9048 2478 9060 2512
rect 9094 2478 9106 2512
rect 9048 2440 9106 2478
rect 9048 2406 9060 2440
rect 9094 2406 9106 2440
rect 9048 2368 9106 2406
rect 9048 2334 9060 2368
rect 9094 2334 9106 2368
rect 9048 2328 9106 2334
rect 9904 3664 9962 3670
rect 9904 3637 9916 3664
rect 9950 3637 9962 3664
rect 9904 3585 9907 3637
rect 9959 3585 9962 3637
rect 9904 3573 9916 3585
rect 9950 3573 9962 3585
rect 9904 3521 9907 3573
rect 9959 3521 9962 3573
rect 9904 3520 9962 3521
rect 9904 3509 9916 3520
rect 9950 3509 9962 3520
rect 9904 3457 9907 3509
rect 9959 3457 9962 3509
rect 9904 3448 9962 3457
rect 9904 3445 9916 3448
rect 9950 3445 9962 3448
rect 9904 3393 9907 3445
rect 9959 3393 9962 3445
rect 9904 3381 9962 3393
rect 9904 3329 9907 3381
rect 9959 3329 9962 3381
rect 9904 3317 9962 3329
rect 9904 3265 9907 3317
rect 9959 3265 9962 3317
rect 9904 3253 9962 3265
rect 9904 3201 9907 3253
rect 9959 3201 9962 3253
rect 9904 3198 9916 3201
rect 9950 3198 9962 3201
rect 9904 3189 9962 3198
rect 9904 3137 9907 3189
rect 9959 3137 9962 3189
rect 9904 3126 9916 3137
rect 9950 3126 9962 3137
rect 9904 3125 9962 3126
rect 9904 3073 9907 3125
rect 9959 3073 9962 3125
rect 9904 3061 9916 3073
rect 9950 3061 9962 3073
rect 9904 3009 9907 3061
rect 9959 3009 9962 3061
rect 9904 2997 9916 3009
rect 9950 2997 9962 3009
rect 9904 2945 9907 2997
rect 9959 2945 9962 2997
rect 9904 2944 9962 2945
rect 9904 2933 9916 2944
rect 9950 2933 9962 2944
rect 9904 2881 9907 2933
rect 9959 2881 9962 2933
rect 9904 2872 9962 2881
rect 9904 2869 9916 2872
rect 9950 2869 9962 2872
rect 9904 2817 9907 2869
rect 9959 2817 9962 2869
rect 9904 2805 9962 2817
rect 9904 2753 9907 2805
rect 9959 2753 9962 2805
rect 9904 2728 9962 2753
rect 9904 2694 9916 2728
rect 9950 2694 9962 2728
rect 9904 2656 9962 2694
rect 9904 2622 9916 2656
rect 9950 2622 9962 2656
rect 9904 2584 9962 2622
rect 9904 2550 9916 2584
rect 9950 2550 9962 2584
rect 9904 2512 9962 2550
rect 9904 2478 9916 2512
rect 9950 2478 9962 2512
rect 9904 2440 9962 2478
rect 9904 2406 9916 2440
rect 9950 2406 9962 2440
rect 9904 2368 9962 2406
rect 9904 2334 9916 2368
rect 9950 2334 9962 2368
rect 9904 2328 9962 2334
rect 10760 3664 10818 3670
rect 10760 3637 10772 3664
rect 10806 3637 10818 3664
rect 10760 3585 10763 3637
rect 10815 3585 10818 3637
rect 10760 3573 10772 3585
rect 10806 3573 10818 3585
rect 10760 3521 10763 3573
rect 10815 3521 10818 3573
rect 10760 3520 10818 3521
rect 10760 3509 10772 3520
rect 10806 3509 10818 3520
rect 10760 3457 10763 3509
rect 10815 3457 10818 3509
rect 10760 3448 10818 3457
rect 10760 3445 10772 3448
rect 10806 3445 10818 3448
rect 10760 3393 10763 3445
rect 10815 3393 10818 3445
rect 10760 3381 10818 3393
rect 10760 3329 10763 3381
rect 10815 3329 10818 3381
rect 10760 3317 10818 3329
rect 10760 3265 10763 3317
rect 10815 3265 10818 3317
rect 10760 3253 10818 3265
rect 10760 3201 10763 3253
rect 10815 3201 10818 3253
rect 10760 3198 10772 3201
rect 10806 3198 10818 3201
rect 10760 3189 10818 3198
rect 10760 3137 10763 3189
rect 10815 3137 10818 3189
rect 10760 3126 10772 3137
rect 10806 3126 10818 3137
rect 10760 3125 10818 3126
rect 10760 3073 10763 3125
rect 10815 3073 10818 3125
rect 10760 3061 10772 3073
rect 10806 3061 10818 3073
rect 10760 3009 10763 3061
rect 10815 3009 10818 3061
rect 10760 2997 10772 3009
rect 10806 2997 10818 3009
rect 10760 2945 10763 2997
rect 10815 2945 10818 2997
rect 10760 2944 10818 2945
rect 10760 2933 10772 2944
rect 10806 2933 10818 2944
rect 10760 2881 10763 2933
rect 10815 2881 10818 2933
rect 10760 2872 10818 2881
rect 10760 2869 10772 2872
rect 10806 2869 10818 2872
rect 10760 2817 10763 2869
rect 10815 2817 10818 2869
rect 10760 2805 10818 2817
rect 10760 2753 10763 2805
rect 10815 2753 10818 2805
rect 10760 2728 10818 2753
rect 10760 2694 10772 2728
rect 10806 2694 10818 2728
rect 10760 2656 10818 2694
rect 10760 2622 10772 2656
rect 10806 2622 10818 2656
rect 10760 2584 10818 2622
rect 10760 2550 10772 2584
rect 10806 2550 10818 2584
rect 10760 2512 10818 2550
rect 10760 2478 10772 2512
rect 10806 2478 10818 2512
rect 10760 2440 10818 2478
rect 10760 2406 10772 2440
rect 10806 2406 10818 2440
rect 10760 2368 10818 2406
rect 10760 2334 10772 2368
rect 10806 2334 10818 2368
rect 10760 2328 10818 2334
rect 10900 3646 10958 3684
rect 10900 3612 10912 3646
rect 10946 3612 10958 3646
rect 10900 3574 10958 3612
rect 10900 3540 10912 3574
rect 10946 3540 10958 3574
rect 10900 3502 10958 3540
rect 10900 3468 10912 3502
rect 10946 3468 10958 3502
rect 10900 3430 10958 3468
rect 10900 3396 10912 3430
rect 10946 3396 10958 3430
rect 10900 3358 10958 3396
rect 10900 3324 10912 3358
rect 10946 3324 10958 3358
rect 10900 3286 10958 3324
rect 10900 3252 10912 3286
rect 10946 3252 10958 3286
rect 10900 3214 10958 3252
rect 10900 3180 10912 3214
rect 10946 3180 10958 3214
rect 10900 3142 10958 3180
rect 10900 3108 10912 3142
rect 10946 3108 10958 3142
rect 10900 3070 10958 3108
rect 10900 3036 10912 3070
rect 10946 3036 10958 3070
rect 10900 2998 10958 3036
rect 10900 2964 10912 2998
rect 10946 2964 10958 2998
rect 10900 2926 10958 2964
rect 10900 2892 10912 2926
rect 10946 2892 10958 2926
rect 10900 2854 10958 2892
rect 10900 2820 10912 2854
rect 10946 2820 10958 2854
rect 10900 2782 10958 2820
rect 10900 2748 10912 2782
rect 10946 2748 10958 2782
rect 10900 2710 10958 2748
rect 10900 2679 10912 2710
rect 10946 2679 10958 2710
rect 10900 2627 10904 2679
rect 10956 2627 10958 2679
rect 10900 2615 10912 2627
rect 10946 2615 10958 2627
rect 10900 2563 10904 2615
rect 10956 2563 10958 2615
rect 10900 2550 10912 2563
rect 10946 2550 10958 2563
rect 10900 2498 10904 2550
rect 10956 2498 10958 2550
rect 10900 2494 10958 2498
rect 10900 2485 10912 2494
rect 10946 2485 10958 2494
rect 10900 2433 10904 2485
rect 10956 2433 10958 2485
rect 10900 2422 10958 2433
rect 10900 2420 10912 2422
rect 10946 2420 10958 2422
rect 10900 2368 10904 2420
rect 10956 2368 10958 2420
rect 10900 2355 10958 2368
rect 10900 2303 10904 2355
rect 10956 2303 10958 2355
tri 10879 2260 10900 2281 se
rect 10900 2260 10958 2303
tri 10862 2243 10879 2260 se
rect 10879 2243 10958 2260
tri 10848 2229 10862 2243 se
rect 10862 2229 10958 2243
rect 6570 2177 6576 2229
rect 6628 2223 6640 2229
rect 6692 2223 6704 2229
rect 6628 2189 6629 2223
rect 6692 2189 6701 2223
rect 6628 2177 6640 2189
rect 6692 2177 6704 2189
rect 6756 2177 6768 2229
rect 6820 2177 6832 2229
rect 6884 2177 6896 2229
rect 6948 2223 6960 2229
rect 7012 2223 7024 2229
rect 7076 2223 7088 2229
rect 7140 2223 7152 2229
rect 7204 2223 7216 2229
rect 7268 2223 7280 2229
rect 6951 2189 6960 2223
rect 7023 2189 7024 2223
rect 7204 2189 7205 2223
rect 7268 2189 7277 2223
rect 6948 2177 6960 2189
rect 7012 2177 7024 2189
rect 7076 2177 7088 2189
rect 7140 2177 7152 2189
rect 7204 2177 7216 2189
rect 7268 2177 7280 2189
rect 7332 2177 7344 2229
rect 7396 2177 7408 2229
rect 7460 2177 7472 2229
rect 7524 2223 7536 2229
rect 7588 2223 7600 2229
rect 7652 2223 7664 2229
rect 7716 2223 7728 2229
rect 7780 2223 7792 2229
rect 7844 2223 7856 2229
rect 7527 2189 7536 2223
rect 7599 2189 7600 2223
rect 7780 2189 7781 2223
rect 7844 2189 7853 2223
rect 7524 2177 7536 2189
rect 7588 2177 7600 2189
rect 7652 2177 7664 2189
rect 7716 2177 7728 2189
rect 7780 2177 7792 2189
rect 7844 2177 7856 2189
rect 7908 2177 7920 2229
rect 7972 2177 7984 2229
rect 8036 2177 8048 2229
rect 8100 2223 8112 2229
rect 8164 2223 8176 2229
rect 8228 2223 8240 2229
rect 8292 2223 8304 2229
rect 8356 2223 8368 2229
rect 8420 2223 8432 2229
rect 8103 2189 8112 2223
rect 8175 2189 8176 2223
rect 8356 2189 8357 2223
rect 8420 2189 8429 2223
rect 8100 2177 8112 2189
rect 8164 2177 8176 2189
rect 8228 2177 8240 2189
rect 8292 2177 8304 2189
rect 8356 2177 8368 2189
rect 8420 2177 8432 2189
rect 8484 2177 8496 2229
rect 8548 2177 8560 2229
rect 8612 2177 8624 2229
rect 8676 2223 8688 2229
rect 8740 2223 8752 2229
rect 8804 2223 8816 2229
rect 8868 2223 8880 2229
rect 8932 2223 8944 2229
rect 8996 2223 9008 2229
rect 8679 2189 8688 2223
rect 8751 2189 8752 2223
rect 8932 2189 8933 2223
rect 8996 2189 9005 2223
rect 8676 2177 8688 2189
rect 8740 2177 8752 2189
rect 8804 2177 8816 2189
rect 8868 2177 8880 2189
rect 8932 2177 8944 2189
rect 8996 2177 9008 2189
rect 9060 2177 9072 2229
rect 9124 2177 9136 2229
rect 9188 2177 9200 2229
rect 9252 2223 9264 2229
rect 9316 2223 9328 2229
rect 9380 2223 9392 2229
rect 9444 2223 9456 2229
rect 9508 2223 9520 2229
rect 9572 2223 9584 2229
rect 9255 2189 9264 2223
rect 9327 2189 9328 2223
rect 9508 2189 9509 2223
rect 9572 2189 9581 2223
rect 9252 2177 9264 2189
rect 9316 2177 9328 2189
rect 9380 2177 9392 2189
rect 9444 2177 9456 2189
rect 9508 2177 9520 2189
rect 9572 2177 9584 2189
rect 9636 2177 9648 2229
rect 9700 2177 9712 2229
rect 9764 2177 9776 2229
rect 9828 2223 9840 2229
rect 9892 2223 9904 2229
rect 9956 2223 9968 2229
rect 10020 2223 10032 2229
rect 10084 2223 10096 2229
rect 10148 2223 10160 2229
rect 9831 2189 9840 2223
rect 9903 2189 9904 2223
rect 10084 2189 10085 2223
rect 10148 2189 10157 2223
rect 9828 2177 9840 2189
rect 9892 2177 9904 2189
rect 9956 2177 9968 2189
rect 10020 2177 10032 2189
rect 10084 2177 10096 2189
rect 10148 2177 10160 2189
rect 10212 2177 10224 2229
rect 10276 2177 10288 2229
rect 10340 2177 10352 2229
rect 10404 2223 10416 2229
rect 10468 2223 10480 2229
rect 10532 2223 10544 2229
rect 10596 2223 10608 2229
rect 10660 2223 10672 2229
rect 10724 2223 10736 2229
rect 10407 2189 10416 2223
rect 10479 2189 10480 2223
rect 10660 2189 10661 2223
rect 10724 2189 10733 2223
rect 10404 2177 10416 2189
rect 10468 2177 10480 2189
rect 10532 2177 10544 2189
rect 10596 2177 10608 2189
rect 10660 2177 10672 2189
rect 10724 2177 10736 2189
rect 10788 2177 10800 2229
rect 10852 2177 10864 2229
rect 10916 2177 10958 2229
rect 6570 2102 6576 2154
rect 6628 2144 6641 2154
rect 6693 2144 6706 2154
rect 6693 2110 6698 2144
rect 6628 2102 6641 2110
rect 6693 2102 6706 2110
rect 6758 2102 6771 2154
rect 6823 2102 6836 2154
rect 6888 2102 6901 2154
rect 6953 2102 6966 2154
rect 7018 2144 7031 2154
rect 7083 2144 7096 2154
rect 7148 2144 7161 2154
rect 7213 2144 7226 2154
rect 7278 2144 7291 2154
rect 7024 2110 7031 2144
rect 7278 2110 7282 2144
rect 7018 2102 7031 2110
rect 7083 2102 7096 2110
rect 7148 2102 7161 2110
rect 7213 2102 7226 2110
rect 7278 2102 7291 2110
rect 7343 2102 7355 2154
rect 7407 2102 7419 2154
rect 7471 2102 7483 2154
rect 7535 2102 7547 2154
rect 7599 2144 7611 2154
rect 7663 2144 7675 2154
rect 7727 2144 7739 2154
rect 7791 2144 7803 2154
rect 7855 2144 7867 2154
rect 7608 2110 7611 2144
rect 7791 2110 7792 2144
rect 7855 2110 7864 2144
rect 7599 2102 7611 2110
rect 7663 2102 7675 2110
rect 7727 2102 7739 2110
rect 7791 2102 7803 2110
rect 7855 2102 7867 2110
rect 7919 2102 7931 2154
rect 7983 2102 7995 2154
rect 8047 2102 8059 2154
rect 8111 2144 8123 2154
rect 8175 2144 8187 2154
rect 8239 2144 8251 2154
rect 8303 2144 8315 2154
rect 8367 2144 8379 2154
rect 8431 2144 8443 2154
rect 8114 2110 8123 2144
rect 8186 2110 8187 2144
rect 8367 2110 8368 2144
rect 8431 2110 8440 2144
rect 8111 2102 8123 2110
rect 8175 2102 8187 2110
rect 8239 2102 8251 2110
rect 8303 2102 8315 2110
rect 8367 2102 8379 2110
rect 8431 2102 8443 2110
rect 8495 2102 8507 2154
rect 8559 2102 8571 2154
rect 8623 2102 8635 2154
rect 8687 2144 8699 2154
rect 8751 2144 8763 2154
rect 8815 2144 8827 2154
rect 8879 2144 8891 2154
rect 8943 2144 8955 2154
rect 9007 2144 9019 2154
rect 8690 2110 8699 2144
rect 8762 2110 8763 2144
rect 8943 2110 8944 2144
rect 9007 2110 9016 2144
rect 8687 2102 8699 2110
rect 8751 2102 8763 2110
rect 8815 2102 8827 2110
rect 8879 2102 8891 2110
rect 8943 2102 8955 2110
rect 9007 2102 9019 2110
rect 9071 2102 9083 2154
rect 9135 2102 9147 2154
rect 9199 2102 9211 2154
rect 9263 2144 9275 2154
rect 9327 2144 9339 2154
rect 9391 2144 9403 2154
rect 9455 2144 9467 2154
rect 9519 2144 9531 2154
rect 9583 2144 9595 2154
rect 9266 2110 9275 2144
rect 9338 2110 9339 2144
rect 9519 2110 9520 2144
rect 9583 2110 9592 2144
rect 9263 2102 9275 2110
rect 9327 2102 9339 2110
rect 9391 2102 9403 2110
rect 9455 2102 9467 2110
rect 9519 2102 9531 2110
rect 9583 2102 9595 2110
rect 9647 2102 9659 2154
rect 9711 2102 9723 2154
rect 9775 2102 9787 2154
rect 9839 2144 9851 2154
rect 9903 2144 9915 2154
rect 9967 2144 9979 2154
rect 10031 2144 10043 2154
rect 10095 2144 10107 2154
rect 10159 2144 10171 2154
rect 9842 2110 9851 2144
rect 9914 2110 9915 2144
rect 10095 2110 10096 2144
rect 10159 2110 10168 2144
rect 9839 2102 9851 2110
rect 9903 2102 9915 2110
rect 9967 2102 9979 2110
rect 10031 2102 10043 2110
rect 10095 2102 10107 2110
rect 10159 2102 10171 2110
rect 10223 2102 10235 2154
rect 10287 2102 10299 2154
rect 10351 2102 10363 2154
rect 10415 2144 10427 2154
rect 10479 2144 10491 2154
rect 10543 2144 10555 2154
rect 10607 2144 10619 2154
rect 10671 2144 10683 2154
rect 10735 2144 10747 2154
rect 10418 2110 10427 2144
rect 10490 2110 10491 2144
rect 10671 2110 10672 2144
rect 10735 2110 10744 2144
rect 10415 2102 10427 2110
rect 10479 2102 10491 2110
rect 10543 2102 10555 2110
rect 10607 2102 10619 2110
rect 10671 2102 10683 2110
rect 10735 2102 10747 2110
rect 10799 2102 10811 2154
rect 10863 2102 10875 2154
rect 10927 2150 10933 2154
rect 10927 2104 10934 2150
rect 10927 2102 10933 2104
rect 6576 2023 6582 2075
rect 6634 2069 6646 2075
rect 6698 2069 6710 2075
rect 6762 2069 6774 2075
rect 6698 2035 6701 2069
rect 6762 2035 6773 2069
rect 6634 2023 6646 2035
rect 6698 2023 6710 2035
rect 6762 2023 6774 2035
rect 6826 2023 6838 2075
rect 6890 2023 6902 2075
rect 6954 2023 6966 2075
rect 7018 2069 7030 2075
rect 7082 2069 7094 2075
rect 7146 2069 7158 2075
rect 7210 2069 7222 2075
rect 7274 2069 7286 2075
rect 7338 2069 7350 2075
rect 7023 2035 7030 2069
rect 7274 2035 7277 2069
rect 7338 2035 7349 2069
rect 7018 2023 7030 2035
rect 7082 2023 7094 2035
rect 7146 2023 7158 2035
rect 7210 2023 7222 2035
rect 7274 2023 7286 2035
rect 7338 2023 7350 2035
rect 7402 2023 7414 2075
rect 7466 2023 7478 2075
rect 7530 2023 7542 2075
rect 7594 2069 7606 2075
rect 7658 2069 7670 2075
rect 7722 2069 7734 2075
rect 7786 2069 7798 2075
rect 7850 2069 7862 2075
rect 7914 2069 7926 2075
rect 7599 2035 7606 2069
rect 7850 2035 7853 2069
rect 7914 2035 7925 2069
rect 7594 2023 7606 2035
rect 7658 2023 7670 2035
rect 7722 2023 7734 2035
rect 7786 2023 7798 2035
rect 7850 2023 7862 2035
rect 7914 2023 7926 2035
rect 7978 2023 7990 2075
rect 8042 2023 8054 2075
rect 8106 2023 8118 2075
rect 8170 2069 8182 2075
rect 8234 2069 8246 2075
rect 8298 2069 8310 2075
rect 8362 2069 8374 2075
rect 8426 2069 8438 2075
rect 8490 2069 8502 2075
rect 8175 2035 8182 2069
rect 8426 2035 8429 2069
rect 8490 2035 8501 2069
rect 8170 2023 8182 2035
rect 8234 2023 8246 2035
rect 8298 2023 8310 2035
rect 8362 2023 8374 2035
rect 8426 2023 8438 2035
rect 8490 2023 8502 2035
rect 8554 2023 8566 2075
rect 8618 2023 8630 2075
rect 8682 2023 8694 2075
rect 8746 2069 8758 2075
rect 8810 2069 8822 2075
rect 8874 2069 8886 2075
rect 8938 2069 8950 2075
rect 9002 2069 9014 2075
rect 9066 2069 9078 2075
rect 8751 2035 8758 2069
rect 9002 2035 9005 2069
rect 9066 2035 9077 2069
rect 8746 2023 8758 2035
rect 8810 2023 8822 2035
rect 8874 2023 8886 2035
rect 8938 2023 8950 2035
rect 9002 2023 9014 2035
rect 9066 2023 9078 2035
rect 9130 2023 9142 2075
rect 9194 2023 9206 2075
rect 9258 2023 9270 2075
rect 9322 2069 9334 2075
rect 9386 2069 9398 2075
rect 9450 2069 9462 2075
rect 9514 2069 9526 2075
rect 9578 2069 9590 2075
rect 9642 2069 9654 2075
rect 9327 2035 9334 2069
rect 9578 2035 9581 2069
rect 9642 2035 9653 2069
rect 9322 2023 9334 2035
rect 9386 2023 9398 2035
rect 9450 2023 9462 2035
rect 9514 2023 9526 2035
rect 9578 2023 9590 2035
rect 9642 2023 9654 2035
rect 9706 2023 9718 2075
rect 9770 2023 9782 2075
rect 9834 2023 9846 2075
rect 9898 2069 9910 2075
rect 9962 2069 9974 2075
rect 10026 2069 10038 2075
rect 10090 2069 10102 2075
rect 10154 2069 10166 2075
rect 10218 2069 10230 2075
rect 9903 2035 9910 2069
rect 10154 2035 10157 2069
rect 10218 2035 10229 2069
rect 9898 2023 9910 2035
rect 9962 2023 9974 2035
rect 10026 2023 10038 2035
rect 10090 2023 10102 2035
rect 10154 2023 10166 2035
rect 10218 2023 10230 2035
rect 10282 2023 10294 2075
rect 10346 2023 10358 2075
rect 10410 2023 10422 2075
rect 10474 2069 10486 2075
rect 10538 2069 10550 2075
rect 10602 2069 10614 2075
rect 10666 2069 10678 2075
rect 10730 2069 10742 2075
rect 10794 2069 10806 2075
rect 10479 2035 10486 2069
rect 10730 2035 10733 2069
rect 10794 2035 10805 2069
rect 10474 2023 10486 2035
rect 10538 2023 10550 2035
rect 10602 2023 10614 2035
rect 10666 2023 10678 2035
rect 10730 2023 10742 2035
rect 10794 2023 10806 2035
rect 10858 2023 10870 2075
rect 10922 2023 10928 2075
tri 10960 1779 10986 1805 se
rect 10986 1779 11114 5910
tri 12053 5897 12066 5910 ne
rect 12066 5897 12115 5910
tri 12115 5897 12140 5922 sw
tri 14645 5897 14670 5922 se
rect 14670 5897 14742 5922
tri 12066 5888 12075 5897 ne
rect 12075 5888 14298 5897
tri 12075 5882 12081 5888 ne
rect 12081 5882 14298 5888
rect 11612 5830 11619 5882
rect 11671 5830 11683 5882
rect 11735 5830 11742 5882
tri 12081 5854 12109 5882 ne
rect 12109 5854 14298 5882
tri 12109 5850 12113 5854 ne
rect 12113 5850 14298 5854
tri 12113 5845 12118 5850 ne
rect 12118 5845 14298 5850
rect 14299 5846 14300 5896
rect 14328 5846 14329 5896
rect 14330 5845 14355 5897
rect 14407 5845 14419 5897
rect 14471 5845 14479 5897
rect 14480 5846 14481 5896
rect 14509 5846 14510 5896
rect 14511 5892 14742 5897
rect 14511 5888 14738 5892
tri 14738 5888 14742 5892 nw
rect 14511 5854 14526 5888
rect 14560 5854 14598 5888
rect 14632 5854 14700 5888
rect 14511 5850 14700 5854
tri 14700 5850 14738 5888 nw
rect 14511 5848 14698 5850
tri 14698 5848 14700 5850 nw
rect 14511 5845 14695 5848
tri 14695 5845 14698 5848 nw
tri 14788 5845 14791 5848 se
rect 14791 5845 14843 6282
tri 14779 5836 14788 5845 se
rect 14788 5836 14843 5845
rect 11612 5810 11742 5830
tri 14759 5816 14779 5836 se
rect 14779 5826 14843 5836
rect 14779 5816 14833 5826
tri 14833 5816 14843 5826 nw
tri 14753 5810 14759 5816 se
rect 14759 5810 14795 5816
tri 14752 5809 14753 5810 se
rect 14753 5809 14795 5810
rect 11613 5808 11741 5809
tri 14751 5808 14752 5809 se
rect 14752 5808 14795 5809
tri 14723 5780 14751 5808 se
rect 14751 5780 14795 5808
rect 11613 5779 11741 5780
tri 14722 5779 14723 5780 se
rect 14723 5779 14795 5780
tri 14721 5778 14722 5779 se
rect 14722 5778 14795 5779
tri 14795 5778 14833 5816 nw
rect 11612 5743 11742 5778
tri 14717 5774 14721 5778 se
rect 14721 5774 14791 5778
tri 14791 5774 14795 5778 nw
tri 14695 5752 14717 5774 se
rect 14717 5752 14761 5774
tri 14687 5744 14695 5752 se
rect 14695 5744 14761 5752
tri 14761 5744 14791 5774 nw
tri 14686 5743 14687 5744 se
rect 14687 5743 14760 5744
tri 14760 5743 14761 5744 nw
rect 11612 5691 11619 5743
rect 11671 5691 11683 5743
rect 11735 5691 11742 5743
rect 14353 5691 14359 5743
rect 14411 5691 14423 5743
rect 14475 5741 14483 5743
rect 14484 5742 14510 5743
rect 14511 5741 14755 5743
rect 14475 5738 14755 5741
tri 14755 5738 14760 5743 nw
rect 14475 5734 14723 5738
rect 14475 5700 14526 5734
rect 14560 5700 14598 5734
rect 14632 5706 14723 5734
tri 14723 5706 14755 5738 nw
tri 14839 5706 14871 5738 se
rect 14871 5716 14923 6342
rect 14871 5706 14913 5716
tri 14913 5706 14923 5716 nw
rect 14632 5700 14708 5706
rect 14475 5693 14708 5700
rect 14475 5691 14483 5693
rect 14484 5691 14510 5692
rect 14511 5691 14708 5693
tri 14708 5691 14723 5706 nw
tri 14824 5691 14839 5706 se
rect 14839 5691 14879 5706
rect 11494 5599 11540 5611
rect 11494 5565 11500 5599
rect 11534 5565 11540 5599
rect 11494 5525 11540 5565
rect 11494 5491 11500 5525
rect 11534 5491 11540 5525
rect 11612 5589 11742 5691
tri 14805 5672 14824 5691 se
rect 14824 5672 14879 5691
tri 14879 5672 14913 5706 nw
tri 14797 5664 14805 5672 se
rect 14805 5664 14871 5672
tri 14871 5664 14879 5672 nw
tri 14767 5634 14797 5664 se
rect 14797 5634 14841 5664
tri 14841 5634 14871 5664 nw
tri 14733 5600 14767 5634 se
rect 14767 5600 14807 5634
tri 14807 5600 14841 5634 nw
tri 14723 5590 14733 5600 se
rect 14733 5590 14797 5600
tri 14797 5590 14807 5600 nw
tri 14722 5589 14723 5590 se
rect 14723 5589 14796 5590
tri 14796 5589 14797 5590 nw
rect 11612 5537 11619 5589
rect 11671 5537 11683 5589
rect 11735 5537 11742 5589
rect 14349 5537 14355 5589
rect 14407 5537 14419 5589
rect 14471 5537 14479 5589
rect 14480 5538 14481 5588
rect 14509 5538 14510 5588
rect 14511 5580 14769 5589
rect 14511 5546 14526 5580
rect 14560 5546 14598 5580
rect 14632 5562 14769 5580
tri 14769 5562 14796 5589 nw
tri 14924 5562 14951 5589 se
rect 14951 5567 15003 6392
rect 14951 5562 14998 5567
tri 14998 5562 15003 5567 nw
rect 14632 5546 14744 5562
rect 14511 5537 14744 5546
tri 14744 5537 14769 5562 nw
tri 14899 5537 14924 5562 se
rect 14924 5537 14964 5562
rect 11612 5502 11742 5537
tri 14890 5528 14899 5537 se
rect 14899 5528 14964 5537
tri 14964 5528 14998 5562 nw
tri 14877 5515 14890 5528 se
rect 14890 5515 14951 5528
tri 14951 5515 14964 5528 nw
tri 14864 5502 14877 5515 se
rect 14877 5502 14926 5515
tri 14863 5501 14864 5502 se
rect 14864 5501 14926 5502
rect 11613 5500 11741 5501
tri 14862 5500 14863 5501 se
rect 14863 5500 14926 5501
rect 11494 5451 11540 5491
tri 14852 5490 14862 5500 se
rect 14862 5490 14926 5500
tri 14926 5490 14951 5515 nw
tri 14834 5472 14852 5490 se
rect 14852 5472 14892 5490
rect 11494 5417 11500 5451
rect 11534 5417 11540 5451
rect 11494 5377 11540 5417
rect 11494 5343 11500 5377
rect 11534 5343 11540 5377
rect 11494 5303 11540 5343
rect 11494 5269 11500 5303
rect 11534 5269 11540 5303
rect 11494 5229 11540 5269
rect 11494 5195 11500 5229
rect 11534 5195 11540 5229
rect 11494 5155 11540 5195
rect 11494 5121 11500 5155
rect 11534 5121 11540 5155
rect 11494 5081 11540 5121
rect 11494 5047 11500 5081
rect 11534 5047 11540 5081
rect 11494 5007 11540 5047
rect 11494 4973 11500 5007
rect 11534 4973 11540 5007
rect 11494 4933 11540 4973
rect 11494 4899 11500 4933
rect 11534 4899 11540 4933
rect 11494 4859 11540 4899
rect 11613 5471 11741 5472
tri 14833 5471 14834 5472 se
rect 14834 5471 14892 5472
tri 14832 5470 14833 5471 se
rect 14833 5470 14892 5471
rect 11612 5435 11742 5470
tri 14818 5456 14832 5470 se
rect 14832 5456 14892 5470
tri 14892 5456 14926 5490 nw
tri 14811 5449 14818 5456 se
rect 14818 5449 14885 5456
tri 14885 5449 14892 5456 nw
tri 14806 5444 14811 5449 se
rect 14811 5444 14880 5449
tri 14880 5444 14885 5449 nw
tri 15026 5444 15031 5449 se
rect 15031 5444 15083 6532
tri 14803 5441 14806 5444 se
rect 14806 5441 14877 5444
tri 14877 5441 14880 5444 nw
tri 15023 5441 15026 5444 se
rect 15026 5441 15083 5444
tri 14797 5435 14803 5441 se
rect 14803 5435 14871 5441
tri 14871 5435 14877 5441 nw
tri 15017 5435 15023 5441 se
rect 15023 5435 15083 5441
rect 11612 5383 11619 5435
rect 11671 5383 11683 5435
rect 11735 5383 11742 5435
rect 14353 5383 14359 5435
rect 14411 5383 14423 5435
rect 14475 5433 14483 5435
rect 14484 5434 14510 5435
rect 14511 5433 14854 5435
rect 14475 5426 14854 5433
rect 14475 5392 14526 5426
rect 14560 5392 14598 5426
rect 14632 5418 14854 5426
tri 14854 5418 14871 5435 nw
tri 15000 5418 15017 5435 se
rect 15017 5427 15083 5435
rect 15017 5418 15074 5427
tri 15074 5418 15083 5427 nw
rect 14632 5392 14820 5418
rect 14475 5385 14820 5392
rect 14475 5383 14483 5385
rect 14511 5384 14820 5385
tri 14820 5384 14854 5418 nw
tri 14966 5384 15000 5418 se
rect 15000 5384 15040 5418
tri 15040 5384 15074 5418 nw
rect 14484 5383 14510 5384
rect 14511 5383 14819 5384
tri 14819 5383 14820 5384 nw
tri 14965 5383 14966 5384 se
rect 14966 5383 15031 5384
rect 11612 5281 11742 5383
tri 14957 5375 14965 5383 se
rect 14965 5375 15031 5383
tri 15031 5375 15040 5384 nw
tri 14928 5346 14957 5375 se
rect 14957 5346 15002 5375
tri 15002 5346 15031 5375 nw
tri 14894 5312 14928 5346 se
rect 14928 5312 14968 5346
tri 14968 5312 15002 5346 nw
tri 14891 5309 14894 5312 se
rect 14894 5309 14965 5312
tri 14965 5309 14968 5312 nw
tri 14883 5301 14891 5309 se
rect 14891 5301 14957 5309
tri 14957 5301 14965 5309 nw
tri 15103 5301 15111 5309 se
rect 15111 5301 15163 6672
tri 14863 5281 14883 5301 se
rect 14883 5281 14937 5301
tri 14937 5281 14957 5301 nw
tri 15083 5281 15103 5301 se
rect 15103 5287 15163 5301
rect 15103 5281 15150 5287
rect 11612 5229 11619 5281
rect 11671 5229 11683 5281
rect 11735 5229 11742 5281
rect 14349 5229 14355 5281
rect 14407 5229 14419 5281
rect 14471 5229 14479 5281
rect 14480 5230 14481 5280
rect 14509 5230 14510 5280
rect 14511 5274 14930 5281
tri 14930 5274 14937 5281 nw
tri 15076 5274 15083 5281 se
rect 15083 5274 15150 5281
tri 15150 5274 15163 5287 nw
rect 14511 5272 14896 5274
rect 14511 5238 14526 5272
rect 14560 5238 14598 5272
rect 14632 5240 14896 5272
tri 14896 5240 14930 5274 nw
tri 15042 5240 15076 5274 se
rect 15076 5240 15116 5274
tri 15116 5240 15150 5274 nw
rect 14632 5238 14891 5240
rect 14511 5235 14891 5238
tri 14891 5235 14896 5240 nw
tri 15037 5235 15042 5240 se
rect 15042 5235 15111 5240
tri 15111 5235 15116 5240 nw
rect 14511 5229 14885 5235
tri 14885 5229 14891 5235 nw
tri 15031 5229 15037 5235 se
rect 15037 5229 15078 5235
rect 11612 5196 11742 5229
tri 15022 5220 15031 5229 se
rect 15031 5220 15078 5229
tri 15004 5202 15022 5220 se
rect 15022 5202 15078 5220
tri 15078 5202 15111 5235 nw
tri 14998 5196 15004 5202 se
rect 15004 5196 15045 5202
rect 11612 5169 11613 5195
rect 11614 5168 11740 5196
tri 14997 5195 14998 5196 se
rect 14998 5195 15045 5196
rect 11741 5169 11742 5195
tri 14971 5169 14997 5195 se
rect 14997 5169 15045 5195
tri 15045 5169 15078 5202 nw
tri 14970 5168 14971 5169 se
rect 14971 5168 15044 5169
tri 15044 5168 15045 5169 nw
tri 15190 5168 15191 5169 se
rect 15191 5168 15243 6804
rect 11612 5127 11742 5168
tri 14963 5161 14970 5168 se
rect 14970 5161 15037 5168
tri 15037 5161 15044 5168 nw
tri 15183 5161 15190 5168 se
rect 15190 5161 15243 5168
tri 14938 5136 14963 5161 se
rect 14963 5136 15012 5161
tri 15012 5136 15037 5161 nw
tri 15158 5136 15183 5161 se
rect 15183 5147 15243 5161
rect 15183 5136 15226 5147
tri 14932 5130 14938 5136 se
rect 14938 5130 15006 5136
tri 15006 5130 15012 5136 nw
tri 15152 5130 15158 5136 se
rect 15158 5130 15226 5136
tri 15226 5130 15243 5147 nw
tri 14929 5127 14932 5130 se
rect 14932 5127 15003 5130
tri 15003 5127 15006 5130 nw
tri 15149 5127 15152 5130 se
rect 15152 5127 15192 5130
rect 11612 5075 11619 5127
rect 11671 5075 11683 5127
rect 11735 5075 11742 5127
rect 14353 5075 14359 5127
rect 14411 5075 14423 5127
rect 14475 5125 14483 5127
rect 14484 5126 14510 5127
rect 14511 5125 14972 5127
rect 14475 5118 14972 5125
rect 14475 5084 14526 5118
rect 14560 5084 14598 5118
rect 14632 5096 14972 5118
tri 14972 5096 15003 5127 nw
tri 15118 5096 15149 5127 se
rect 15149 5096 15192 5127
tri 15192 5096 15226 5130 nw
rect 14632 5095 14971 5096
tri 14971 5095 14972 5096 nw
tri 15117 5095 15118 5096 se
rect 15118 5095 15191 5096
tri 15191 5095 15192 5096 nw
rect 14632 5084 14951 5095
rect 14475 5077 14951 5084
rect 14475 5075 14483 5077
rect 14484 5075 14510 5076
rect 14511 5075 14951 5077
tri 14951 5075 14971 5095 nw
tri 15097 5075 15117 5095 se
rect 15117 5075 15154 5095
rect 11612 4973 11742 5075
tri 15080 5058 15097 5075 se
rect 15097 5058 15154 5075
tri 15154 5058 15191 5095 nw
tri 15051 5029 15080 5058 se
rect 15080 5029 15125 5058
tri 15125 5029 15154 5058 nw
tri 15046 5024 15051 5029 se
rect 15051 5024 15120 5029
tri 15120 5024 15125 5029 nw
tri 15266 5024 15271 5029 se
rect 15271 5024 15323 6952
tri 15043 5021 15046 5024 se
rect 15046 5021 15117 5024
tri 15117 5021 15120 5024 nw
tri 15263 5021 15266 5024 se
rect 15266 5021 15323 5024
tri 15008 4986 15043 5021 se
rect 15043 4986 15082 5021
tri 15082 4986 15117 5021 nw
tri 15228 4986 15263 5021 se
rect 15263 5007 15323 5021
rect 15263 4986 15302 5007
tri 15302 4986 15323 5007 nw
tri 14995 4973 15008 4986 se
rect 15008 4973 15069 4986
tri 15069 4973 15082 4986 nw
tri 15215 4973 15228 4986 se
rect 15228 4973 15271 4986
rect 11612 4921 11619 4973
rect 11671 4921 11683 4973
rect 11735 4921 11742 4973
rect 14349 4921 14355 4973
rect 14407 4921 14419 4973
rect 14471 4921 14479 4973
rect 14480 4922 14481 4972
rect 14509 4922 14510 4972
rect 14511 4964 15051 4973
rect 14511 4930 14526 4964
rect 14560 4930 14598 4964
rect 14632 4955 15051 4964
tri 15051 4955 15069 4973 nw
tri 15197 4955 15215 4973 se
rect 15215 4955 15271 4973
tri 15271 4955 15302 4986 nw
rect 14632 4952 15048 4955
tri 15048 4952 15051 4955 nw
tri 15194 4952 15197 4955 se
rect 15197 4952 15268 4955
tri 15268 4952 15271 4955 nw
rect 14632 4930 15017 4952
rect 14511 4921 15017 4930
tri 15017 4921 15048 4952 nw
tri 15163 4921 15194 4952 se
rect 15194 4921 15230 4952
rect 11612 4886 11742 4921
tri 15156 4914 15163 4921 se
rect 15163 4914 15230 4921
tri 15230 4914 15268 4952 nw
tri 15154 4912 15156 4914 se
rect 15156 4912 15205 4914
tri 15131 4889 15154 4912 se
rect 15154 4889 15205 4912
tri 15205 4889 15230 4914 nw
tri 15128 4886 15131 4889 se
rect 15131 4886 15197 4889
tri 15127 4885 15128 4886 se
rect 15128 4885 15197 4886
rect 11613 4884 11741 4885
tri 15126 4884 15127 4885 se
rect 15127 4884 15197 4885
tri 15123 4881 15126 4884 se
rect 15126 4881 15197 4884
tri 15197 4881 15205 4889 nw
tri 15343 4881 15351 4889 se
rect 15351 4881 15403 7074
tri 15122 4880 15123 4881 se
rect 15123 4880 15196 4881
tri 15196 4880 15197 4881 nw
tri 15342 4880 15343 4881 se
rect 15343 4880 15403 4881
rect 11494 4825 11500 4859
rect 11534 4825 11540 4859
tri 15098 4856 15122 4880 se
rect 15122 4856 15158 4880
rect 11494 4786 11540 4825
rect 11494 4752 11500 4786
rect 11534 4752 11540 4786
rect 11494 4713 11540 4752
rect 11494 4679 11500 4713
rect 11534 4679 11540 4713
rect 11494 4640 11540 4679
rect 11494 4606 11500 4640
rect 11534 4606 11540 4640
rect 11494 4567 11540 4606
rect 11613 4855 11741 4856
tri 15097 4855 15098 4856 se
rect 15098 4855 15158 4856
tri 15096 4854 15097 4855 se
rect 15097 4854 15158 4855
rect 11612 4819 11742 4854
tri 15084 4842 15096 4854 se
rect 15096 4842 15158 4854
tri 15158 4842 15196 4880 nw
tri 15304 4842 15342 4880 se
rect 15342 4867 15403 4880
rect 15342 4842 15378 4867
tri 15378 4842 15403 4867 nw
tri 15070 4828 15084 4842 se
rect 15084 4828 15144 4842
tri 15144 4828 15158 4842 nw
tri 15290 4828 15304 4842 se
rect 15304 4828 15351 4842
tri 15061 4819 15070 4828 se
rect 15070 4819 15135 4828
tri 15135 4819 15144 4828 nw
tri 15281 4819 15290 4828 se
rect 15290 4819 15351 4828
rect 11612 4767 11619 4819
rect 11671 4767 11683 4819
rect 11735 4767 11742 4819
rect 14353 4767 14359 4819
rect 14411 4767 14423 4819
rect 14475 4817 14483 4819
rect 14484 4818 14510 4819
rect 14511 4817 15131 4819
rect 14475 4815 15131 4817
tri 15131 4815 15135 4819 nw
tri 15277 4815 15281 4819 se
rect 15281 4815 15351 4819
tri 15351 4815 15378 4842 nw
rect 14475 4810 15124 4815
rect 14475 4776 14526 4810
rect 14560 4776 14598 4810
rect 14632 4808 15124 4810
tri 15124 4808 15131 4815 nw
tri 15270 4808 15277 4815 se
rect 15277 4808 15344 4815
tri 15344 4808 15351 4815 nw
rect 14632 4776 15086 4808
rect 14475 4770 15086 4776
tri 15086 4770 15124 4808 nw
tri 15232 4770 15270 4808 se
rect 15270 4770 15306 4808
tri 15306 4770 15344 4808 nw
rect 14475 4769 15083 4770
rect 14475 4767 14483 4769
rect 14484 4767 14510 4768
rect 14511 4767 15083 4769
tri 15083 4767 15086 4770 nw
tri 15229 4767 15232 4770 se
rect 15232 4767 15277 4770
rect 11612 4665 11742 4767
tri 15203 4741 15229 4767 se
rect 15229 4741 15277 4767
tri 15277 4741 15306 4770 nw
tri 15423 4741 15431 4749 se
rect 15431 4741 15483 7214
tri 15198 4736 15203 4741 se
rect 15203 4736 15272 4741
tri 15272 4736 15277 4741 nw
tri 15418 4736 15423 4741 se
rect 15423 4736 15483 4741
tri 15160 4698 15198 4736 se
rect 15198 4698 15234 4736
tri 15234 4698 15272 4736 nw
tri 15395 4713 15418 4736 se
rect 15418 4727 15483 4736
rect 15418 4713 15469 4727
tri 15469 4713 15483 4727 nw
tri 15380 4698 15395 4713 se
rect 15395 4698 15454 4713
tri 15454 4698 15469 4713 nw
tri 15496 4698 15511 4713 se
rect 15511 4698 15563 7354
tri 15129 4667 15160 4698 se
rect 15160 4667 15203 4698
tri 15203 4667 15234 4698 nw
tri 15357 4675 15380 4698 se
rect 15380 4685 15441 4698
tri 15441 4685 15454 4698 nw
tri 15483 4685 15496 4698 se
rect 15496 4691 15563 4698
rect 15496 4685 15536 4691
rect 15380 4675 15431 4685
tri 15431 4675 15441 4685 nw
tri 15473 4675 15483 4685 se
rect 15483 4675 15536 4685
tri 15349 4667 15357 4675 se
rect 15357 4667 15423 4675
tri 15423 4667 15431 4675 nw
tri 15465 4667 15473 4675 se
rect 15473 4667 15536 4675
tri 15127 4665 15129 4667 se
rect 15129 4665 15201 4667
tri 15201 4665 15203 4667 nw
tri 15347 4665 15349 4667 se
rect 15349 4665 15421 4667
tri 15421 4665 15423 4667 nw
tri 15463 4665 15465 4667 se
rect 15465 4665 15536 4667
rect 11612 4613 11619 4665
rect 11671 4613 11683 4665
rect 11735 4613 11742 4665
rect 14349 4613 14355 4665
rect 14407 4613 14419 4665
rect 14471 4613 14479 4665
rect 14480 4614 14481 4664
rect 14511 4664 15200 4665
tri 15200 4664 15201 4665 nw
tri 15346 4664 15347 4665 se
rect 15347 4664 15420 4665
tri 15420 4664 15421 4665 nw
tri 15462 4664 15463 4665 se
rect 15463 4664 15536 4665
tri 15536 4664 15563 4691 nw
rect 14509 4614 14510 4664
rect 14511 4656 15162 4664
rect 14511 4622 14526 4656
rect 14560 4622 14598 4656
rect 14632 4626 15162 4656
tri 15162 4626 15200 4664 nw
tri 15321 4639 15346 4664 se
rect 15346 4639 15395 4664
tri 15395 4639 15420 4664 nw
tri 15437 4639 15462 4664 se
rect 15462 4639 15511 4664
tri 15511 4639 15536 4664 nw
tri 15308 4626 15321 4639 se
rect 15321 4633 15389 4639
tri 15389 4633 15395 4639 nw
tri 15431 4633 15437 4639 se
rect 15437 4633 15498 4639
rect 15321 4626 15382 4633
tri 15382 4626 15389 4633 nw
tri 15424 4626 15431 4633 se
rect 15431 4626 15498 4633
tri 15498 4626 15511 4639 nw
rect 14632 4622 15149 4626
rect 14511 4613 15149 4622
tri 15149 4613 15162 4626 nw
tri 15295 4613 15308 4626 se
rect 15308 4613 15369 4626
tri 15369 4613 15382 4626 nw
tri 15411 4613 15424 4626 se
rect 15424 4613 15464 4626
rect 11612 4578 11742 4613
tri 15286 4604 15295 4613 se
rect 15295 4604 15360 4613
tri 15360 4604 15369 4613 nw
tri 15402 4604 15411 4613 se
rect 15411 4604 15464 4613
tri 15283 4601 15286 4604 se
rect 15286 4601 15357 4604
tri 15357 4601 15360 4604 nw
tri 15399 4601 15402 4604 se
rect 15402 4601 15464 4604
tri 15274 4592 15283 4601 se
rect 15283 4592 15348 4601
tri 15348 4592 15357 4601 nw
tri 15390 4592 15399 4601 se
rect 15399 4592 15464 4601
tri 15464 4592 15498 4626 nw
tri 15582 4592 15591 4601 se
rect 15591 4592 15643 7494
tri 15260 4578 15274 4592 se
rect 15274 4578 15321 4592
tri 15259 4577 15260 4578 se
rect 15260 4577 15321 4578
rect 11613 4576 11741 4577
tri 15258 4576 15259 4577 se
rect 15259 4576 15321 4577
rect 11494 4533 11500 4567
rect 11534 4533 11540 4567
tri 15247 4565 15258 4576 se
rect 15258 4565 15321 4576
tri 15321 4565 15348 4592 nw
tri 15363 4565 15390 4592 se
rect 15390 4565 15437 4592
tri 15437 4565 15464 4592 nw
tri 15555 4565 15582 4592 se
rect 15582 4579 15643 4592
rect 15582 4565 15618 4579
tri 15236 4554 15247 4565 se
rect 15247 4559 15315 4565
tri 15315 4559 15321 4565 nw
tri 15357 4559 15363 4565 se
rect 15363 4559 15426 4565
rect 15247 4554 15310 4559
tri 15310 4554 15315 4559 nw
tri 15352 4554 15357 4559 se
rect 15357 4554 15426 4559
tri 15426 4554 15437 4565 nw
tri 15544 4554 15555 4565 se
rect 15555 4554 15618 4565
tri 15618 4554 15643 4579 nw
rect 15725 7472 15733 7506
rect 15767 7472 15819 7506
rect 15853 7472 15905 7506
rect 15939 7472 15991 7506
rect 16025 7472 16033 7506
rect 15725 7434 16033 7472
rect 15725 7400 15733 7434
rect 15767 7400 15819 7434
rect 15853 7400 15905 7434
rect 15939 7400 15991 7434
rect 16025 7400 16033 7434
rect 15725 7362 16033 7400
rect 15725 7328 15733 7362
rect 15767 7328 15819 7362
rect 15853 7328 15905 7362
rect 15939 7328 15991 7362
rect 16025 7328 16033 7362
rect 15725 7290 16033 7328
rect 15725 7256 15733 7290
rect 15767 7256 15819 7290
rect 15853 7256 15905 7290
rect 15939 7256 15991 7290
rect 16025 7256 16033 7290
rect 15725 7218 16033 7256
rect 15725 7184 15733 7218
rect 15767 7184 15819 7218
rect 15853 7184 15905 7218
rect 15939 7184 15991 7218
rect 16025 7184 16033 7218
rect 15725 7146 16033 7184
rect 15725 7112 15733 7146
rect 15767 7112 15819 7146
rect 15853 7112 15905 7146
rect 15939 7112 15991 7146
rect 16025 7112 16033 7146
rect 15725 7074 16033 7112
rect 15725 7040 15733 7074
rect 15767 7040 15819 7074
rect 15853 7040 15905 7074
rect 15939 7040 15991 7074
rect 16025 7040 16033 7074
rect 15725 7002 16033 7040
rect 15725 6968 15733 7002
rect 15767 6968 15819 7002
rect 15853 6968 15905 7002
rect 15939 6968 15991 7002
rect 16025 6968 16033 7002
rect 15725 6930 16033 6968
rect 15725 6896 15733 6930
rect 15767 6896 15819 6930
rect 15853 6896 15905 6930
rect 15939 6896 15991 6930
rect 16025 6896 16033 6930
rect 15725 6858 16033 6896
rect 15725 6824 15733 6858
rect 15767 6824 15819 6858
rect 15853 6824 15905 6858
rect 15939 6824 15991 6858
rect 16025 6824 16033 6858
rect 15725 6786 16033 6824
rect 15725 6752 15733 6786
rect 15767 6752 15819 6786
rect 15853 6752 15905 6786
rect 15939 6752 15991 6786
rect 16025 6752 16033 6786
rect 15725 6714 16033 6752
rect 15725 6680 15733 6714
rect 15767 6680 15819 6714
rect 15853 6680 15905 6714
rect 15939 6680 15991 6714
rect 16025 6680 16033 6714
rect 15725 6642 16033 6680
rect 15725 6608 15733 6642
rect 15767 6608 15819 6642
rect 15853 6608 15905 6642
rect 15939 6608 15991 6642
rect 16025 6608 16033 6642
rect 15725 6570 16033 6608
rect 15725 6536 15733 6570
rect 15767 6536 15819 6570
rect 15853 6536 15905 6570
rect 15939 6536 15991 6570
rect 16025 6536 16033 6570
rect 15725 6498 16033 6536
rect 15725 6464 15733 6498
rect 15767 6464 15819 6498
rect 15853 6464 15905 6498
rect 15939 6464 15991 6498
rect 16025 6464 16033 6498
rect 15725 6426 16033 6464
rect 15725 6392 15733 6426
rect 15767 6392 15819 6426
rect 15853 6392 15905 6426
rect 15939 6392 15991 6426
rect 16025 6392 16033 6426
rect 15725 6354 16033 6392
rect 15725 6320 15733 6354
rect 15767 6320 15819 6354
rect 15853 6320 15905 6354
rect 15939 6320 15991 6354
rect 16025 6320 16033 6354
rect 15725 6282 16033 6320
rect 15725 6248 15733 6282
rect 15767 6248 15819 6282
rect 15853 6248 15905 6282
rect 15939 6248 15991 6282
rect 16025 6248 16033 6282
rect 15725 6210 16033 6248
rect 15725 6176 15733 6210
rect 15767 6176 15819 6210
rect 15853 6176 15905 6210
rect 15939 6176 15991 6210
rect 16025 6176 16033 6210
rect 15725 6138 16033 6176
rect 15725 6104 15733 6138
rect 15767 6104 15819 6138
rect 15853 6104 15905 6138
rect 15939 6104 15991 6138
rect 16025 6104 16033 6138
rect 15725 6066 16033 6104
rect 15725 6032 15733 6066
rect 15767 6032 15819 6066
rect 15853 6032 15905 6066
rect 15939 6032 15991 6066
rect 16025 6032 16033 6066
rect 15725 5994 16033 6032
rect 15725 5960 15733 5994
rect 15767 5960 15819 5994
rect 15853 5960 15905 5994
rect 15939 5960 15991 5994
rect 16025 5960 16033 5994
rect 15725 5922 16033 5960
rect 15725 5888 15733 5922
rect 15767 5888 15819 5922
rect 15853 5888 15905 5922
rect 15939 5888 15991 5922
rect 16025 5888 16033 5922
rect 15725 5850 16033 5888
rect 15725 5816 15733 5850
rect 15767 5816 15819 5850
rect 15853 5816 15905 5850
rect 15939 5816 15991 5850
rect 16025 5816 16033 5850
rect 15725 5778 16033 5816
rect 15725 5744 15733 5778
rect 15767 5744 15819 5778
rect 15853 5744 15905 5778
rect 15939 5744 15991 5778
rect 16025 5744 16033 5778
rect 15725 5706 16033 5744
rect 15725 5672 15733 5706
rect 15767 5672 15819 5706
rect 15853 5672 15905 5706
rect 15939 5672 15991 5706
rect 16025 5672 16033 5706
rect 15725 5634 16033 5672
rect 15725 5600 15733 5634
rect 15767 5600 15819 5634
rect 15853 5600 15905 5634
rect 15939 5600 15991 5634
rect 16025 5600 16033 5634
rect 15725 5562 16033 5600
rect 15725 5528 15733 5562
rect 15767 5528 15819 5562
rect 15853 5528 15905 5562
rect 15939 5528 15991 5562
rect 16025 5528 16033 5562
rect 15725 5490 16033 5528
rect 15725 5456 15733 5490
rect 15767 5456 15819 5490
rect 15853 5456 15905 5490
rect 15939 5456 15991 5490
rect 16025 5456 16033 5490
rect 15725 5418 16033 5456
rect 15725 5384 15733 5418
rect 15767 5384 15819 5418
rect 15853 5384 15905 5418
rect 15939 5384 15991 5418
rect 16025 5384 16033 5418
rect 15725 5346 16033 5384
rect 15725 5312 15733 5346
rect 15767 5312 15819 5346
rect 15853 5312 15905 5346
rect 15939 5312 15991 5346
rect 16025 5312 16033 5346
rect 15725 5274 16033 5312
rect 15725 5240 15733 5274
rect 15767 5240 15819 5274
rect 15853 5240 15905 5274
rect 15939 5240 15991 5274
rect 16025 5240 16033 5274
rect 15725 5202 16033 5240
rect 15725 5168 15733 5202
rect 15767 5168 15819 5202
rect 15853 5168 15905 5202
rect 15939 5168 15991 5202
rect 16025 5168 16033 5202
rect 15725 5130 16033 5168
rect 15725 5096 15733 5130
rect 15767 5096 15819 5130
rect 15853 5096 15905 5130
rect 15939 5096 15991 5130
rect 16025 5096 16033 5130
rect 15725 5058 16033 5096
rect 15725 5024 15733 5058
rect 15767 5024 15819 5058
rect 15853 5024 15905 5058
rect 15939 5024 15991 5058
rect 16025 5024 16033 5058
rect 15725 4986 16033 5024
rect 15725 4952 15733 4986
rect 15767 4952 15819 4986
rect 15853 4952 15905 4986
rect 15939 4952 15991 4986
rect 16025 4952 16033 4986
rect 15725 4914 16033 4952
rect 15725 4880 15733 4914
rect 15767 4880 15819 4914
rect 15853 4880 15905 4914
rect 15939 4880 15991 4914
rect 16025 4880 16033 4914
rect 15725 4842 16033 4880
rect 15725 4808 15733 4842
rect 15767 4808 15819 4842
rect 15853 4808 15905 4842
rect 15939 4808 15991 4842
rect 16025 4808 16033 4842
rect 15725 4770 16033 4808
rect 15725 4736 15733 4770
rect 15767 4736 15819 4770
rect 15853 4736 15905 4770
rect 15939 4736 15991 4770
rect 16025 4736 16033 4770
rect 15725 4698 16033 4736
rect 15725 4664 15733 4698
rect 15767 4664 15819 4698
rect 15853 4664 15905 4698
rect 15939 4664 15991 4698
rect 16025 4664 16033 4698
rect 15725 4626 16033 4664
rect 15725 4592 15733 4626
rect 15767 4592 15819 4626
rect 15853 4592 15905 4626
rect 15939 4592 15991 4626
rect 16025 4592 16033 4626
rect 15725 4554 16033 4592
tri 15230 4548 15236 4554 se
rect 15236 4548 15283 4554
rect 11494 4494 11540 4533
rect 11494 4460 11500 4494
rect 11534 4460 11540 4494
rect 11494 4421 11540 4460
rect 11494 4387 11500 4421
rect 11534 4387 11540 4421
rect 11494 4348 11540 4387
rect 11494 4314 11500 4348
rect 11534 4314 11540 4348
rect 11494 4275 11540 4314
rect 11613 4547 11741 4548
tri 15229 4547 15230 4548 se
rect 15230 4547 15283 4548
tri 15228 4546 15229 4547 se
rect 15229 4546 15283 4547
rect 11612 4511 11742 4546
tri 15209 4527 15228 4546 se
rect 15228 4527 15283 4546
tri 15283 4527 15310 4554 nw
tri 15325 4527 15352 4554 se
rect 15352 4527 15392 4554
tri 15202 4520 15209 4527 se
rect 15209 4520 15276 4527
tri 15276 4520 15283 4527 nw
tri 15318 4520 15325 4527 se
rect 15325 4520 15392 4527
tri 15392 4520 15426 4554 nw
tri 15517 4527 15544 4554 se
rect 15544 4527 15591 4554
tri 15591 4527 15618 4554 nw
tri 15510 4520 15517 4527 se
rect 15517 4520 15584 4527
tri 15584 4520 15591 4527 nw
rect 15725 4520 15733 4554
rect 15767 4520 15819 4554
rect 15853 4520 15905 4554
rect 15939 4520 15991 4554
rect 16025 4520 16033 4554
tri 15193 4511 15202 4520 se
rect 15202 4511 15267 4520
tri 15267 4511 15276 4520 nw
tri 15309 4511 15318 4520 se
rect 15318 4511 15363 4520
rect 11612 4459 11619 4511
rect 11671 4459 11683 4511
rect 11735 4459 11742 4511
rect 14353 4459 14359 4511
rect 14411 4459 14423 4511
rect 14475 4509 14483 4511
rect 14484 4510 14510 4511
rect 14511 4509 15247 4511
rect 14475 4502 15247 4509
rect 14475 4468 14526 4502
rect 14560 4468 14598 4502
rect 14632 4491 15247 4502
tri 15247 4491 15267 4511 nw
tri 15289 4491 15309 4511 se
rect 15309 4491 15363 4511
tri 15363 4491 15392 4520 nw
tri 15481 4491 15510 4520 se
rect 15510 4491 15546 4520
rect 14632 4485 15241 4491
tri 15241 4485 15247 4491 nw
tri 15283 4485 15289 4491 se
rect 15289 4485 15354 4491
rect 14632 4482 15238 4485
tri 15238 4482 15241 4485 nw
tri 15280 4482 15283 4485 se
rect 15283 4482 15354 4485
tri 15354 4482 15363 4491 nw
tri 15472 4482 15481 4491 se
rect 15481 4482 15546 4491
tri 15546 4482 15584 4520 nw
rect 15725 4482 16033 4520
rect 14632 4468 15215 4482
rect 14475 4461 15215 4468
rect 14475 4459 14483 4461
rect 14484 4459 14510 4460
rect 14511 4459 15215 4461
tri 15215 4459 15238 4482 nw
tri 15257 4459 15280 4482 se
rect 15280 4459 15320 4482
rect 11612 4357 11742 4459
tri 15246 4448 15257 4459 se
rect 15257 4448 15320 4459
tri 15320 4448 15354 4482 nw
tri 15443 4453 15472 4482 se
rect 15472 4453 15517 4482
tri 15517 4453 15546 4482 nw
tri 15438 4448 15443 4453 se
rect 15443 4448 15512 4453
tri 15512 4448 15517 4453 nw
rect 15725 4448 15733 4482
rect 15767 4448 15819 4482
rect 15853 4448 15905 4482
rect 15939 4448 15991 4482
rect 16025 4448 16033 4482
tri 15215 4417 15246 4448 se
rect 15246 4435 15307 4448
tri 15307 4435 15320 4448 nw
tri 15425 4435 15438 4448 se
rect 15438 4435 15499 4448
tri 15499 4435 15512 4448 nw
rect 15246 4417 15289 4435
tri 15289 4417 15307 4435 nw
tri 15407 4417 15425 4435 se
rect 15425 4417 15474 4435
tri 15208 4410 15215 4417 se
rect 15215 4410 15282 4417
tri 15282 4410 15289 4417 nw
tri 15400 4410 15407 4417 se
rect 15407 4410 15474 4417
tri 15474 4410 15499 4435 nw
tri 15700 4410 15725 4435 se
rect 15725 4410 16033 4448
tri 15174 4376 15208 4410 se
rect 15208 4376 15248 4410
tri 15248 4376 15282 4410 nw
tri 15369 4379 15400 4410 se
rect 15400 4379 15443 4410
tri 15443 4379 15474 4410 nw
tri 15669 4379 15700 4410 se
rect 15700 4379 15733 4410
tri 15366 4376 15369 4379 se
rect 15369 4376 15440 4379
tri 15440 4376 15443 4379 nw
tri 15666 4376 15669 4379 se
rect 15669 4376 15733 4379
rect 15767 4376 15819 4410
rect 15853 4376 15905 4410
rect 15939 4376 15991 4410
rect 16025 4376 16033 4410
tri 15155 4357 15174 4376 se
rect 15174 4357 15229 4376
tri 15229 4357 15248 4376 nw
tri 15347 4357 15366 4376 se
rect 15366 4357 15402 4376
rect 11612 4305 11619 4357
rect 11671 4305 11683 4357
rect 11735 4305 11742 4357
rect 14349 4305 14355 4357
rect 14407 4305 14419 4357
rect 14471 4305 14479 4357
rect 14480 4306 14481 4356
rect 14509 4306 14510 4356
rect 14511 4348 15210 4357
rect 14511 4314 14526 4348
rect 14560 4314 14598 4348
rect 14632 4338 15210 4348
tri 15210 4338 15229 4357 nw
tri 15328 4338 15347 4357 se
rect 15347 4338 15402 4357
tri 15402 4338 15440 4376 nw
tri 15628 4338 15666 4376 se
rect 15666 4338 16033 4376
rect 14632 4314 15177 4338
rect 14511 4305 15177 4314
tri 15177 4305 15210 4338 nw
tri 15324 4334 15328 4338 se
rect 15328 4334 15369 4338
tri 15295 4305 15324 4334 se
rect 15324 4305 15369 4334
tri 15369 4305 15402 4338 nw
tri 15595 4305 15628 4338 se
rect 15628 4305 15733 4338
tri 15294 4304 15295 4305 se
rect 15295 4304 15368 4305
tri 15368 4304 15369 4305 nw
tri 15594 4304 15595 4305 se
rect 15595 4304 15733 4305
rect 15767 4304 15819 4338
rect 15853 4304 15905 4338
rect 15939 4304 15991 4338
rect 16025 4304 16033 4338
rect 11494 4241 11500 4275
rect 11534 4241 11540 4275
tri 15256 4266 15294 4304 se
rect 15294 4266 15330 4304
tri 15330 4266 15368 4304 nw
tri 15556 4266 15594 4304 se
rect 15594 4266 16033 4304
tri 15236 4246 15256 4266 se
rect 15256 4260 15324 4266
tri 15324 4260 15330 4266 nw
tri 15550 4260 15556 4266 se
rect 15556 4260 15733 4266
rect 15256 4246 15310 4260
tri 15310 4246 15324 4260 nw
tri 15542 4252 15550 4260 se
rect 15550 4252 15733 4260
tri 15536 4246 15542 4252 se
rect 15542 4246 15733 4252
rect 11494 4202 11540 4241
tri 15221 4231 15236 4246 se
rect 15236 4231 15295 4246
tri 15295 4231 15310 4246 nw
tri 15521 4231 15536 4246 se
rect 15536 4231 15554 4246
tri 15202 4212 15221 4231 se
rect 15221 4212 15276 4231
tri 15276 4212 15295 4231 nw
tri 15502 4212 15521 4231 se
rect 15521 4212 15554 4231
rect 15588 4212 15626 4246
rect 15660 4232 15733 4246
rect 15767 4232 15819 4266
rect 15853 4232 15905 4266
rect 15939 4232 15991 4266
rect 16025 4232 16033 4266
rect 15660 4212 16033 4232
tri 15193 4203 15202 4212 se
rect 15202 4203 15267 4212
tri 15267 4203 15276 4212 nw
tri 15493 4203 15502 4212 se
rect 15502 4203 16033 4212
rect 11494 4168 11500 4202
rect 11534 4168 11540 4202
rect 11494 4129 11540 4168
rect 11612 4151 11619 4203
rect 11671 4151 11683 4203
rect 11735 4151 11742 4203
rect 14353 4151 14359 4203
rect 14411 4151 14423 4203
rect 14475 4201 14483 4203
rect 14484 4202 14510 4203
rect 14511 4201 15258 4203
rect 14475 4194 15258 4201
tri 15258 4194 15267 4203 nw
tri 15484 4194 15493 4203 se
rect 15493 4194 16033 4203
rect 14475 4160 14526 4194
rect 14560 4160 14598 4194
rect 14632 4173 15237 4194
tri 15237 4173 15258 4194 nw
tri 15475 4185 15484 4194 se
rect 15484 4185 15733 4194
tri 15463 4173 15475 4185 se
rect 15475 4173 15733 4185
rect 14632 4160 15215 4173
rect 14475 4153 15215 4160
rect 14475 4151 14483 4153
rect 14484 4151 14510 4152
rect 14511 4151 15215 4153
tri 15215 4151 15237 4173 nw
tri 15441 4151 15463 4173 se
rect 15463 4151 15484 4173
tri 15429 4139 15441 4151 se
rect 15441 4139 15484 4151
rect 15518 4139 15560 4173
rect 15594 4139 15636 4173
rect 15670 4160 15733 4173
rect 15767 4160 15819 4194
rect 15853 4160 15905 4194
rect 15939 4160 15991 4194
rect 16025 4160 16033 4194
rect 15670 4139 16033 4160
rect 11494 4095 11500 4129
rect 11534 4100 11540 4129
tri 15412 4122 15429 4139 se
rect 15429 4122 16033 4139
tri 15399 4109 15412 4122 se
rect 15412 4109 15733 4122
tri 11540 4100 11549 4109 sw
tri 15390 4100 15399 4109 se
rect 15399 4100 15733 4109
rect 11534 4095 11549 4100
rect 11494 4092 11549 4095
tri 11549 4092 11557 4100 sw
tri 15382 4092 15390 4100 se
rect 15390 4092 15733 4100
rect 11494 4088 11557 4092
tri 11557 4088 11561 4092 sw
tri 15378 4088 15382 4092 se
rect 15382 4088 15484 4092
rect 11494 4057 11561 4088
tri 11561 4057 11592 4088 sw
tri 15347 4057 15378 4088 se
rect 15378 4057 15405 4088
rect 11494 4056 15405 4057
rect 11494 4022 11500 4056
rect 11534 4054 15405 4056
rect 15439 4058 15484 4088
rect 15518 4058 15560 4092
rect 15594 4058 15636 4092
rect 15670 4088 15733 4092
rect 15767 4088 15819 4122
rect 15853 4088 15905 4122
rect 15939 4088 15991 4122
rect 16025 4088 16033 4122
rect 15670 4058 16033 4088
rect 15439 4054 16033 4058
rect 11534 4051 16033 4054
rect 11534 4022 11583 4051
rect 11494 4017 11583 4022
rect 11617 4017 11656 4051
rect 11690 4017 11729 4051
rect 11763 4017 11801 4051
rect 11835 4017 11873 4051
rect 11907 4017 11945 4051
rect 11979 4017 12017 4051
rect 12051 4017 12089 4051
rect 12123 4017 12161 4051
rect 12195 4017 12233 4051
rect 12267 4017 12305 4051
rect 12339 4017 12377 4051
rect 12411 4017 12449 4051
rect 12483 4017 12521 4051
rect 12555 4017 12593 4051
rect 12627 4017 12665 4051
rect 12699 4017 12737 4051
rect 12771 4017 12809 4051
rect 12843 4017 12881 4051
rect 12915 4017 12953 4051
rect 12987 4017 13025 4051
rect 13059 4017 13097 4051
rect 13131 4017 13169 4051
rect 13203 4017 13241 4051
rect 13275 4017 13313 4051
rect 13347 4017 13385 4051
rect 13419 4017 13457 4051
rect 13491 4017 13529 4051
rect 13563 4017 13601 4051
rect 13635 4017 13673 4051
rect 13707 4017 13745 4051
rect 13779 4017 13817 4051
rect 13851 4017 13889 4051
rect 13923 4017 13961 4051
rect 13995 4017 14033 4051
rect 14067 4017 14105 4051
rect 14139 4017 14177 4051
rect 14211 4017 14249 4051
rect 14283 4017 14321 4051
rect 14355 4017 14393 4051
rect 14427 4017 14465 4051
rect 14499 4017 14537 4051
rect 14571 4017 14609 4051
rect 14643 4017 14681 4051
rect 14715 4017 14753 4051
rect 14787 4017 14825 4051
rect 14859 4017 14897 4051
rect 14931 4017 14969 4051
rect 15003 4017 15041 4051
rect 15075 4017 15113 4051
rect 15147 4017 15185 4051
rect 15219 4017 15257 4051
rect 15291 4017 15329 4051
rect 15363 4050 16033 4051
rect 15363 4017 15733 4050
rect 11494 4016 15733 4017
rect 15767 4016 15819 4050
rect 15853 4016 15905 4050
rect 15939 4016 15991 4050
rect 16025 4016 16033 4050
rect 11494 4011 15405 4016
rect 11494 4010 11577 4011
tri 11577 4010 11578 4011 nw
tri 15347 4010 15348 4011 ne
rect 15348 4010 15405 4011
rect 11494 3950 11552 4010
tri 11552 3985 11577 4010 nw
tri 15348 3985 15373 4010 ne
rect 15373 3985 15405 4010
tri 15373 3982 15376 3985 ne
rect 15376 3982 15405 3985
rect 15439 4012 16033 4016
rect 15439 3982 15484 4012
tri 15376 3978 15380 3982 ne
rect 15380 3978 15484 3982
rect 15518 3978 15560 4012
rect 15594 3978 15636 4012
rect 15670 3978 16033 4012
tri 15380 3970 15388 3978 ne
rect 15388 3970 15733 3978
rect 11494 3916 11506 3950
rect 11540 3916 11552 3950
tri 15388 3944 15414 3970 ne
rect 15414 3944 15733 3970
rect 15767 3944 15819 3978
rect 15853 3944 15905 3978
rect 15939 3944 15991 3978
rect 16025 3944 16033 3978
tri 15414 3932 15426 3944 ne
rect 15426 3932 16033 3944
tri 15426 3917 15441 3932 ne
rect 15441 3917 15484 3932
rect 11494 3878 11552 3916
rect 11494 3844 11506 3878
rect 11540 3844 11552 3878
rect 11494 3806 11552 3844
rect 11494 3772 11506 3806
rect 11540 3772 11552 3806
rect 11494 3734 11552 3772
rect 11494 3700 11506 3734
rect 11540 3700 11552 3734
rect 11612 3865 11619 3917
rect 11671 3865 11683 3917
rect 11735 3865 11742 3917
rect 14353 3865 14359 3917
rect 14411 3865 14423 3917
rect 14475 3915 14483 3917
rect 14484 3916 14510 3917
rect 14511 3915 15173 3917
rect 14475 3908 15173 3915
rect 14475 3874 14526 3908
rect 14560 3874 14598 3908
rect 14632 3874 15173 3908
rect 14475 3867 15173 3874
rect 14475 3865 14483 3867
rect 14484 3865 14510 3866
rect 14511 3865 15173 3867
rect 15225 3865 15237 3917
rect 15289 3865 15295 3917
tri 15441 3898 15460 3917 ne
rect 15460 3898 15484 3917
rect 15518 3898 15560 3932
rect 15594 3898 15636 3932
rect 15670 3906 16033 3932
rect 15670 3898 15733 3906
tri 15460 3886 15472 3898 ne
rect 15472 3886 15733 3898
tri 15472 3872 15486 3886 ne
rect 15486 3872 15733 3886
rect 15767 3872 15819 3906
rect 15853 3872 15905 3906
rect 15939 3872 15991 3906
rect 16025 3872 16033 3906
tri 15486 3865 15493 3872 ne
rect 15493 3865 16033 3872
rect 11612 3763 11742 3865
tri 15493 3859 15499 3865 ne
rect 15499 3859 16033 3865
tri 15499 3825 15533 3859 ne
rect 15533 3825 15554 3859
rect 15588 3825 15626 3859
rect 15660 3834 16033 3859
rect 15660 3825 15733 3834
tri 15533 3819 15539 3825 ne
rect 15539 3819 15733 3825
tri 15539 3800 15558 3819 ne
rect 15558 3800 15733 3819
rect 15767 3800 15819 3834
rect 15853 3800 15905 3834
rect 15939 3800 15991 3834
rect 16025 3800 16033 3834
tri 15558 3763 15595 3800 ne
rect 15595 3763 16033 3800
rect 11612 3711 11619 3763
rect 11671 3711 11683 3763
rect 11735 3711 11742 3763
rect 14349 3711 14355 3763
rect 14407 3711 14419 3763
rect 14471 3711 14479 3763
rect 14480 3712 14481 3762
rect 14509 3712 14510 3762
rect 14511 3754 15005 3763
rect 14511 3720 14526 3754
rect 14560 3720 14598 3754
rect 14632 3720 15005 3754
rect 14511 3711 15005 3720
rect 15057 3711 15069 3763
rect 15121 3711 15127 3763
tri 15595 3762 15596 3763 ne
rect 15596 3762 16033 3763
tri 15596 3728 15630 3762 ne
rect 15630 3728 15733 3762
rect 15767 3728 15819 3762
rect 15853 3728 15905 3762
rect 15939 3728 15991 3762
rect 16025 3728 16033 3762
tri 15630 3711 15647 3728 ne
rect 15647 3711 16033 3728
rect 11494 3662 11552 3700
tri 15647 3690 15668 3711 ne
rect 15668 3690 16033 3711
rect 11494 3628 11506 3662
rect 11540 3628 11552 3662
tri 15668 3656 15702 3690 ne
rect 15702 3656 15733 3690
rect 15767 3656 15819 3690
rect 15853 3656 15905 3690
rect 15939 3656 15991 3690
rect 16025 3656 16033 3690
tri 15702 3633 15725 3656 ne
rect 11494 3590 11552 3628
rect 15725 3618 16033 3656
rect 11494 3556 11506 3590
rect 11540 3556 11552 3590
rect 11494 3518 11552 3556
rect 11494 3484 11506 3518
rect 11540 3484 11552 3518
rect 11494 3446 11552 3484
rect 11494 3412 11506 3446
rect 11540 3412 11552 3446
rect 11494 3374 11552 3412
rect 11612 3557 11619 3609
rect 11671 3557 11683 3609
rect 11735 3557 11742 3609
rect 14353 3557 14359 3609
rect 14411 3557 14423 3609
rect 14475 3607 14483 3609
rect 14484 3608 14510 3609
rect 14511 3607 15467 3609
rect 14475 3600 15467 3607
rect 14475 3566 14526 3600
rect 14560 3566 14598 3600
rect 14632 3584 15467 3600
tri 15467 3584 15492 3609 sw
rect 15725 3584 15733 3618
rect 15767 3584 15819 3618
rect 15853 3584 15905 3618
rect 15939 3584 15991 3618
rect 16025 3584 16033 3618
rect 14632 3581 15492 3584
tri 15492 3581 15495 3584 sw
rect 14632 3566 15495 3581
rect 14475 3559 15495 3566
rect 14475 3557 14483 3559
rect 14484 3557 14510 3558
rect 14511 3557 15495 3559
tri 15495 3557 15519 3581 sw
rect 11612 3455 11742 3557
tri 15445 3546 15456 3557 ne
rect 15456 3546 15519 3557
tri 15519 3546 15530 3557 sw
rect 15725 3546 16033 3584
tri 15456 3512 15490 3546 ne
rect 15490 3512 15530 3546
tri 15530 3512 15564 3546 sw
rect 15725 3512 15733 3546
rect 15767 3512 15819 3546
rect 15853 3512 15905 3546
rect 15939 3512 15991 3546
rect 16025 3512 16033 3546
tri 15490 3507 15495 3512 ne
rect 15495 3507 15564 3512
tri 15564 3507 15569 3512 sw
tri 15495 3474 15528 3507 ne
rect 15528 3474 15569 3507
tri 15569 3474 15602 3507 sw
rect 15725 3474 16033 3512
tri 15528 3455 15547 3474 ne
rect 15547 3455 15602 3474
tri 15602 3455 15621 3474 sw
rect 11612 3403 11619 3455
rect 11671 3403 11683 3455
rect 11735 3403 11742 3455
rect 14349 3403 14355 3455
rect 14407 3403 14419 3455
rect 14471 3403 14479 3455
rect 14480 3404 14481 3454
rect 14509 3404 14510 3454
rect 14511 3446 15401 3455
rect 14511 3412 14526 3446
rect 14560 3412 14598 3446
rect 14632 3441 15401 3446
tri 15401 3441 15415 3455 sw
tri 15547 3441 15561 3455 ne
rect 15561 3441 15621 3455
tri 15621 3441 15635 3455 sw
rect 14632 3440 15415 3441
tri 15415 3440 15416 3441 sw
tri 15561 3440 15562 3441 ne
rect 15562 3440 15635 3441
tri 15635 3440 15636 3441 sw
rect 15725 3440 15733 3474
rect 15767 3440 15819 3474
rect 15853 3440 15905 3474
rect 15939 3440 15991 3474
rect 16025 3440 16033 3474
rect 14632 3412 15416 3440
rect 14511 3403 15416 3412
tri 15416 3403 15453 3440 sw
tri 15562 3433 15569 3440 ne
rect 15569 3433 15636 3440
tri 15636 3433 15643 3440 sw
tri 15569 3411 15591 3433 ne
tri 15379 3402 15380 3403 ne
rect 15380 3402 15453 3403
tri 15453 3402 15454 3403 sw
rect 11494 3340 11506 3374
rect 11540 3340 11552 3374
tri 15380 3368 15414 3402 ne
rect 15414 3368 15454 3402
tri 15454 3368 15488 3402 sw
tri 15414 3367 15415 3368 ne
rect 15415 3367 15488 3368
tri 15488 3367 15489 3368 sw
rect 11494 3302 11552 3340
tri 15415 3330 15452 3367 ne
rect 15452 3330 15489 3367
tri 15489 3330 15526 3367 sw
rect 11494 3268 11506 3302
rect 11540 3268 11552 3302
tri 15452 3301 15481 3330 ne
rect 15481 3301 15526 3330
tri 15526 3301 15555 3330 sw
rect 11494 3230 11552 3268
rect 11494 3196 11506 3230
rect 11540 3196 11552 3230
rect 11494 3158 11552 3196
rect 11494 3124 11506 3158
rect 11540 3124 11552 3158
rect 11494 3086 11552 3124
rect 11612 3249 11619 3301
rect 11671 3249 11683 3301
rect 11735 3249 11742 3301
rect 14353 3249 14359 3301
rect 14411 3249 14423 3301
rect 14475 3299 14483 3301
rect 14484 3300 14510 3301
rect 14511 3299 15335 3301
rect 14475 3296 15335 3299
tri 15335 3296 15340 3301 sw
tri 15481 3296 15486 3301 ne
rect 15486 3296 15555 3301
tri 15555 3296 15560 3301 sw
rect 14475 3292 15340 3296
rect 14475 3258 14526 3292
rect 14560 3258 14598 3292
rect 14632 3258 15340 3292
tri 15340 3258 15378 3296 sw
tri 15486 3293 15489 3296 ne
rect 15489 3293 15560 3296
tri 15560 3293 15563 3296 sw
tri 15489 3271 15511 3293 ne
rect 14475 3251 15378 3258
rect 14475 3249 14483 3251
rect 14484 3249 14510 3250
rect 14511 3249 15378 3251
tri 15378 3249 15387 3258 sw
rect 11612 3147 11742 3249
tri 15313 3227 15335 3249 ne
rect 15335 3227 15387 3249
tri 15387 3227 15409 3249 sw
tri 15335 3224 15338 3227 ne
rect 15338 3224 15409 3227
tri 15409 3224 15412 3227 sw
tri 15338 3186 15376 3224 ne
rect 15376 3186 15412 3224
tri 15412 3186 15450 3224 sw
tri 15376 3153 15409 3186 ne
rect 15409 3153 15450 3186
tri 15450 3153 15483 3186 sw
tri 15409 3152 15410 3153 ne
rect 15410 3152 15483 3153
tri 15410 3147 15415 3152 ne
rect 15415 3147 15483 3152
rect 11612 3095 11619 3147
rect 11671 3095 11683 3147
rect 11735 3095 11742 3147
rect 14349 3095 14355 3147
rect 14407 3095 14419 3147
rect 14471 3095 14479 3147
rect 14480 3096 14481 3146
rect 14509 3096 14510 3146
rect 14511 3138 15269 3147
rect 14511 3104 14526 3138
rect 14560 3104 14598 3138
rect 14632 3131 15269 3138
tri 15269 3131 15285 3147 sw
tri 15415 3131 15431 3147 ne
rect 14632 3114 15285 3131
tri 15285 3114 15302 3131 sw
rect 14632 3104 15302 3114
rect 14511 3095 15302 3104
tri 15302 3095 15321 3114 sw
tri 15247 3087 15255 3095 ne
rect 15255 3087 15321 3095
tri 15321 3087 15329 3095 sw
rect 11494 3052 11506 3086
rect 11540 3052 11552 3086
tri 15255 3080 15262 3087 ne
rect 15262 3080 15329 3087
tri 15329 3080 15336 3087 sw
tri 15262 3073 15269 3080 ne
rect 15269 3073 15336 3080
rect 11494 3014 11552 3052
tri 15269 3042 15300 3073 ne
rect 15300 3042 15336 3073
tri 15336 3042 15374 3080 sw
rect 11494 2980 11506 3014
rect 11540 2980 11552 3014
tri 15300 3013 15329 3042 ne
rect 15329 3013 15374 3042
tri 15374 3013 15403 3042 sw
tri 15329 3008 15334 3013 ne
rect 15334 3008 15403 3013
tri 15334 2993 15349 3008 ne
rect 15349 2993 15403 3008
rect 11494 2942 11552 2980
rect 11494 2908 11506 2942
rect 11540 2908 11552 2942
rect 11494 2870 11552 2908
rect 11494 2836 11506 2870
rect 11540 2836 11552 2870
rect 11494 2798 11552 2836
rect 11494 2764 11506 2798
rect 11540 2764 11552 2798
rect 11612 2941 11619 2993
rect 11671 2941 11683 2993
rect 11735 2941 11742 2993
rect 14353 2941 14359 2993
rect 14411 2941 14423 2993
rect 14475 2991 14483 2993
rect 14484 2992 14510 2993
rect 14511 2991 15203 2993
rect 14475 2984 15203 2991
rect 14475 2950 14526 2984
rect 14560 2950 14598 2984
rect 14632 2970 15203 2984
tri 15203 2970 15226 2993 sw
tri 15349 2991 15351 2993 ne
rect 14632 2950 15226 2970
rect 14475 2947 15226 2950
tri 15226 2947 15249 2970 sw
rect 14475 2943 15249 2947
rect 14475 2941 14483 2943
rect 14484 2941 14510 2942
rect 14511 2941 15249 2943
tri 15249 2941 15255 2947 sw
rect 11612 2839 11742 2941
tri 15181 2936 15186 2941 ne
rect 15186 2936 15255 2941
tri 15255 2936 15260 2941 sw
tri 15186 2898 15224 2936 ne
rect 15224 2898 15260 2936
tri 15260 2898 15298 2936 sw
tri 15224 2873 15249 2898 ne
rect 15249 2873 15298 2898
tri 15298 2873 15323 2898 sw
tri 15249 2864 15258 2873 ne
rect 15258 2864 15323 2873
tri 15258 2851 15271 2864 ne
rect 11612 2787 11619 2839
rect 11671 2787 11683 2839
rect 11735 2787 11742 2839
rect 14349 2787 14355 2839
rect 14407 2787 14419 2839
rect 14471 2787 14479 2839
rect 14480 2788 14481 2838
rect 14509 2788 14510 2838
rect 14511 2830 15137 2839
rect 14511 2796 14526 2830
rect 14560 2796 14598 2830
rect 14632 2826 15137 2830
tri 15137 2826 15150 2839 sw
rect 14632 2807 15150 2826
tri 15150 2807 15169 2826 sw
rect 14632 2796 15169 2807
rect 14511 2792 15169 2796
tri 15169 2792 15184 2807 sw
rect 14511 2787 15184 2792
tri 15184 2787 15189 2792 sw
rect 11494 2726 11552 2764
tri 15115 2754 15148 2787 ne
rect 15148 2754 15189 2787
tri 15189 2754 15222 2787 sw
tri 15148 2733 15169 2754 ne
rect 15169 2733 15222 2754
tri 15222 2733 15243 2754 sw
rect 11494 2692 11506 2726
rect 11540 2692 11552 2726
tri 15169 2720 15182 2733 ne
rect 15182 2720 15243 2733
tri 15182 2711 15191 2720 ne
rect 11494 2654 11552 2692
rect 11494 2620 11506 2654
rect 11540 2620 11552 2654
rect 11494 2582 11552 2620
rect 11494 2548 11506 2582
rect 11540 2548 11552 2582
rect 11494 2510 11552 2548
rect 11494 2476 11506 2510
rect 11540 2476 11552 2510
rect 11612 2633 11619 2685
rect 11671 2633 11683 2685
rect 11735 2633 11742 2685
rect 14353 2633 14359 2685
rect 14411 2633 14423 2685
rect 14475 2683 14483 2685
rect 14484 2684 14510 2685
rect 14511 2683 15071 2685
rect 14475 2681 15071 2683
tri 15071 2681 15075 2685 sw
rect 14475 2676 15075 2681
rect 14475 2642 14526 2676
rect 14560 2642 14598 2676
rect 14632 2667 15075 2676
tri 15075 2667 15089 2681 sw
rect 14632 2647 15089 2667
tri 15089 2647 15109 2667 sw
rect 14632 2642 15109 2647
rect 14475 2635 15109 2642
rect 14475 2633 14483 2635
rect 14484 2633 14510 2634
rect 14511 2633 15109 2635
tri 15109 2633 15123 2647 sw
rect 11612 2531 11742 2633
tri 15049 2608 15074 2633 ne
rect 15074 2608 15123 2633
tri 15123 2608 15148 2633 sw
tri 15074 2593 15089 2608 ne
rect 15089 2593 15148 2608
tri 15148 2593 15163 2608 sw
tri 15089 2574 15108 2593 ne
rect 15108 2574 15163 2593
tri 15108 2571 15111 2574 ne
rect 11612 2479 11619 2531
rect 11671 2479 11683 2531
rect 11735 2479 11742 2531
rect 14349 2479 14355 2531
rect 14407 2479 14419 2531
rect 14471 2479 14479 2531
rect 14480 2480 14481 2530
rect 14511 2530 14859 2531
tri 14859 2530 14860 2531 sw
rect 14509 2480 14510 2530
rect 14511 2522 14860 2530
rect 14511 2488 14526 2522
rect 14560 2488 14598 2522
rect 14632 2501 14860 2522
tri 14860 2501 14889 2530 sw
rect 14632 2488 14889 2501
rect 14511 2479 14889 2488
tri 14889 2479 14911 2501 sw
rect 11494 2438 11552 2476
tri 14837 2462 14854 2479 ne
rect 14854 2462 14911 2479
tri 14911 2462 14928 2479 sw
tri 14854 2456 14860 2462 ne
rect 14860 2456 14928 2462
tri 14928 2456 14934 2462 sw
rect 11494 2404 11506 2438
rect 11540 2404 11552 2438
tri 14860 2428 14888 2456 ne
rect 14888 2428 14934 2456
tri 14934 2428 14962 2456 sw
rect 11494 2366 11552 2404
tri 14888 2389 14927 2428 ne
rect 14927 2389 14962 2428
tri 14962 2389 15001 2428 sw
tri 14927 2382 14934 2389 ne
rect 14934 2382 15001 2389
tri 15001 2382 15008 2389 sw
tri 14934 2377 14939 2382 ne
rect 14939 2377 15008 2382
tri 15008 2377 15013 2382 sw
rect 11494 2332 11506 2366
rect 11540 2332 11552 2366
rect 11494 2294 11552 2332
rect 11494 2260 11506 2294
rect 11540 2260 11552 2294
rect 11494 2222 11552 2260
rect 11494 2188 11506 2222
rect 11540 2188 11552 2222
rect 11494 2150 11552 2188
rect 11612 2325 11619 2377
rect 11671 2325 11683 2377
rect 11735 2325 11742 2377
rect 14353 2325 14359 2377
rect 14411 2325 14423 2377
rect 14475 2375 14483 2377
rect 14484 2376 14510 2377
rect 14511 2375 14866 2377
rect 14475 2368 14866 2375
rect 14475 2334 14526 2368
rect 14560 2334 14598 2368
rect 14632 2355 14866 2368
tri 14866 2355 14888 2377 sw
tri 14939 2355 14961 2377 ne
rect 14961 2355 15013 2377
tri 15013 2355 15035 2377 sw
rect 14632 2334 14888 2355
rect 14475 2327 14888 2334
rect 14475 2325 14483 2327
rect 14484 2325 14510 2326
rect 14511 2325 14888 2327
tri 14888 2325 14918 2355 sw
tri 14961 2325 14991 2355 ne
rect 14991 2325 15035 2355
tri 15035 2325 15065 2355 sw
rect 11612 2223 11742 2325
tri 14844 2316 14853 2325 ne
rect 14853 2316 14918 2325
tri 14918 2316 14927 2325 sw
tri 14991 2316 15000 2325 ne
rect 15000 2316 15065 2325
tri 15065 2316 15074 2325 sw
tri 14853 2303 14866 2316 ne
rect 14866 2315 14927 2316
tri 14927 2315 14928 2316 sw
tri 15000 2315 15001 2316 ne
rect 15001 2315 15074 2316
rect 14866 2308 14928 2315
tri 14928 2308 14935 2315 sw
tri 15001 2308 15008 2315 ne
rect 15008 2308 15074 2315
tri 15074 2308 15082 2316 sw
rect 14866 2303 14935 2308
tri 14866 2282 14887 2303 ne
rect 14887 2286 14935 2303
tri 14935 2286 14957 2308 sw
tri 15008 2286 15030 2308 ne
rect 14887 2282 14957 2286
tri 14957 2282 14961 2286 sw
tri 14887 2243 14926 2282 ne
rect 14926 2243 14961 2282
tri 14961 2243 15000 2282 sw
tri 14926 2242 14927 2243 ne
rect 14927 2242 15000 2243
tri 15000 2242 15001 2243 sw
tri 14927 2223 14946 2242 ne
rect 14946 2223 15001 2242
rect 11612 2171 11619 2223
rect 11671 2171 11683 2223
rect 11735 2171 11742 2223
rect 14349 2171 14355 2223
rect 14407 2171 14419 2223
rect 14471 2171 14479 2223
rect 14480 2172 14481 2222
rect 14509 2172 14510 2222
rect 14511 2220 14873 2223
tri 14873 2220 14876 2223 sw
tri 14946 2220 14949 2223 ne
rect 14511 2214 14876 2220
rect 14511 2180 14526 2214
rect 14560 2180 14598 2214
rect 14632 2209 14876 2214
tri 14876 2209 14887 2220 sw
rect 14632 2180 14887 2209
rect 14511 2176 14887 2180
tri 14887 2176 14920 2209 sw
rect 14511 2171 14920 2176
tri 14815 2170 14816 2171 ne
rect 14816 2170 14920 2171
rect 11494 2116 11506 2150
rect 11540 2116 11552 2150
tri 14816 2136 14850 2170 ne
rect 14850 2136 14920 2170
tri 14850 2118 14868 2136 ne
rect 11494 2097 11552 2116
tri 11552 2097 11559 2104 sw
rect 11494 2078 11559 2097
tri 11559 2078 11578 2097 sw
rect 11494 2044 11506 2078
rect 11540 2044 11585 2078
rect 11637 2069 11649 2078
rect 11701 2069 11713 2078
rect 11765 2069 11777 2078
rect 11829 2069 11841 2078
rect 11893 2069 11905 2078
rect 11957 2069 11969 2078
rect 11494 2026 11585 2044
rect 11642 2035 11649 2069
rect 11893 2035 11896 2069
rect 11957 2035 11968 2069
rect 11637 2026 11649 2035
rect 11701 2026 11713 2035
rect 11765 2026 11777 2035
rect 11829 2026 11841 2035
rect 11893 2026 11905 2035
rect 11957 2026 11969 2035
rect 12021 2026 12033 2078
rect 12085 2026 12097 2078
rect 12149 2026 12161 2078
rect 12213 2069 12225 2078
rect 12277 2069 12289 2078
rect 12341 2069 12353 2078
rect 12405 2069 12417 2078
rect 12469 2069 12481 2078
rect 12533 2069 12545 2078
rect 12218 2035 12225 2069
rect 12469 2035 12472 2069
rect 12533 2035 12544 2069
rect 12213 2026 12225 2035
rect 12277 2026 12289 2035
rect 12341 2026 12353 2035
rect 12405 2026 12417 2035
rect 12469 2026 12481 2035
rect 12533 2026 12545 2035
rect 12597 2026 12609 2078
rect 12661 2026 12673 2078
rect 12725 2026 12737 2078
rect 12789 2069 12801 2078
rect 12853 2069 12865 2078
rect 12917 2069 12929 2078
rect 12981 2069 12993 2078
rect 13045 2069 13057 2078
rect 13109 2069 13121 2078
rect 12794 2035 12801 2069
rect 13045 2035 13048 2069
rect 13109 2035 13120 2069
rect 12789 2026 12801 2035
rect 12853 2026 12865 2035
rect 12917 2026 12929 2035
rect 12981 2026 12993 2035
rect 13045 2026 13057 2035
rect 13109 2026 13121 2035
rect 13173 2026 13185 2078
rect 13237 2026 13249 2078
rect 13301 2026 13313 2078
rect 13365 2069 13377 2078
rect 13429 2069 13441 2078
rect 13493 2069 13505 2078
rect 13557 2069 13569 2078
rect 13621 2069 13633 2078
rect 13685 2069 13697 2078
rect 13370 2035 13377 2069
rect 13621 2035 13624 2069
rect 13685 2035 13696 2069
rect 13365 2026 13377 2035
rect 13429 2026 13441 2035
rect 13493 2026 13505 2035
rect 13557 2026 13569 2035
rect 13621 2026 13633 2035
rect 13685 2026 13697 2035
rect 13749 2026 13761 2078
rect 13813 2026 13825 2078
rect 13877 2026 13889 2078
rect 13941 2069 13953 2078
rect 14005 2069 14017 2078
rect 14069 2069 14081 2078
rect 14133 2069 14145 2078
rect 14197 2069 14209 2078
rect 14261 2069 14273 2078
rect 13946 2035 13953 2069
rect 14197 2035 14200 2069
rect 14261 2035 14272 2069
rect 13941 2026 13953 2035
rect 14005 2026 14017 2035
rect 14069 2026 14081 2035
rect 14133 2026 14145 2035
rect 14197 2026 14209 2035
rect 14261 2026 14273 2035
rect 14325 2026 14337 2078
rect 14389 2026 14401 2078
rect 14453 2026 14465 2078
rect 14517 2069 14529 2078
rect 14581 2069 14593 2078
rect 14645 2069 14657 2078
rect 14709 2069 14721 2078
rect 14522 2035 14529 2069
rect 14517 2026 14529 2035
rect 14581 2026 14593 2035
rect 14645 2026 14657 2035
rect 14709 2026 14721 2035
rect 14773 2026 14779 2078
tri 14834 1990 14868 2024 se
rect 14868 2002 14920 2136
rect 14868 1990 14908 2002
tri 14908 1990 14920 2002 nw
tri 14802 1958 14834 1990 se
rect 14834 1958 14876 1990
tri 14876 1958 14908 1990 nw
tri 14795 1951 14802 1958 se
rect 14802 1951 14869 1958
tri 14869 1951 14876 1958 nw
tri 14942 1951 14949 1958 se
rect 14949 1951 15001 2223
tri 14794 1950 14795 1951 se
rect 14795 1950 14868 1951
tri 14868 1950 14869 1951 nw
tri 14941 1950 14942 1951 se
rect 14942 1950 15001 1951
tri 14777 1933 14794 1950 se
rect 14794 1933 14851 1950
tri 14851 1933 14868 1950 nw
tri 14924 1933 14941 1950 se
rect 14941 1936 15001 1950
rect 14941 1933 14982 1936
rect 12870 1924 14835 1933
rect 12870 1890 12882 1924
rect 12916 1890 12954 1924
rect 12988 1917 14835 1924
tri 14835 1917 14851 1933 nw
tri 14908 1917 14924 1933 se
rect 14924 1917 14982 1933
tri 14982 1917 15001 1936 nw
rect 12988 1892 14810 1917
tri 14810 1892 14835 1917 nw
tri 14883 1892 14908 1917 se
rect 14908 1892 14957 1917
tri 14957 1892 14982 1917 nw
rect 12988 1890 14804 1892
rect 12870 1886 14804 1890
tri 14804 1886 14810 1892 nw
tri 14877 1886 14883 1892 se
rect 14883 1886 14949 1892
rect 12870 1884 13196 1886
tri 13196 1884 13198 1886 nw
tri 13837 1884 13839 1886 ne
rect 13839 1884 14802 1886
tri 14802 1884 14804 1886 nw
tri 14875 1884 14877 1886 se
rect 14877 1884 14949 1886
tri 14949 1884 14957 1892 nw
tri 15022 1884 15030 1892 se
rect 15030 1884 15082 2308
rect 12870 1881 13193 1884
tri 13193 1881 13196 1884 nw
tri 13839 1881 13842 1884 ne
rect 13842 1881 14799 1884
tri 14799 1881 14802 1884 nw
tri 14872 1881 14875 1884 se
rect 14875 1881 14946 1884
tri 14946 1881 14949 1884 nw
tri 15019 1881 15022 1884 se
rect 15022 1881 15082 1884
tri 14869 1878 14872 1881 se
rect 14872 1878 14943 1881
tri 14943 1878 14946 1881 nw
tri 15016 1878 15019 1881 se
rect 15019 1878 15082 1881
tri 14847 1856 14869 1878 se
rect 14869 1856 14921 1878
tri 14921 1856 14943 1878 nw
tri 14994 1856 15016 1878 se
rect 15016 1870 15082 1878
rect 15016 1856 15056 1870
tri 13245 1853 13248 1856 se
rect 13248 1853 13254 1856
rect 13156 1847 13254 1853
rect 13306 1847 13322 1856
rect 13156 1813 13168 1847
rect 13202 1813 13244 1847
rect 13306 1813 13320 1847
rect 13156 1807 13254 1813
tri 13245 1805 13247 1807 ne
rect 13247 1805 13254 1807
tri 13247 1804 13248 1805 ne
rect 13248 1804 13254 1805
rect 13306 1804 13322 1813
rect 13374 1804 13390 1856
rect 13442 1804 13458 1856
rect 13510 1804 13526 1856
rect 13578 1847 13594 1856
rect 13646 1847 13662 1856
rect 13714 1847 13730 1856
rect 13782 1853 13788 1856
tri 13788 1853 13791 1856 sw
tri 14844 1853 14847 1856 se
rect 14847 1853 14918 1856
tri 14918 1853 14921 1856 nw
tri 14991 1853 14994 1856 se
rect 14994 1853 15056 1856
rect 13782 1847 14647 1853
rect 13582 1813 13594 1847
rect 13658 1813 13662 1847
rect 13810 1813 13851 1847
rect 13885 1813 13926 1847
rect 13960 1813 14001 1847
rect 14035 1813 14076 1847
rect 14110 1813 14151 1847
rect 14185 1813 14226 1847
rect 14260 1813 14301 1847
rect 14335 1813 14376 1847
rect 14410 1813 14451 1847
rect 14485 1813 14526 1847
rect 14560 1813 14601 1847
rect 14635 1813 14647 1847
tri 14835 1844 14844 1853 se
rect 14844 1844 14909 1853
tri 14909 1844 14918 1853 nw
tri 14982 1844 14991 1853 se
rect 14991 1844 15056 1853
tri 15056 1844 15082 1870 nw
tri 14809 1818 14835 1844 se
rect 14835 1818 14883 1844
tri 14883 1818 14909 1844 nw
tri 14956 1818 14982 1844 se
rect 14982 1818 15030 1844
tri 15030 1818 15056 1844 nw
rect 13578 1804 13594 1813
rect 13646 1804 13662 1813
rect 13714 1804 13730 1813
rect 13782 1807 14647 1813
tri 14801 1810 14809 1818 se
rect 14809 1811 14876 1818
tri 14876 1811 14883 1818 nw
tri 14949 1811 14956 1818 se
rect 14956 1811 15017 1818
rect 14809 1810 14875 1811
tri 14875 1810 14876 1811 nw
tri 14948 1810 14949 1811 se
rect 14949 1810 15017 1811
tri 14798 1807 14801 1810 se
rect 14801 1807 14872 1810
tri 14872 1807 14875 1810 nw
tri 14945 1807 14948 1810 se
rect 14948 1807 15017 1810
rect 13782 1805 13789 1807
tri 13789 1805 13791 1807 nw
tri 14796 1805 14798 1807 se
rect 14798 1805 14870 1807
tri 14870 1805 14872 1807 nw
tri 14943 1805 14945 1807 se
rect 14945 1805 15017 1807
tri 15017 1805 15030 1818 nw
rect 13782 1804 13788 1805
tri 13788 1804 13789 1805 nw
tri 14795 1804 14796 1805 se
rect 14796 1804 14869 1805
tri 14869 1804 14870 1805 nw
tri 14942 1804 14943 1805 se
rect 14943 1804 14983 1805
tri 14770 1779 14795 1804 se
rect 14795 1779 14844 1804
tri 14844 1779 14869 1804 nw
tri 14917 1779 14942 1804 se
rect 14942 1779 14983 1804
rect 10783 1727 10789 1779
rect 10841 1727 10853 1779
rect 10905 1727 10928 1779
rect 10929 1728 10930 1778
rect 10958 1728 10959 1778
rect 10960 1727 11114 1779
rect 12870 1772 13217 1779
tri 13217 1772 13224 1779 sw
tri 13818 1772 13825 1779 se
rect 13825 1772 14837 1779
tri 14837 1772 14844 1779 nw
tri 14910 1772 14917 1779 se
rect 14917 1772 14983 1779
rect 12870 1771 14836 1772
tri 14836 1771 14837 1772 nw
tri 14909 1771 14910 1772 se
rect 14910 1771 14983 1772
tri 14983 1771 15017 1805 nw
rect 12870 1770 14809 1771
rect 12870 1736 12882 1770
rect 12916 1736 12954 1770
rect 12988 1744 14809 1770
tri 14809 1744 14836 1771 nw
tri 14882 1744 14909 1771 se
rect 14909 1744 14956 1771
tri 14956 1744 14983 1771 nw
rect 12988 1736 14797 1744
rect 12870 1732 14797 1736
tri 14797 1732 14809 1744 nw
tri 14870 1732 14882 1744 se
rect 14882 1732 14944 1744
tri 14944 1732 14956 1744 nw
rect 12870 1727 14792 1732
tri 14792 1727 14797 1732 nw
tri 14865 1727 14870 1732 se
rect 14870 1727 14910 1732
tri 10960 1701 10986 1727 ne
tri 10968 1479 10986 1497 se
rect 10986 1479 11114 1727
tri 14836 1698 14865 1727 se
rect 14865 1698 14910 1727
tri 14910 1698 14944 1732 nw
tri 14808 1670 14836 1698 se
rect 14836 1670 14882 1698
tri 14882 1670 14910 1698 nw
tri 14797 1659 14808 1670 se
rect 14808 1659 14871 1670
tri 14871 1659 14882 1670 nw
tri 14763 1625 14797 1659 se
rect 14797 1625 14837 1659
tri 14837 1625 14871 1659 nw
rect 12870 1616 14819 1625
rect 12870 1582 12882 1616
rect 12916 1582 12954 1616
rect 12988 1607 14819 1616
tri 14819 1607 14837 1625 nw
rect 12988 1586 14798 1607
tri 14798 1586 14819 1607 nw
tri 15090 1586 15111 1607 se
rect 15111 1586 15163 2574
rect 12988 1582 14785 1586
rect 12870 1573 14785 1582
tri 14785 1573 14798 1586 nw
tri 15077 1573 15090 1586 se
rect 15090 1585 15163 1586
rect 15090 1573 15130 1585
tri 15056 1552 15077 1573 se
rect 15077 1552 15130 1573
tri 15130 1552 15163 1585 nw
tri 15037 1533 15056 1552 se
rect 15056 1533 15111 1552
tri 15111 1533 15130 1552 nw
tri 15017 1513 15037 1533 se
rect 15037 1513 15091 1533
tri 15091 1513 15111 1533 nw
tri 14983 1479 15017 1513 se
rect 15017 1479 15057 1513
tri 15057 1479 15091 1513 nw
tri 10960 1471 10968 1479 se
rect 10968 1471 11114 1479
tri 14975 1471 14983 1479 se
rect 14983 1471 15049 1479
tri 15049 1471 15057 1479 nw
rect 10783 1419 10789 1471
rect 10841 1419 10853 1471
rect 10905 1469 10926 1471
rect 10927 1470 10953 1471
rect 10954 1469 11114 1471
rect 10905 1421 11114 1469
rect 10905 1419 10926 1421
rect 10927 1419 10953 1420
rect 10954 1419 11114 1421
rect 12870 1462 15018 1471
rect 12870 1428 12882 1462
rect 12916 1428 12954 1462
rect 12988 1440 15018 1462
tri 15018 1440 15049 1471 nw
tri 15164 1440 15191 1467 se
rect 15191 1445 15243 2720
rect 15191 1440 15238 1445
tri 15238 1440 15243 1445 nw
rect 12988 1428 15000 1440
rect 12870 1422 15000 1428
tri 15000 1422 15018 1440 nw
tri 15146 1422 15164 1440 se
rect 15164 1422 15204 1440
rect 12870 1419 13233 1422
tri 13233 1419 13236 1422 nw
tri 13813 1419 13816 1422 ne
rect 13816 1419 14997 1422
tri 14997 1419 15000 1422 nw
tri 15143 1419 15146 1422 se
rect 15146 1419 15204 1422
tri 10960 1406 10973 1419 ne
rect 10973 1406 11114 1419
tri 15130 1406 15143 1419 se
rect 15143 1406 15204 1419
tri 15204 1406 15238 1440 nw
tri 10973 1393 10986 1406 ne
tri 10984 1187 10986 1189 se
rect 10986 1187 11114 1406
tri 15118 1394 15130 1406 se
rect 15130 1394 15191 1406
tri 13245 1391 13248 1394 se
rect 13248 1391 13254 1394
rect 13156 1385 13254 1391
rect 13306 1385 13322 1394
rect 13156 1351 13168 1385
rect 13202 1351 13244 1385
rect 13306 1351 13320 1385
rect 13156 1345 13254 1351
tri 13245 1342 13248 1345 ne
rect 13248 1342 13254 1345
rect 13306 1342 13322 1351
rect 13374 1342 13390 1394
rect 13442 1342 13458 1394
rect 13510 1342 13526 1394
rect 13578 1385 13594 1394
rect 13646 1385 13662 1394
rect 13714 1385 13730 1394
rect 13782 1393 13788 1394
tri 13788 1393 13789 1394 sw
tri 15117 1393 15118 1394 se
rect 15118 1393 15191 1394
tri 15191 1393 15204 1406 nw
rect 13782 1391 13789 1393
tri 13789 1391 13791 1393 sw
tri 15115 1391 15117 1393 se
rect 15117 1391 15165 1393
rect 13782 1385 14647 1391
rect 13582 1351 13594 1385
rect 13658 1351 13662 1385
rect 13810 1351 13851 1385
rect 13885 1351 13926 1385
rect 13960 1351 14001 1385
rect 14035 1351 14076 1385
rect 14110 1351 14151 1385
rect 14185 1351 14226 1385
rect 14260 1351 14301 1385
rect 14335 1351 14376 1385
rect 14410 1351 14451 1385
rect 14485 1351 14526 1385
rect 14560 1351 14601 1385
rect 14635 1351 14647 1385
tri 15091 1367 15115 1391 se
rect 15115 1367 15165 1391
tri 15165 1367 15191 1393 nw
rect 13578 1342 13594 1351
rect 13646 1342 13662 1351
rect 13714 1342 13730 1351
rect 13782 1345 14647 1351
tri 15069 1345 15091 1367 se
rect 15091 1345 15131 1367
rect 13782 1342 13788 1345
tri 13788 1342 13791 1345 nw
tri 15066 1342 15069 1345 se
rect 15069 1342 15131 1345
tri 15057 1333 15066 1342 se
rect 15066 1333 15131 1342
tri 15131 1333 15165 1367 nw
tri 15043 1319 15057 1333 se
rect 15057 1319 15117 1333
tri 15117 1319 15131 1333 nw
tri 15263 1319 15271 1327 se
rect 15271 1319 15323 2864
tri 15041 1317 15043 1319 se
rect 15043 1317 15115 1319
tri 15115 1317 15117 1319 nw
tri 15261 1317 15263 1319 se
rect 15263 1317 15323 1319
rect 12870 1313 13206 1317
tri 13206 1313 13210 1317 sw
tri 13821 1313 13825 1317 se
rect 13825 1313 15111 1317
tri 15111 1313 15115 1317 nw
tri 15257 1313 15261 1317 se
rect 15261 1313 15323 1317
rect 12870 1308 15092 1313
rect 12870 1274 12882 1308
rect 12916 1274 12954 1308
rect 12988 1294 15092 1308
tri 15092 1294 15111 1313 nw
tri 15238 1294 15257 1313 se
rect 15257 1305 15323 1313
rect 15257 1294 15312 1305
tri 15312 1294 15323 1305 nw
rect 12988 1274 15063 1294
rect 12870 1265 15063 1274
tri 15063 1265 15092 1294 nw
tri 15209 1265 15238 1294 se
rect 15238 1265 15278 1294
tri 15204 1260 15209 1265 se
rect 15209 1260 15278 1265
tri 15278 1260 15312 1294 nw
tri 15197 1253 15204 1260 se
rect 15204 1253 15271 1260
tri 15271 1253 15278 1260 nw
tri 15165 1221 15197 1253 se
rect 15197 1221 15239 1253
tri 15239 1221 15271 1253 nw
tri 15131 1187 15165 1221 se
rect 15165 1187 15205 1221
tri 15205 1187 15239 1221 nw
tri 10960 1163 10984 1187 se
rect 10984 1163 11114 1187
tri 15123 1179 15131 1187 se
rect 15131 1179 15197 1187
tri 15197 1179 15205 1187 nw
tri 15343 1179 15351 1187 se
rect 15351 1179 15403 2993
tri 15107 1163 15123 1179 se
rect 15123 1163 15181 1179
tri 15181 1163 15197 1179 nw
tri 15327 1163 15343 1179 se
rect 15343 1165 15403 1179
rect 15343 1163 15386 1165
rect 10783 1111 10789 1163
rect 10841 1111 10853 1163
rect 10905 1111 10928 1163
rect 10929 1112 10930 1162
rect 10958 1112 10959 1162
rect 10960 1111 11114 1163
rect 12870 1154 15166 1163
rect 12870 1120 12882 1154
rect 12916 1120 12954 1154
rect 12988 1148 15166 1154
tri 15166 1148 15181 1163 nw
tri 15312 1148 15327 1163 se
rect 15327 1148 15386 1163
tri 15386 1148 15403 1165 nw
rect 12988 1120 15133 1148
rect 12870 1115 15133 1120
tri 15133 1115 15166 1148 nw
tri 15279 1115 15312 1148 se
rect 15312 1115 15352 1148
rect 12870 1114 13221 1115
tri 13221 1114 13222 1115 nw
tri 13825 1114 13826 1115 ne
rect 13826 1114 15132 1115
tri 15132 1114 15133 1115 nw
tri 15278 1114 15279 1115 se
rect 15279 1114 15352 1115
tri 15352 1114 15386 1148 nw
rect 12870 1111 13218 1114
tri 13218 1111 13221 1114 nw
tri 13826 1111 13829 1114 ne
rect 13829 1111 15129 1114
tri 15129 1111 15132 1114 nw
tri 15277 1113 15278 1114 se
rect 15278 1113 15351 1114
tri 15351 1113 15352 1114 nw
tri 15275 1111 15277 1113 se
rect 15277 1111 15313 1113
tri 10960 1085 10986 1111 ne
tri 10961 856 10986 881 se
rect 10986 856 11114 1111
tri 15250 1086 15275 1111 se
rect 15275 1086 15313 1111
tri 13245 1083 13248 1086 se
rect 13248 1083 13254 1086
rect 13156 1077 13254 1083
rect 13306 1077 13322 1086
rect 13156 1043 13168 1077
rect 13202 1043 13244 1077
rect 13306 1043 13320 1077
rect 13156 1037 13254 1043
tri 13245 1034 13248 1037 ne
rect 13248 1034 13254 1037
rect 13306 1034 13322 1043
rect 13374 1034 13390 1086
rect 13442 1034 13458 1086
rect 13510 1034 13526 1086
rect 13578 1077 13594 1086
rect 13646 1077 13662 1086
rect 13714 1077 13730 1086
rect 13782 1083 13788 1086
tri 13788 1083 13791 1086 sw
tri 15247 1083 15250 1086 se
rect 15250 1083 15313 1086
rect 13782 1077 14647 1083
rect 13582 1043 13594 1077
rect 13658 1043 13662 1077
rect 13810 1043 13851 1077
rect 13885 1043 13926 1077
rect 13960 1043 14001 1077
rect 14035 1043 14076 1077
rect 14110 1043 14151 1077
rect 14185 1043 14226 1077
rect 14260 1043 14301 1077
rect 14335 1043 14376 1077
rect 14410 1043 14451 1077
rect 14485 1043 14526 1077
rect 14560 1043 14601 1077
rect 14635 1043 14647 1077
tri 15239 1075 15247 1083 se
rect 15247 1075 15313 1083
tri 15313 1075 15351 1113 nw
tri 15211 1047 15239 1075 se
rect 15239 1047 15285 1075
tri 15285 1047 15313 1075 nw
rect 13578 1034 13594 1043
rect 13646 1034 13662 1043
rect 13714 1034 13730 1043
rect 13782 1037 14647 1043
tri 15205 1041 15211 1047 se
rect 15211 1041 15279 1047
tri 15279 1041 15285 1047 nw
tri 15425 1041 15431 1047 se
rect 15431 1041 15483 3147
tri 15203 1039 15205 1041 se
rect 15205 1039 15277 1041
tri 15277 1039 15279 1041 nw
tri 15423 1039 15425 1041 se
rect 15425 1039 15483 1041
tri 15201 1037 15203 1039 se
rect 15203 1037 15247 1039
rect 13782 1034 13788 1037
tri 13788 1034 13791 1037 nw
tri 15198 1034 15201 1037 se
rect 15201 1034 15247 1037
tri 15173 1009 15198 1034 se
rect 15198 1009 15247 1034
tri 15247 1009 15277 1039 nw
tri 15393 1009 15423 1039 se
rect 15423 1025 15483 1039
rect 15423 1009 15460 1025
rect 12870 1004 13215 1009
tri 13215 1004 13220 1009 sw
tri 13812 1004 13817 1009 se
rect 13817 1004 15242 1009
tri 15242 1004 15247 1009 nw
tri 15388 1004 15393 1009 se
rect 15393 1004 15460 1009
rect 12870 1002 15240 1004
tri 15240 1002 15242 1004 nw
tri 15386 1002 15388 1004 se
rect 15388 1002 15460 1004
tri 15460 1002 15483 1025 nw
rect 12870 1000 15211 1002
rect 12870 966 12882 1000
rect 12916 966 12954 1000
rect 12988 973 15211 1000
tri 15211 973 15240 1002 nw
tri 15357 973 15386 1002 se
rect 15386 973 15431 1002
tri 15431 973 15460 1002 nw
rect 12988 968 15206 973
tri 15206 968 15211 973 nw
tri 15352 968 15357 973 se
rect 15357 968 15426 973
tri 15426 968 15431 973 nw
rect 12988 966 15195 968
rect 12870 957 15195 966
tri 15195 957 15206 968 nw
tri 15341 957 15352 968 se
rect 15352 957 15387 968
tri 15313 929 15341 957 se
rect 15341 929 15387 957
tri 15387 929 15426 968 nw
tri 15283 899 15313 929 se
rect 15313 899 15357 929
tri 15357 899 15387 929 nw
tri 15503 899 15511 907 se
rect 15511 899 15563 3293
tri 15279 895 15283 899 se
rect 15283 895 15353 899
tri 15353 895 15357 899 nw
tri 15499 895 15503 899 se
rect 15503 895 15563 899
tri 15240 856 15279 895 se
rect 15279 856 15314 895
tri 15314 856 15353 895 nw
tri 15460 856 15499 895 se
rect 15499 885 15563 895
rect 15499 856 15534 885
tri 15534 856 15563 885 nw
tri 10960 855 10961 856 se
rect 10961 855 11114 856
tri 15239 855 15240 856 se
rect 15240 855 15313 856
tri 15313 855 15314 856 nw
tri 15459 855 15460 856 se
rect 15460 855 15511 856
rect 10783 803 10789 855
rect 10841 803 10853 855
rect 10905 803 10928 855
rect 10929 804 10930 854
rect 10958 804 10959 854
rect 10960 803 11114 855
rect 12870 846 15280 855
rect 12870 812 12882 846
rect 12916 812 12954 846
rect 12988 822 15280 846
tri 15280 822 15313 855 nw
tri 15437 833 15459 855 se
rect 15459 833 15511 855
tri 15511 833 15534 856 nw
tri 15426 822 15437 833 se
rect 15437 822 15500 833
tri 15500 822 15511 833 nw
rect 12988 812 15264 822
rect 12870 806 15264 812
tri 15264 806 15280 822 nw
tri 15410 806 15426 822 se
rect 15426 806 15461 822
rect 12870 803 13227 806
tri 13227 803 13230 806 nw
tri 13818 803 13821 806 ne
rect 13821 803 15261 806
tri 15261 803 15264 806 nw
tri 15407 803 15410 806 se
rect 15410 803 15461 806
tri 10960 783 10980 803 ne
rect 10980 783 11114 803
tri 15387 783 15407 803 se
rect 15407 783 15461 803
tri 15461 783 15500 822 nw
tri 10980 777 10986 783 ne
tri 10977 564 10986 573 se
rect 10986 564 11114 783
tri 15382 778 15387 783 se
rect 15387 778 15437 783
tri 13245 775 13248 778 se
rect 13248 775 13254 778
rect 13156 769 13254 775
rect 13306 769 13322 778
rect 13156 735 13168 769
rect 13202 735 13244 769
rect 13306 735 13320 769
rect 13156 729 13254 735
tri 13245 726 13248 729 ne
rect 13248 726 13254 729
rect 13306 726 13322 735
rect 13374 726 13390 778
rect 13442 726 13458 778
rect 13510 726 13526 778
rect 13578 769 13594 778
rect 13646 769 13662 778
rect 13714 769 13730 778
rect 13782 775 13788 778
tri 13788 775 13791 778 sw
tri 15379 775 15382 778 se
rect 15382 775 15437 778
rect 13782 769 14647 775
rect 13582 735 13594 769
rect 13658 735 13662 769
rect 13810 735 13851 769
rect 13885 735 13926 769
rect 13960 735 14001 769
rect 14035 735 14076 769
rect 14110 735 14151 769
rect 14185 735 14226 769
rect 14260 735 14301 769
rect 14335 735 14376 769
rect 14410 735 14451 769
rect 14485 735 14526 769
rect 14560 735 14601 769
rect 14635 735 14647 769
tri 15363 759 15379 775 se
rect 15379 759 15437 775
tri 15437 759 15461 783 nw
tri 15583 759 15591 767 se
rect 15591 759 15643 3433
tri 15353 749 15363 759 se
rect 15363 749 15427 759
tri 15427 749 15437 759 nw
tri 15573 749 15583 759 se
rect 15583 749 15643 759
rect 13578 726 13594 735
rect 13646 726 13662 735
rect 13714 726 13730 735
rect 13782 729 14647 735
tri 15333 729 15353 749 se
rect 15353 729 15388 749
rect 13782 726 13788 729
tri 13788 726 13791 729 nw
tri 15330 726 15333 729 se
rect 15333 726 15388 729
tri 15314 710 15330 726 se
rect 15330 710 15388 726
tri 15388 710 15427 749 nw
tri 15534 710 15573 749 se
rect 15573 745 15643 749
rect 15573 710 15608 745
tri 15608 710 15643 745 nw
rect 15725 3402 16033 3440
rect 15725 3368 15733 3402
rect 15767 3368 15819 3402
rect 15853 3368 15905 3402
rect 15939 3368 15991 3402
rect 16025 3368 16033 3402
rect 15725 3330 16033 3368
rect 15725 3296 15733 3330
rect 15767 3296 15819 3330
rect 15853 3296 15905 3330
rect 15939 3296 15991 3330
rect 16025 3296 16033 3330
rect 15725 3258 16033 3296
rect 15725 3224 15733 3258
rect 15767 3224 15819 3258
rect 15853 3224 15905 3258
rect 15939 3224 15991 3258
rect 16025 3224 16033 3258
rect 15725 3186 16033 3224
rect 15725 3152 15733 3186
rect 15767 3152 15819 3186
rect 15853 3152 15905 3186
rect 15939 3152 15991 3186
rect 16025 3152 16033 3186
rect 15725 3114 16033 3152
rect 15725 3080 15733 3114
rect 15767 3080 15819 3114
rect 15853 3080 15905 3114
rect 15939 3080 15991 3114
rect 16025 3080 16033 3114
rect 15725 3042 16033 3080
rect 15725 3008 15733 3042
rect 15767 3008 15819 3042
rect 15853 3008 15905 3042
rect 15939 3008 15991 3042
rect 16025 3008 16033 3042
rect 15725 2970 16033 3008
rect 15725 2936 15733 2970
rect 15767 2936 15819 2970
rect 15853 2936 15905 2970
rect 15939 2936 15991 2970
rect 16025 2936 16033 2970
rect 15725 2898 16033 2936
rect 15725 2864 15733 2898
rect 15767 2864 15819 2898
rect 15853 2864 15905 2898
rect 15939 2864 15991 2898
rect 16025 2864 16033 2898
rect 15725 2826 16033 2864
rect 15725 2792 15733 2826
rect 15767 2792 15819 2826
rect 15853 2792 15905 2826
rect 15939 2792 15991 2826
rect 16025 2792 16033 2826
rect 15725 2754 16033 2792
rect 15725 2720 15733 2754
rect 15767 2720 15819 2754
rect 15853 2720 15905 2754
rect 15939 2720 15991 2754
rect 16025 2720 16033 2754
rect 15725 2681 16033 2720
rect 15725 2647 15733 2681
rect 15767 2647 15819 2681
rect 15853 2647 15905 2681
rect 15939 2647 15991 2681
rect 16025 2647 16033 2681
rect 15725 2608 16033 2647
rect 15725 2574 15733 2608
rect 15767 2574 15819 2608
rect 15853 2574 15905 2608
rect 15939 2574 15991 2608
rect 16025 2574 16033 2608
rect 15725 2535 16033 2574
rect 15725 2501 15733 2535
rect 15767 2501 15819 2535
rect 15853 2501 15905 2535
rect 15939 2501 15991 2535
rect 16025 2501 16033 2535
rect 15725 2462 16033 2501
rect 15725 2428 15733 2462
rect 15767 2428 15819 2462
rect 15853 2428 15905 2462
rect 15939 2428 15991 2462
rect 16025 2428 16033 2462
rect 15725 2389 16033 2428
rect 15725 2355 15733 2389
rect 15767 2355 15819 2389
rect 15853 2355 15905 2389
rect 15939 2355 15991 2389
rect 16025 2355 16033 2389
rect 15725 2316 16033 2355
rect 15725 2282 15733 2316
rect 15767 2282 15819 2316
rect 15853 2282 15905 2316
rect 15939 2282 15991 2316
rect 16025 2282 16033 2316
rect 15725 2243 16033 2282
rect 15725 2209 15733 2243
rect 15767 2209 15819 2243
rect 15853 2209 15905 2243
rect 15939 2209 15991 2243
rect 16025 2209 16033 2243
rect 15725 2170 16033 2209
rect 15725 2136 15733 2170
rect 15767 2136 15819 2170
rect 15853 2136 15905 2170
rect 15939 2136 15991 2170
rect 16025 2136 16033 2170
rect 15725 2097 16033 2136
rect 15725 2063 15733 2097
rect 15767 2063 15819 2097
rect 15853 2063 15905 2097
rect 15939 2063 15991 2097
rect 16025 2063 16033 2097
rect 15725 2024 16033 2063
rect 15725 1990 15733 2024
rect 15767 1990 15819 2024
rect 15853 1990 15905 2024
rect 15939 1990 15991 2024
rect 16025 1990 16033 2024
rect 15725 1951 16033 1990
rect 15725 1917 15733 1951
rect 15767 1917 15819 1951
rect 15853 1917 15905 1951
rect 15939 1917 15991 1951
rect 16025 1917 16033 1951
rect 15725 1878 16033 1917
rect 15725 1844 15733 1878
rect 15767 1844 15819 1878
rect 15853 1844 15905 1878
rect 15939 1844 15991 1878
rect 16025 1844 16033 1878
rect 15725 1805 16033 1844
rect 15725 1771 15733 1805
rect 15767 1771 15819 1805
rect 15853 1771 15905 1805
rect 15939 1771 15991 1805
rect 16025 1771 16033 1805
rect 15725 1732 16033 1771
rect 15725 1698 15733 1732
rect 15767 1698 15819 1732
rect 15853 1698 15905 1732
rect 15939 1698 15991 1732
rect 16025 1698 16033 1732
rect 15725 1659 16033 1698
rect 15725 1625 15733 1659
rect 15767 1625 15819 1659
rect 15853 1625 15905 1659
rect 15939 1625 15991 1659
rect 16025 1625 16033 1659
rect 15725 1586 16033 1625
rect 15725 1552 15733 1586
rect 15767 1552 15819 1586
rect 15853 1552 15905 1586
rect 15939 1552 15991 1586
rect 16025 1552 16033 1586
rect 15725 1513 16033 1552
rect 15725 1479 15733 1513
rect 15767 1479 15819 1513
rect 15853 1479 15905 1513
rect 15939 1479 15991 1513
rect 16025 1479 16033 1513
rect 15725 1440 16033 1479
rect 15725 1406 15733 1440
rect 15767 1406 15819 1440
rect 15853 1406 15905 1440
rect 15939 1406 15991 1440
rect 16025 1406 16033 1440
rect 15725 1367 16033 1406
rect 15725 1333 15733 1367
rect 15767 1333 15819 1367
rect 15853 1333 15905 1367
rect 15939 1333 15991 1367
rect 16025 1333 16033 1367
rect 15725 1294 16033 1333
rect 15725 1260 15733 1294
rect 15767 1260 15819 1294
rect 15853 1260 15905 1294
rect 15939 1260 15991 1294
rect 16025 1260 16033 1294
rect 15725 1221 16033 1260
rect 15725 1187 15733 1221
rect 15767 1187 15819 1221
rect 15853 1187 15905 1221
rect 15939 1187 15991 1221
rect 16025 1187 16033 1221
rect 15725 1148 16033 1187
rect 15725 1114 15733 1148
rect 15767 1114 15819 1148
rect 15853 1114 15905 1148
rect 15939 1114 15991 1148
rect 16025 1114 16033 1148
rect 15725 1075 16033 1114
rect 15725 1041 15733 1075
rect 15767 1041 15819 1075
rect 15853 1041 15905 1075
rect 15939 1041 15991 1075
rect 16025 1041 16033 1075
rect 15725 1002 16033 1041
rect 15725 968 15733 1002
rect 15767 968 15819 1002
rect 15853 968 15905 1002
rect 15939 968 15991 1002
rect 16025 968 16033 1002
rect 15725 929 16033 968
rect 15725 895 15733 929
rect 15767 895 15819 929
rect 15853 895 15905 929
rect 15939 895 15991 929
rect 16025 895 16033 929
rect 15725 856 16033 895
rect 15725 822 15733 856
rect 15767 822 15819 856
rect 15853 822 15905 856
rect 15939 822 15991 856
rect 16025 822 16033 856
rect 15725 783 16033 822
rect 15725 749 15733 783
rect 15767 749 15819 783
rect 15853 749 15905 783
rect 15939 749 15991 783
rect 16025 749 16033 783
rect 15725 710 16033 749
tri 15305 701 15314 710 se
rect 15314 701 15379 710
tri 15379 701 15388 710 nw
tri 15525 701 15534 710 se
rect 15534 701 15591 710
rect 12870 698 13222 701
tri 13222 698 13225 701 sw
tri 13849 698 13852 701 se
rect 13852 698 15376 701
tri 15376 698 15379 701 nw
tri 15522 698 15525 701 se
rect 15525 698 15591 701
rect 12870 692 15354 698
rect 12870 658 12882 692
rect 12916 658 12954 692
rect 12988 676 15354 692
tri 15354 676 15376 698 nw
tri 15517 693 15522 698 se
rect 15522 693 15591 698
tri 15591 693 15608 710 nw
tri 15500 676 15517 693 se
rect 15517 676 15574 693
tri 15574 676 15591 693 nw
rect 15725 676 15733 710
rect 15767 676 15819 710
rect 15853 676 15905 710
rect 15939 676 15991 710
rect 16025 676 16033 710
rect 12988 658 15327 676
rect 12870 649 15327 658
tri 15327 649 15354 676 nw
tri 15473 649 15500 676 se
rect 15500 649 15535 676
tri 15461 637 15473 649 se
rect 15473 637 15535 649
tri 15535 637 15574 676 nw
rect 15725 637 16033 676
tri 15443 619 15461 637 se
rect 15461 619 15517 637
tri 15517 619 15535 637 nw
tri 15427 603 15443 619 se
rect 15443 603 15501 619
tri 15501 603 15517 619 nw
rect 15725 603 15733 637
rect 15767 603 15819 637
rect 15853 603 15905 637
rect 15939 603 15991 637
rect 16025 603 16033 637
tri 15388 564 15427 603 se
rect 15427 564 15462 603
tri 15462 564 15501 603 nw
rect 15725 564 16033 603
tri 10960 547 10977 564 se
rect 10977 547 11114 564
tri 15371 547 15388 564 se
rect 15388 547 15445 564
tri 15445 547 15462 564 nw
rect 10783 495 10789 547
rect 10841 495 10853 547
rect 10905 495 10928 547
rect 10929 496 10930 546
rect 10958 496 10959 546
rect 10960 495 11114 547
rect 12870 538 15428 547
rect 12870 504 12882 538
rect 12916 504 12954 538
rect 12988 530 15428 538
tri 15428 530 15445 547 nw
rect 15725 530 15733 564
rect 15767 530 15819 564
rect 15853 530 15905 564
rect 15939 530 15991 564
rect 16025 530 16033 564
rect 12988 522 15420 530
tri 15420 522 15428 530 nw
rect 12988 504 15397 522
rect 12870 499 15397 504
tri 15397 499 15420 522 nw
tri 15702 499 15725 522 se
rect 15725 499 16033 530
rect 12870 495 13132 499
tri 13132 495 13136 499 nw
tri 13998 495 14002 499 ne
rect 14002 495 15393 499
tri 15393 495 15397 499 nw
tri 15698 495 15702 499 se
rect 15702 495 16033 499
tri 10960 491 10964 495 ne
rect 10964 491 11114 495
tri 15694 491 15698 495 se
rect 15698 491 16033 495
tri 10964 469 10986 491 ne
rect 6480 426 6481 452
rect 6482 425 6536 453
rect 6537 426 6538 452
tri 6479 418 6480 419 se
rect 6480 418 6538 425
tri 6538 418 6539 419 sw
tri 6454 393 6479 418 se
rect 6479 393 6539 418
tri 6539 393 6564 418 sw
rect 6445 341 6451 393
rect 6503 341 6515 393
rect 6567 341 6573 393
tri 10960 239 10986 265 se
rect 10986 239 11114 491
tri 15673 470 15694 491 se
rect 15694 470 15733 491
rect 13156 418 13162 470
rect 13214 418 13232 470
rect 13284 418 13302 470
rect 13354 418 13372 470
rect 13424 418 13442 470
rect 13494 418 13511 470
rect 13563 461 13580 470
rect 13632 461 13649 470
rect 13701 461 13718 470
rect 13770 461 13787 470
rect 13839 461 13856 470
rect 13908 461 13925 470
rect 13977 467 13983 470
tri 13983 467 13986 470 sw
tri 15670 467 15673 470 se
rect 15673 467 15733 470
rect 13977 461 15733 467
rect 13567 427 13580 461
rect 13640 427 13649 461
rect 13713 427 13718 461
rect 13786 427 13787 461
rect 14005 427 14044 461
rect 14078 427 14117 461
rect 14151 427 14190 461
rect 14224 427 14263 461
rect 14297 427 14336 461
rect 14370 427 14409 461
rect 14443 427 14482 461
rect 14516 427 14555 461
rect 14589 427 14628 461
rect 14662 427 14701 461
rect 14735 427 14774 461
rect 14808 427 14847 461
rect 14881 427 14920 461
rect 14954 427 14993 461
rect 15027 427 15065 461
rect 15099 427 15137 461
rect 15171 427 15209 461
rect 15243 427 15281 461
rect 15315 427 15353 461
rect 15387 427 15425 461
rect 15459 427 15497 461
rect 15531 427 15569 461
rect 15603 427 15641 461
rect 15675 457 15733 461
rect 15767 457 15819 491
rect 15853 457 15905 491
rect 15939 457 15991 491
rect 16025 457 16033 491
rect 15675 427 16033 457
rect 13563 418 13580 427
rect 13632 418 13649 427
rect 13701 418 13718 427
rect 13770 418 13787 427
rect 13839 418 13856 427
rect 13908 418 13925 427
rect 13977 421 16033 427
rect 13977 418 13983 421
tri 13983 418 13986 421 nw
tri 15670 418 15673 421 ne
rect 15673 418 16033 421
tri 15673 393 15698 418 ne
rect 15698 393 15733 418
rect 12867 390 13101 393
tri 13101 390 13104 393 sw
tri 14030 390 14033 393 se
rect 14033 390 15005 393
rect 12867 384 15005 390
rect 12867 350 12882 384
rect 12916 350 12954 384
rect 12988 350 15005 384
rect 12867 341 15005 350
rect 15057 341 15069 393
rect 15121 341 15127 393
tri 15698 384 15707 393 ne
rect 15707 384 15733 393
rect 15767 384 15819 418
rect 15853 384 15905 418
rect 15939 384 15991 418
rect 16025 384 16033 418
tri 15707 366 15725 384 ne
rect 15725 345 16033 384
rect 15725 311 15733 345
rect 15767 311 15819 345
rect 15853 311 15905 345
rect 15939 311 15991 345
rect 16025 311 16033 345
rect 15725 272 16033 311
rect 348 188 406 226
rect 348 154 360 188
rect 394 154 406 188
rect 466 187 473 239
rect 525 187 537 239
rect 589 187 596 239
rect 3203 187 3209 239
rect 3261 187 3273 239
rect 3325 187 3333 239
rect 3334 188 3335 238
rect 3363 188 3364 238
rect 3365 230 3498 239
rect 3365 196 3380 230
rect 3414 196 3452 230
rect 3486 196 3498 230
rect 3365 187 3498 196
rect 5142 187 5149 239
rect 5201 187 5213 239
rect 5265 187 5272 239
rect 10783 187 10789 239
rect 10841 187 10853 239
rect 10905 187 10928 239
rect 10929 188 10930 238
rect 10958 188 10959 238
rect 10960 233 11114 239
rect 10960 230 11111 233
tri 11111 230 11114 233 nw
rect 12870 230 15173 239
rect 10960 196 11077 230
tri 11077 196 11111 230 nw
rect 12870 196 12882 230
rect 12916 196 12954 230
rect 12988 196 15173 230
rect 10960 187 11068 196
tri 11068 187 11077 196 nw
rect 12870 187 15173 196
rect 15225 187 15237 239
rect 15289 187 15295 239
rect 15725 238 15733 272
rect 15767 238 15819 272
rect 15853 238 15905 272
rect 15939 238 15991 272
rect 16025 238 16033 272
rect 15725 199 16033 238
rect 348 126 406 154
rect 15725 165 15733 199
rect 15767 165 15819 199
rect 15853 165 15905 199
rect 15939 165 15991 199
rect 16025 165 16033 199
tri 406 126 425 145 sw
tri 15718 126 15725 133 se
rect 15725 126 16033 165
rect 348 93 425 126
tri 425 93 458 126 sw
tri 15685 93 15718 126 se
rect 15718 93 15733 126
rect 348 41 363 93
rect 415 84 427 93
rect 479 84 491 93
rect 543 84 555 93
rect 607 84 619 93
rect 671 84 683 93
rect 423 50 427 84
rect 671 50 677 84
rect 415 41 427 50
rect 479 41 491 50
rect 543 41 555 50
rect 607 41 619 50
rect 671 41 683 50
rect 735 41 886 93
rect 938 84 950 93
rect 1002 84 1014 93
rect 1066 84 1078 93
rect 1130 84 1142 93
rect 1194 84 1206 93
rect 949 50 950 84
rect 1130 50 1131 84
rect 1194 50 1203 84
rect 938 41 950 50
rect 1002 41 1014 50
rect 1066 41 1078 50
rect 1130 41 1142 50
rect 1194 41 1206 50
rect 1258 41 1270 93
rect 1322 41 1334 93
rect 1386 41 1398 93
rect 1450 84 1462 93
rect 1514 84 1526 93
rect 1578 84 1590 93
rect 1642 84 1654 93
rect 1706 84 1718 93
rect 1770 84 1782 93
rect 1453 50 1462 84
rect 1525 50 1526 84
rect 1706 50 1707 84
rect 1770 50 1779 84
rect 1450 41 1462 50
rect 1514 41 1526 50
rect 1578 41 1590 50
rect 1642 41 1654 50
rect 1706 41 1718 50
rect 1770 41 1782 50
rect 1834 41 1846 93
rect 1898 41 1910 93
rect 1962 41 1974 93
rect 2026 84 2038 93
rect 2090 84 2102 93
rect 2154 84 2166 93
rect 2218 84 2230 93
rect 2282 84 2294 93
rect 2346 84 2358 93
rect 2029 50 2038 84
rect 2101 50 2102 84
rect 2282 50 2283 84
rect 2346 50 2355 84
rect 2026 41 2038 50
rect 2090 41 2102 50
rect 2154 41 2166 50
rect 2218 41 2230 50
rect 2282 41 2294 50
rect 2346 41 2358 50
rect 2410 41 2422 93
rect 2474 41 2486 93
rect 2538 41 2550 93
rect 2602 84 2614 93
rect 2666 84 2678 93
rect 2730 84 2742 93
rect 2794 84 2806 93
rect 2858 84 2870 93
rect 2922 84 2934 93
rect 2605 50 2614 84
rect 2677 50 2678 84
rect 2858 50 2859 84
rect 2922 50 2931 84
rect 2602 41 2614 50
rect 2666 41 2678 50
rect 2730 41 2742 50
rect 2794 41 2806 50
rect 2858 41 2870 50
rect 2922 41 2934 50
rect 2986 41 2998 93
rect 3050 41 3062 93
rect 3114 41 3126 93
rect 3178 84 3190 93
rect 3242 84 3254 93
rect 3306 84 3318 93
rect 3370 84 3382 93
rect 3434 84 3446 93
rect 3498 84 3510 93
rect 3181 50 3190 84
rect 3253 50 3254 84
rect 3434 50 3435 84
rect 3498 50 3507 84
rect 3178 41 3190 50
rect 3242 41 3254 50
rect 3306 41 3318 50
rect 3370 41 3382 50
rect 3434 41 3446 50
rect 3498 41 3510 50
rect 3562 41 3574 93
rect 3626 41 3638 93
rect 3690 41 3702 93
rect 3754 84 3766 93
rect 3818 84 3830 93
rect 3882 84 3894 93
rect 3946 84 3958 93
rect 4010 84 4022 93
rect 4074 84 4086 93
rect 3757 50 3766 84
rect 3829 50 3830 84
rect 4010 50 4011 84
rect 4074 50 4083 84
rect 3754 41 3766 50
rect 3818 41 3830 50
rect 3882 41 3894 50
rect 3946 41 3958 50
rect 4010 41 4022 50
rect 4074 41 4086 50
rect 4138 41 4150 93
rect 4202 41 4214 93
rect 4266 41 4278 93
rect 4330 84 4342 93
rect 4394 84 4406 93
rect 4458 84 4470 93
rect 4522 84 4534 93
rect 4586 84 4598 93
rect 4650 84 4662 93
rect 4333 50 4342 84
rect 4405 50 4406 84
rect 4586 50 4587 84
rect 4650 50 4659 84
rect 4330 41 4342 50
rect 4394 41 4406 50
rect 4458 41 4470 50
rect 4522 41 4534 50
rect 4586 41 4598 50
rect 4650 41 4662 50
rect 4714 41 4726 93
rect 4778 41 4790 93
rect 4842 41 4854 93
rect 4906 84 4918 93
rect 4970 84 4982 93
rect 5034 84 5046 93
rect 5098 84 5110 93
rect 5162 84 5174 93
rect 5226 84 5238 93
rect 4909 50 4918 84
rect 4981 50 4982 84
rect 5162 50 5163 84
rect 5226 50 5235 84
rect 4906 41 4918 50
rect 4970 41 4982 50
rect 5034 41 5046 50
rect 5098 41 5110 50
rect 5162 41 5174 50
rect 5226 41 5238 50
rect 5290 41 5302 93
rect 5354 41 5366 93
rect 5418 41 5430 93
rect 5482 84 5494 93
rect 5546 84 5558 93
rect 5610 84 5622 93
rect 5674 84 5686 93
rect 5738 84 5750 93
rect 5802 84 5814 93
rect 5485 50 5494 84
rect 5557 50 5558 84
rect 5738 50 5739 84
rect 5802 50 5811 84
rect 5482 41 5494 50
rect 5546 41 5558 50
rect 5610 41 5622 50
rect 5674 41 5686 50
rect 5738 41 5750 50
rect 5802 41 5814 50
rect 5866 41 5878 93
rect 5930 41 5942 93
rect 5994 41 6006 93
rect 6058 84 6070 93
rect 6122 84 6134 93
rect 6186 84 6198 93
rect 6250 84 6262 93
rect 6314 84 6326 93
rect 6378 84 6390 93
rect 6061 50 6070 84
rect 6133 50 6134 84
rect 6314 50 6315 84
rect 6378 50 6387 84
rect 6058 41 6070 50
rect 6122 41 6134 50
rect 6186 41 6198 50
rect 6250 41 6262 50
rect 6314 41 6326 50
rect 6378 41 6390 50
rect 6442 41 6454 93
rect 6506 41 6518 93
rect 6570 41 6582 93
rect 6634 84 6646 93
rect 6698 84 6710 93
rect 6762 84 6774 93
rect 6826 84 6838 93
rect 6890 84 6902 93
rect 6954 84 6966 93
rect 6637 50 6646 84
rect 6709 50 6710 84
rect 6890 50 6891 84
rect 6954 50 6963 84
rect 6634 41 6646 50
rect 6698 41 6710 50
rect 6762 41 6774 50
rect 6826 41 6838 50
rect 6890 41 6902 50
rect 6954 41 6966 50
rect 7018 41 7030 93
rect 7082 41 7094 93
rect 7146 41 7158 93
rect 7210 84 7222 93
rect 7274 84 7286 93
rect 7338 84 7350 93
rect 7402 84 7414 93
rect 7466 84 7478 93
rect 7530 84 7542 93
rect 7213 50 7222 84
rect 7285 50 7286 84
rect 7466 50 7467 84
rect 7530 50 7539 84
rect 7210 41 7222 50
rect 7274 41 7286 50
rect 7338 41 7350 50
rect 7402 41 7414 50
rect 7466 41 7478 50
rect 7530 41 7542 50
rect 7594 41 7606 93
rect 7658 41 7670 93
rect 7722 41 7734 93
rect 7786 84 7798 93
rect 7850 84 7862 93
rect 7914 84 7926 93
rect 7978 84 7990 93
rect 8042 84 8054 93
rect 8106 84 8118 93
rect 7789 50 7798 84
rect 7861 50 7862 84
rect 8042 50 8043 84
rect 8106 50 8115 84
rect 7786 41 7798 50
rect 7850 41 7862 50
rect 7914 41 7926 50
rect 7978 41 7990 50
rect 8042 41 8054 50
rect 8106 41 8118 50
rect 8170 41 8182 93
rect 8234 41 8246 93
rect 8298 41 8310 93
rect 8362 84 8374 93
rect 8426 84 8438 93
rect 8490 84 8502 93
rect 8554 84 8566 93
rect 8618 84 8630 93
rect 8682 84 8694 93
rect 8365 50 8374 84
rect 8437 50 8438 84
rect 8618 50 8619 84
rect 8682 50 8691 84
rect 8362 41 8374 50
rect 8426 41 8438 50
rect 8490 41 8502 50
rect 8554 41 8566 50
rect 8618 41 8630 50
rect 8682 41 8694 50
rect 8746 41 8758 93
rect 8810 41 8822 93
rect 8874 41 8886 93
rect 8938 84 8950 93
rect 9002 84 9014 93
rect 9066 84 9078 93
rect 9130 84 9142 93
rect 9194 84 9206 93
rect 9258 84 9270 93
rect 8941 50 8950 84
rect 9013 50 9014 84
rect 9194 50 9195 84
rect 9258 50 9267 84
rect 8938 41 8950 50
rect 9002 41 9014 50
rect 9066 41 9078 50
rect 9130 41 9142 50
rect 9194 41 9206 50
rect 9258 41 9270 50
rect 9322 41 9334 93
rect 9386 41 9398 93
rect 9450 41 9462 93
rect 9514 84 9526 93
rect 9578 84 9590 93
rect 9642 84 9654 93
rect 9706 84 9718 93
rect 9770 84 9782 93
rect 9834 84 9846 93
rect 9517 50 9526 84
rect 9589 50 9590 84
rect 9770 50 9771 84
rect 9834 50 9843 84
rect 9514 41 9526 50
rect 9578 41 9590 50
rect 9642 41 9654 50
rect 9706 41 9718 50
rect 9770 41 9782 50
rect 9834 41 9846 50
rect 9898 41 9910 93
rect 9962 41 9974 93
rect 10026 41 10038 93
rect 10090 84 10102 93
rect 10154 84 10166 93
rect 10218 84 10230 93
rect 10282 84 10294 93
rect 10346 84 10358 93
rect 10410 84 10422 93
rect 10093 50 10102 84
rect 10165 50 10166 84
rect 10346 50 10347 84
rect 10410 50 10419 84
rect 10090 41 10102 50
rect 10154 41 10166 50
rect 10218 41 10230 50
rect 10282 41 10294 50
rect 10346 41 10358 50
rect 10410 41 10422 50
rect 10474 41 10486 93
rect 10538 41 10550 93
rect 10602 41 10614 93
rect 10666 84 10678 93
rect 10730 84 10742 93
rect 10794 84 10806 93
rect 10858 84 10870 93
rect 10922 84 10934 93
rect 10986 84 10998 93
rect 10669 50 10678 84
rect 10741 50 10742 84
rect 10922 50 10923 84
rect 10986 50 10995 84
rect 10666 41 10678 50
rect 10730 41 10742 50
rect 10794 41 10806 50
rect 10858 41 10870 50
rect 10922 41 10934 50
rect 10986 41 10998 50
rect 11050 41 11062 93
rect 11114 41 11126 93
rect 11178 41 11190 93
rect 11242 84 11254 93
rect 11306 84 11318 93
rect 11370 84 11382 93
rect 11434 84 11446 93
rect 11498 84 11510 93
rect 11562 84 11574 93
rect 11245 50 11254 84
rect 11317 50 11318 84
rect 11498 50 11499 84
rect 11562 50 11571 84
rect 11242 41 11254 50
rect 11306 41 11318 50
rect 11370 41 11382 50
rect 11434 41 11446 50
rect 11498 41 11510 50
rect 11562 41 11574 50
rect 11626 41 11638 93
rect 11690 41 11702 93
rect 11754 41 11766 93
rect 11818 84 11830 93
rect 11882 84 11894 93
rect 11946 84 11958 93
rect 12010 84 12022 93
rect 12074 84 12086 93
rect 12138 84 12150 93
rect 11821 50 11830 84
rect 11893 50 11894 84
rect 12074 50 12075 84
rect 12138 50 12147 84
rect 11818 41 11830 50
rect 11882 41 11894 50
rect 11946 41 11958 50
rect 12010 41 12022 50
rect 12074 41 12086 50
rect 12138 41 12150 50
rect 12202 41 12214 93
rect 12266 41 12278 93
rect 12330 41 12342 93
rect 12394 84 12406 93
rect 12458 84 12470 93
rect 12522 84 12534 93
rect 12586 84 12598 93
rect 12650 84 12662 93
rect 12714 84 12726 93
rect 12397 50 12406 84
rect 12469 50 12470 84
rect 12650 50 12651 84
rect 12714 50 12723 84
rect 12394 41 12406 50
rect 12458 41 12470 50
rect 12522 41 12534 50
rect 12586 41 12598 50
rect 12650 41 12662 50
rect 12714 41 12726 50
rect 12778 41 12790 93
rect 12842 41 12854 93
rect 12906 41 12918 93
rect 12970 84 12982 93
rect 13034 84 13046 93
rect 13098 84 13110 93
rect 13162 84 13174 93
rect 13226 84 13238 93
rect 13290 84 13302 93
rect 12973 50 12982 84
rect 13045 50 13046 84
rect 13226 50 13227 84
rect 13290 50 13299 84
rect 12970 41 12982 50
rect 13034 41 13046 50
rect 13098 41 13110 50
rect 13162 41 13174 50
rect 13226 41 13238 50
rect 13290 41 13302 50
rect 13354 41 13366 93
rect 13418 41 13430 93
rect 13482 41 13494 93
rect 13546 84 13558 93
rect 13610 84 13622 93
rect 13674 84 13686 93
rect 13738 84 13750 93
rect 13802 84 13814 93
rect 13866 84 13878 93
rect 13549 50 13558 84
rect 13621 50 13622 84
rect 13802 50 13803 84
rect 13866 50 13875 84
rect 13546 41 13558 50
rect 13610 41 13622 50
rect 13674 41 13686 50
rect 13738 41 13750 50
rect 13802 41 13814 50
rect 13866 41 13878 50
rect 13930 41 13942 93
rect 13994 41 14006 93
rect 14058 41 14070 93
rect 14122 84 14134 93
rect 14186 84 14198 93
rect 14250 84 14262 93
rect 14314 84 14326 93
rect 14125 50 14134 84
rect 14197 50 14198 84
rect 14122 41 14134 50
rect 14186 41 14198 50
rect 14250 41 14262 50
rect 14314 41 14326 50
rect 14378 41 14384 93
tri 15684 92 15685 93 se
rect 15685 92 15733 93
rect 15767 92 15819 126
rect 15853 92 15905 126
rect 15939 92 15991 126
rect 16025 92 16033 126
tri 15645 53 15684 92 se
rect 15684 53 16033 92
tri 15633 41 15645 53 se
rect 15645 41 15733 53
tri 15611 19 15633 41 se
rect 15633 19 15733 41
rect 15767 19 15819 53
rect 15853 19 15905 53
rect 15939 19 15991 53
rect 16025 19 16033 53
tri 15576 -16 15611 19 se
rect 15611 -13 16033 19
rect 15611 -16 15726 -13
<< rmetal1 >>
rect 3333 7881 3335 7882
rect 3333 7831 3334 7881
rect 3333 7830 3335 7831
rect 3363 7881 3365 7882
rect 3364 7831 3365 7881
rect 3363 7830 3365 7831
rect 3337 7727 3338 7728
rect 3364 7727 3365 7728
rect 3337 7726 3365 7727
rect 3337 7677 3365 7678
rect 3337 7676 3338 7677
rect 3364 7676 3365 7677
rect 3333 7573 3335 7574
rect 3333 7523 3334 7573
rect 3333 7522 3335 7523
rect 3363 7573 3365 7574
rect 3364 7523 3365 7573
rect 3363 7522 3365 7523
rect 3337 7419 3338 7420
rect 3364 7419 3365 7420
rect 3337 7418 3365 7419
rect 3337 7369 3365 7370
rect 3337 7368 3338 7369
rect 3364 7368 3365 7369
rect 3333 7265 3335 7266
rect 3333 7215 3334 7265
rect 3333 7214 3335 7215
rect 3363 7265 3365 7266
rect 3364 7215 3365 7265
rect 3363 7214 3365 7215
rect 3337 7111 3338 7112
rect 3364 7111 3365 7112
rect 3337 7110 3365 7111
rect 3337 7061 3365 7062
rect 3337 7060 3338 7061
rect 3364 7060 3365 7061
rect 3333 6957 3335 6958
rect 3333 6907 3334 6957
rect 3333 6906 3335 6907
rect 3363 6957 3365 6958
rect 3364 6907 3365 6957
rect 3363 6906 3365 6907
rect 3337 6803 3338 6804
rect 3364 6803 3365 6804
rect 3337 6802 3365 6803
rect 3337 6753 3365 6754
rect 3337 6752 3338 6753
rect 3364 6752 3365 6753
rect 3333 6649 3335 6650
rect 3333 6599 3334 6649
rect 3333 6598 3335 6599
rect 3363 6649 3365 6650
rect 3364 6599 3365 6649
rect 3363 6598 3365 6599
rect 3337 6495 3338 6496
rect 3364 6495 3365 6496
rect 3337 6494 3365 6495
rect 3337 6445 3365 6446
rect 3337 6444 3338 6445
rect 3364 6444 3365 6445
rect 3333 6341 3335 6342
rect 3333 6291 3334 6341
rect 3333 6290 3335 6291
rect 3363 6341 3365 6342
rect 3364 6291 3365 6341
rect 3363 6290 3365 6291
rect 3337 6187 3338 6188
rect 3364 6187 3365 6188
rect 3337 6186 3365 6187
rect 3337 6137 3365 6138
rect 3337 6136 3338 6137
rect 3364 6136 3365 6137
rect 1344 1990 1402 1991
rect 1344 1989 1345 1990
rect 1401 1989 1402 1990
rect 1344 1960 1345 1961
rect 1401 1960 1402 1961
rect 1344 1959 1402 1960
rect 466 1690 468 1691
rect 467 1664 468 1690
rect 466 1663 468 1664
rect 594 1690 596 1691
rect 594 1664 595 1690
rect 594 1663 596 1664
rect 2200 1682 2258 1683
rect 2200 1681 2201 1682
rect 2257 1681 2258 1682
rect 2200 1652 2201 1653
rect 2257 1652 2258 1653
rect 2200 1651 2258 1652
rect 466 1385 596 1386
rect 466 1384 467 1385
rect 595 1384 596 1385
rect 466 1355 467 1356
rect 595 1355 596 1356
rect 466 1354 596 1355
rect 3337 1932 3338 1933
rect 3364 1932 3365 1933
rect 3337 1931 3365 1932
rect 3337 1882 3365 1883
rect 3337 1881 3338 1882
rect 3364 1881 3365 1882
rect 3333 1778 3335 1779
rect 3333 1728 3334 1778
rect 3333 1727 3335 1728
rect 3363 1778 3365 1779
rect 3364 1728 3365 1778
rect 3363 1727 3365 1728
rect 3337 1624 3338 1625
rect 3364 1624 3365 1625
rect 3337 1623 3365 1624
rect 3337 1574 3365 1575
rect 3337 1573 3338 1574
rect 3364 1573 3365 1574
rect 3333 1470 3335 1471
rect 3333 1420 3334 1470
rect 3333 1419 3335 1420
rect 3363 1470 3365 1471
rect 3364 1420 3365 1470
rect 3363 1419 3365 1420
rect 3056 1376 3058 1377
rect 3057 1350 3058 1376
rect 3056 1349 3058 1350
rect 3112 1376 3114 1377
rect 3112 1350 3113 1376
rect 3112 1349 3114 1350
rect 3337 1316 3338 1317
rect 3364 1316 3365 1317
rect 3337 1315 3365 1316
rect 3337 1266 3365 1267
rect 3337 1265 3338 1266
rect 3364 1265 3365 1266
rect 3333 1162 3335 1163
rect 3333 1112 3334 1162
rect 3333 1111 3335 1112
rect 3363 1162 3365 1163
rect 3364 1112 3365 1162
rect 3363 1111 3365 1112
rect 466 1077 596 1078
rect 466 1076 467 1077
rect 595 1076 596 1077
rect 466 1047 467 1048
rect 595 1047 596 1048
rect 466 1046 596 1047
rect 3337 1008 3338 1009
rect 3364 1008 3365 1009
rect 3337 1007 3365 1008
rect 3337 958 3365 959
rect 3337 957 3338 958
rect 3364 957 3365 958
rect 3333 854 3335 855
rect 3333 804 3334 854
rect 3333 803 3335 804
rect 3363 854 3365 855
rect 3364 804 3365 854
rect 3363 803 3365 804
rect 466 770 596 771
rect 466 769 467 770
rect 595 769 596 770
rect 466 740 467 741
rect 595 740 596 741
rect 466 739 596 740
rect 3337 700 3338 701
rect 3364 700 3365 701
rect 3337 699 3365 700
rect 3337 650 3365 651
rect 3337 649 3338 650
rect 3364 649 3365 650
rect 4768 1068 4770 1069
rect 4769 1042 4770 1068
rect 4768 1041 4770 1042
rect 4824 1068 4826 1069
rect 4824 1042 4825 1068
rect 4824 1041 4826 1042
rect 3333 546 3335 547
rect 3333 496 3334 546
rect 3333 495 3335 496
rect 3363 546 3365 547
rect 3364 496 3365 546
rect 3363 495 3365 496
rect 466 462 596 463
rect 466 461 467 462
rect 595 461 596 462
rect 466 432 467 433
rect 595 432 596 433
rect 466 431 596 432
rect 3337 392 3338 393
rect 3364 392 3365 393
rect 3337 391 3365 392
rect 3337 342 3365 343
rect 3337 341 3338 342
rect 3364 341 3365 342
rect 5938 1932 5939 1933
rect 5965 1932 5966 1933
rect 5938 1931 5966 1932
rect 5938 1882 5966 1883
rect 5938 1881 5939 1882
rect 5965 1881 5966 1882
rect 5624 760 5626 761
rect 5625 734 5626 760
rect 5624 733 5626 734
rect 5680 760 5682 761
rect 5680 734 5681 760
rect 5680 733 5682 734
rect 14298 5896 14300 5897
rect 14298 5846 14299 5896
rect 14298 5845 14300 5846
rect 14328 5896 14330 5897
rect 14329 5846 14330 5896
rect 14328 5845 14330 5846
rect 14479 5896 14481 5897
rect 14479 5846 14480 5896
rect 14479 5845 14481 5846
rect 14509 5896 14511 5897
rect 14510 5846 14511 5896
rect 14509 5845 14511 5846
rect 11612 5809 11742 5810
rect 11612 5808 11613 5809
rect 11741 5808 11742 5809
rect 11612 5779 11613 5780
rect 11741 5779 11742 5780
rect 11612 5778 11742 5779
rect 14483 5742 14484 5743
rect 14510 5742 14511 5743
rect 14483 5741 14511 5742
rect 14483 5692 14511 5693
rect 14483 5691 14484 5692
rect 14510 5691 14511 5692
rect 14479 5588 14481 5589
rect 14479 5538 14480 5588
rect 14479 5537 14481 5538
rect 14509 5588 14511 5589
rect 14510 5538 14511 5588
rect 14509 5537 14511 5538
rect 11612 5501 11742 5502
rect 11612 5500 11613 5501
rect 11741 5500 11742 5501
rect 11612 5471 11613 5472
rect 11741 5471 11742 5472
rect 11612 5470 11742 5471
rect 14483 5434 14484 5435
rect 14510 5434 14511 5435
rect 14483 5433 14511 5434
rect 14483 5384 14511 5385
rect 14483 5383 14484 5384
rect 14510 5383 14511 5384
rect 14479 5280 14481 5281
rect 14479 5230 14480 5280
rect 14479 5229 14481 5230
rect 14509 5280 14511 5281
rect 14510 5230 14511 5280
rect 14509 5229 14511 5230
rect 11612 5195 11614 5196
rect 11613 5169 11614 5195
rect 11612 5168 11614 5169
rect 11740 5195 11742 5196
rect 11740 5169 11741 5195
rect 11740 5168 11742 5169
rect 14483 5126 14484 5127
rect 14510 5126 14511 5127
rect 14483 5125 14511 5126
rect 14483 5076 14511 5077
rect 14483 5075 14484 5076
rect 14510 5075 14511 5076
rect 14479 4972 14481 4973
rect 14479 4922 14480 4972
rect 14479 4921 14481 4922
rect 14509 4972 14511 4973
rect 14510 4922 14511 4972
rect 14509 4921 14511 4922
rect 11612 4885 11742 4886
rect 11612 4884 11613 4885
rect 11741 4884 11742 4885
rect 11612 4855 11613 4856
rect 11741 4855 11742 4856
rect 11612 4854 11742 4855
rect 14483 4818 14484 4819
rect 14510 4818 14511 4819
rect 14483 4817 14511 4818
rect 14483 4768 14511 4769
rect 14483 4767 14484 4768
rect 14510 4767 14511 4768
rect 14479 4664 14481 4665
rect 14479 4614 14480 4664
rect 14479 4613 14481 4614
rect 14509 4664 14511 4665
rect 14510 4614 14511 4664
rect 14509 4613 14511 4614
rect 11612 4577 11742 4578
rect 11612 4576 11613 4577
rect 11741 4576 11742 4577
rect 11612 4547 11613 4548
rect 11741 4547 11742 4548
rect 11612 4546 11742 4547
rect 14483 4510 14484 4511
rect 14510 4510 14511 4511
rect 14483 4509 14511 4510
rect 14483 4460 14511 4461
rect 14483 4459 14484 4460
rect 14510 4459 14511 4460
rect 14479 4356 14481 4357
rect 14479 4306 14480 4356
rect 14479 4305 14481 4306
rect 14509 4356 14511 4357
rect 14510 4306 14511 4356
rect 14509 4305 14511 4306
rect 14483 4202 14484 4203
rect 14510 4202 14511 4203
rect 14483 4201 14511 4202
rect 14483 4152 14511 4153
rect 14483 4151 14484 4152
rect 14510 4151 14511 4152
rect 14483 3916 14484 3917
rect 14510 3916 14511 3917
rect 14483 3915 14511 3916
rect 14483 3866 14511 3867
rect 14483 3865 14484 3866
rect 14510 3865 14511 3866
rect 14479 3762 14481 3763
rect 14479 3712 14480 3762
rect 14479 3711 14481 3712
rect 14509 3762 14511 3763
rect 14510 3712 14511 3762
rect 14509 3711 14511 3712
rect 14483 3608 14484 3609
rect 14510 3608 14511 3609
rect 14483 3607 14511 3608
rect 14483 3558 14511 3559
rect 14483 3557 14484 3558
rect 14510 3557 14511 3558
rect 14479 3454 14481 3455
rect 14479 3404 14480 3454
rect 14479 3403 14481 3404
rect 14509 3454 14511 3455
rect 14510 3404 14511 3454
rect 14509 3403 14511 3404
rect 14483 3300 14484 3301
rect 14510 3300 14511 3301
rect 14483 3299 14511 3300
rect 14483 3250 14511 3251
rect 14483 3249 14484 3250
rect 14510 3249 14511 3250
rect 14479 3146 14481 3147
rect 14479 3096 14480 3146
rect 14479 3095 14481 3096
rect 14509 3146 14511 3147
rect 14510 3096 14511 3146
rect 14509 3095 14511 3096
rect 14483 2992 14484 2993
rect 14510 2992 14511 2993
rect 14483 2991 14511 2992
rect 14483 2942 14511 2943
rect 14483 2941 14484 2942
rect 14510 2941 14511 2942
rect 14479 2838 14481 2839
rect 14479 2788 14480 2838
rect 14479 2787 14481 2788
rect 14509 2838 14511 2839
rect 14510 2788 14511 2838
rect 14509 2787 14511 2788
rect 14483 2684 14484 2685
rect 14510 2684 14511 2685
rect 14483 2683 14511 2684
rect 14483 2634 14511 2635
rect 14483 2633 14484 2634
rect 14510 2633 14511 2634
rect 14479 2530 14481 2531
rect 14479 2480 14480 2530
rect 14479 2479 14481 2480
rect 14509 2530 14511 2531
rect 14510 2480 14511 2530
rect 14509 2479 14511 2480
rect 14483 2376 14484 2377
rect 14510 2376 14511 2377
rect 14483 2375 14511 2376
rect 14483 2326 14511 2327
rect 14483 2325 14484 2326
rect 14510 2325 14511 2326
rect 14479 2222 14481 2223
rect 14479 2172 14480 2222
rect 14479 2171 14481 2172
rect 14509 2222 14511 2223
rect 14510 2172 14511 2222
rect 14509 2171 14511 2172
rect 10928 1778 10930 1779
rect 10928 1728 10929 1778
rect 10928 1727 10930 1728
rect 10958 1778 10960 1779
rect 10959 1728 10960 1778
rect 10958 1727 10960 1728
rect 10926 1470 10927 1471
rect 10953 1470 10954 1471
rect 10926 1469 10954 1470
rect 10926 1420 10954 1421
rect 10926 1419 10927 1420
rect 10953 1419 10954 1420
rect 10928 1162 10930 1163
rect 10928 1112 10929 1162
rect 10928 1111 10930 1112
rect 10958 1162 10960 1163
rect 10959 1112 10960 1162
rect 10958 1111 10960 1112
rect 10928 854 10930 855
rect 10928 804 10929 854
rect 10928 803 10930 804
rect 10958 854 10960 855
rect 10959 804 10960 854
rect 10958 803 10960 804
rect 10928 546 10930 547
rect 10928 496 10929 546
rect 10928 495 10930 496
rect 10958 546 10960 547
rect 10959 496 10960 546
rect 10958 495 10960 496
rect 6480 452 6482 453
rect 6481 426 6482 452
rect 6480 425 6482 426
rect 6536 452 6538 453
rect 6536 426 6537 452
rect 6536 425 6538 426
rect 3333 238 3335 239
rect 3333 188 3334 238
rect 3333 187 3335 188
rect 3363 238 3365 239
rect 3364 188 3365 238
rect 3363 187 3365 188
rect 10928 238 10930 239
rect 10928 188 10929 238
rect 10928 187 10930 188
rect 10958 238 10960 239
rect 10959 188 10960 238
rect 10958 187 10960 188
<< via1 >>
rect 354 8000 406 8027
rect 354 7975 360 8000
rect 360 7975 394 8000
rect 394 7975 406 8000
rect 418 8018 470 8027
rect 482 8018 534 8027
rect 546 8018 598 8027
rect 610 8018 662 8027
rect 674 8018 726 8027
rect 857 8018 909 8027
rect 921 8018 973 8027
rect 985 8018 1037 8027
rect 1049 8018 1101 8027
rect 1113 8018 1165 8027
rect 1177 8018 1229 8027
rect 1241 8018 1293 8027
rect 418 7984 445 8018
rect 445 7984 470 8018
rect 482 7984 517 8018
rect 517 7984 534 8018
rect 546 7984 551 8018
rect 551 7984 589 8018
rect 589 7984 598 8018
rect 610 7984 623 8018
rect 623 7984 661 8018
rect 661 7984 662 8018
rect 674 7984 695 8018
rect 695 7984 726 8018
rect 857 7984 876 8018
rect 876 7984 909 8018
rect 921 7984 948 8018
rect 948 7984 973 8018
rect 985 7984 1020 8018
rect 1020 7984 1037 8018
rect 1049 7984 1054 8018
rect 1054 7984 1092 8018
rect 1092 7984 1101 8018
rect 1113 7984 1126 8018
rect 1126 7984 1164 8018
rect 1164 7984 1165 8018
rect 1177 7984 1198 8018
rect 1198 7984 1229 8018
rect 1241 7984 1270 8018
rect 1270 7984 1293 8018
rect 418 7975 470 7984
rect 482 7975 534 7984
rect 546 7975 598 7984
rect 610 7975 662 7984
rect 674 7975 726 7984
rect 857 7975 909 7984
rect 921 7975 973 7984
rect 985 7975 1037 7984
rect 1049 7975 1101 7984
rect 1113 7975 1165 7984
rect 1177 7975 1229 7984
rect 1241 7975 1293 7984
rect 1305 8018 1357 8027
rect 1305 7984 1308 8018
rect 1308 7984 1342 8018
rect 1342 7984 1357 8018
rect 1305 7975 1357 7984
rect 1369 8018 1421 8027
rect 1369 7984 1380 8018
rect 1380 7984 1414 8018
rect 1414 7984 1421 8018
rect 1369 7975 1421 7984
rect 1433 8018 1485 8027
rect 1497 8018 1549 8027
rect 1561 8018 1613 8027
rect 1625 8018 1677 8027
rect 1689 8018 1741 8027
rect 1753 8018 1805 8027
rect 1817 8018 1869 8027
rect 1433 7984 1452 8018
rect 1452 7984 1485 8018
rect 1497 7984 1524 8018
rect 1524 7984 1549 8018
rect 1561 7984 1596 8018
rect 1596 7984 1613 8018
rect 1625 7984 1630 8018
rect 1630 7984 1668 8018
rect 1668 7984 1677 8018
rect 1689 7984 1702 8018
rect 1702 7984 1740 8018
rect 1740 7984 1741 8018
rect 1753 7984 1774 8018
rect 1774 7984 1805 8018
rect 1817 7984 1846 8018
rect 1846 7984 1869 8018
rect 1433 7975 1485 7984
rect 1497 7975 1549 7984
rect 1561 7975 1613 7984
rect 1625 7975 1677 7984
rect 1689 7975 1741 7984
rect 1753 7975 1805 7984
rect 1817 7975 1869 7984
rect 1881 8018 1933 8027
rect 1881 7984 1884 8018
rect 1884 7984 1918 8018
rect 1918 7984 1933 8018
rect 1881 7975 1933 7984
rect 1945 8018 1997 8027
rect 1945 7984 1956 8018
rect 1956 7984 1990 8018
rect 1990 7984 1997 8018
rect 1945 7975 1997 7984
rect 2009 8018 2061 8027
rect 2073 8018 2125 8027
rect 2137 8018 2189 8027
rect 2201 8018 2253 8027
rect 2265 8018 2317 8027
rect 2329 8018 2381 8027
rect 2393 8018 2445 8027
rect 2009 7984 2028 8018
rect 2028 7984 2061 8018
rect 2073 7984 2100 8018
rect 2100 7984 2125 8018
rect 2137 7984 2172 8018
rect 2172 7984 2189 8018
rect 2201 7984 2206 8018
rect 2206 7984 2244 8018
rect 2244 7984 2253 8018
rect 2265 7984 2278 8018
rect 2278 7984 2316 8018
rect 2316 7984 2317 8018
rect 2329 7984 2350 8018
rect 2350 7984 2381 8018
rect 2393 7984 2422 8018
rect 2422 7984 2445 8018
rect 2009 7975 2061 7984
rect 2073 7975 2125 7984
rect 2137 7975 2189 7984
rect 2201 7975 2253 7984
rect 2265 7975 2317 7984
rect 2329 7975 2381 7984
rect 2393 7975 2445 7984
rect 2457 8018 2509 8027
rect 2457 7984 2460 8018
rect 2460 7984 2494 8018
rect 2494 7984 2509 8018
rect 2457 7975 2509 7984
rect 2521 8018 2573 8027
rect 2521 7984 2532 8018
rect 2532 7984 2566 8018
rect 2566 7984 2573 8018
rect 2521 7975 2573 7984
rect 2585 8018 2637 8027
rect 2649 8018 2701 8027
rect 2713 8018 2765 8027
rect 2777 8018 2829 8027
rect 2841 8018 2893 8027
rect 2905 8018 2957 8027
rect 2969 8018 3021 8027
rect 2585 7984 2604 8018
rect 2604 7984 2637 8018
rect 2649 7984 2676 8018
rect 2676 7984 2701 8018
rect 2713 7984 2748 8018
rect 2748 7984 2765 8018
rect 2777 7984 2782 8018
rect 2782 7984 2820 8018
rect 2820 7984 2829 8018
rect 2841 7984 2854 8018
rect 2854 7984 2892 8018
rect 2892 7984 2893 8018
rect 2905 7984 2926 8018
rect 2926 7984 2957 8018
rect 2969 7984 2998 8018
rect 2998 7984 3021 8018
rect 2585 7975 2637 7984
rect 2649 7975 2701 7984
rect 2713 7975 2765 7984
rect 2777 7975 2829 7984
rect 2841 7975 2893 7984
rect 2905 7975 2957 7984
rect 2969 7975 3021 7984
rect 3033 8018 3085 8027
rect 3033 7984 3036 8018
rect 3036 7984 3070 8018
rect 3070 7984 3085 8018
rect 3033 7975 3085 7984
rect 3097 8018 3149 8027
rect 3097 7984 3108 8018
rect 3108 7984 3142 8018
rect 3142 7984 3149 8018
rect 3097 7975 3149 7984
rect 3161 8018 3213 8027
rect 3225 8018 3277 8027
rect 3289 8018 3341 8027
rect 3353 8018 3405 8027
rect 3417 8018 3469 8027
rect 3481 8018 3533 8027
rect 3545 8018 3597 8027
rect 3161 7984 3180 8018
rect 3180 7984 3213 8018
rect 3225 7984 3252 8018
rect 3252 7984 3277 8018
rect 3289 7984 3324 8018
rect 3324 7984 3341 8018
rect 3353 7984 3358 8018
rect 3358 7984 3396 8018
rect 3396 7984 3405 8018
rect 3417 7984 3430 8018
rect 3430 7984 3468 8018
rect 3468 7984 3469 8018
rect 3481 7984 3502 8018
rect 3502 7984 3533 8018
rect 3545 7984 3574 8018
rect 3574 7984 3597 8018
rect 3161 7975 3213 7984
rect 3225 7975 3277 7984
rect 3289 7975 3341 7984
rect 3353 7975 3405 7984
rect 3417 7975 3469 7984
rect 3481 7975 3533 7984
rect 3545 7975 3597 7984
rect 3609 8018 3661 8027
rect 3609 7984 3612 8018
rect 3612 7984 3646 8018
rect 3646 7984 3661 8018
rect 3609 7975 3661 7984
rect 3673 8018 3725 8027
rect 3673 7984 3684 8018
rect 3684 7984 3718 8018
rect 3718 7984 3725 8018
rect 3673 7975 3725 7984
rect 3737 8018 3789 8027
rect 3801 8018 3853 8027
rect 3865 8018 3917 8027
rect 3929 8018 3981 8027
rect 3993 8018 4045 8027
rect 4057 8018 4109 8027
rect 4121 8018 4173 8027
rect 3737 7984 3756 8018
rect 3756 7984 3789 8018
rect 3801 7984 3828 8018
rect 3828 7984 3853 8018
rect 3865 7984 3900 8018
rect 3900 7984 3917 8018
rect 3929 7984 3934 8018
rect 3934 7984 3972 8018
rect 3972 7984 3981 8018
rect 3993 7984 4006 8018
rect 4006 7984 4044 8018
rect 4044 7984 4045 8018
rect 4057 7984 4078 8018
rect 4078 7984 4109 8018
rect 4121 7984 4150 8018
rect 4150 7984 4173 8018
rect 3737 7975 3789 7984
rect 3801 7975 3853 7984
rect 3865 7975 3917 7984
rect 3929 7975 3981 7984
rect 3993 7975 4045 7984
rect 4057 7975 4109 7984
rect 4121 7975 4173 7984
rect 4185 8018 4237 8027
rect 4185 7984 4188 8018
rect 4188 7984 4222 8018
rect 4222 7984 4237 8018
rect 4185 7975 4237 7984
rect 4249 8018 4301 8027
rect 4249 7984 4260 8018
rect 4260 7984 4294 8018
rect 4294 7984 4301 8018
rect 4249 7975 4301 7984
rect 4313 8018 4365 8027
rect 4377 8018 4429 8027
rect 4441 8018 4493 8027
rect 4505 8018 4557 8027
rect 4722 8018 4774 8027
rect 4786 8018 4838 8027
rect 4850 8018 4902 8027
rect 4914 8018 4966 8027
rect 4313 7984 4332 8018
rect 4332 7984 4365 8018
rect 4377 7984 4404 8018
rect 4404 7984 4429 8018
rect 4441 7984 4476 8018
rect 4476 7984 4493 8018
rect 4505 7984 4510 8018
rect 4510 7984 4557 8018
rect 4722 7984 4766 8018
rect 4766 7984 4774 8018
rect 4786 7984 4800 8018
rect 4800 7984 4838 8018
rect 4850 7984 4872 8018
rect 4872 7984 4902 8018
rect 4914 7984 4944 8018
rect 4944 7984 4966 8018
rect 4313 7975 4365 7984
rect 4377 7975 4429 7984
rect 4441 7975 4493 7984
rect 4505 7975 4557 7984
rect 4722 7975 4774 7984
rect 4786 7975 4838 7984
rect 4850 7975 4902 7984
rect 4914 7975 4966 7984
rect 4978 8018 5030 8027
rect 4978 7984 4982 8018
rect 4982 7984 5016 8018
rect 5016 7984 5030 8018
rect 4978 7975 5030 7984
rect 5042 8018 5094 8027
rect 5042 7984 5054 8018
rect 5054 7984 5088 8018
rect 5088 7984 5094 8018
rect 5042 7975 5094 7984
rect 5106 8018 5158 8027
rect 5170 8018 5222 8027
rect 5234 8018 5286 8027
rect 5298 8018 5350 8027
rect 5362 8018 5414 8027
rect 5426 8018 5478 8027
rect 5490 8018 5542 8027
rect 5106 7984 5126 8018
rect 5126 7984 5158 8018
rect 5170 7984 5198 8018
rect 5198 7984 5222 8018
rect 5234 7984 5270 8018
rect 5270 7984 5286 8018
rect 5298 7984 5304 8018
rect 5304 7984 5342 8018
rect 5342 7984 5350 8018
rect 5362 7984 5376 8018
rect 5376 7984 5414 8018
rect 5426 7984 5448 8018
rect 5448 7984 5478 8018
rect 5490 7984 5520 8018
rect 5520 7984 5542 8018
rect 5106 7975 5158 7984
rect 5170 7975 5222 7984
rect 5234 7975 5286 7984
rect 5298 7975 5350 7984
rect 5362 7975 5414 7984
rect 5426 7975 5478 7984
rect 5490 7975 5542 7984
rect 5554 8018 5606 8027
rect 5554 7984 5558 8018
rect 5558 7984 5592 8018
rect 5592 7984 5606 8018
rect 5554 7975 5606 7984
rect 5618 8018 5670 8027
rect 5618 7984 5630 8018
rect 5630 7984 5664 8018
rect 5664 7984 5670 8018
rect 5618 7975 5670 7984
rect 5682 8018 5734 8027
rect 5746 8018 5798 8027
rect 5810 8018 5862 8027
rect 5874 8018 5926 8027
rect 5938 8018 5990 8027
rect 6002 8018 6054 8027
rect 6066 8018 6118 8027
rect 5682 7984 5702 8018
rect 5702 7984 5734 8018
rect 5746 7984 5774 8018
rect 5774 7984 5798 8018
rect 5810 7984 5846 8018
rect 5846 7984 5862 8018
rect 5874 7984 5880 8018
rect 5880 7984 5918 8018
rect 5918 7984 5926 8018
rect 5938 7984 5952 8018
rect 5952 7984 5990 8018
rect 6002 7984 6024 8018
rect 6024 7984 6054 8018
rect 6066 7984 6096 8018
rect 6096 7984 6118 8018
rect 5682 7975 5734 7984
rect 5746 7975 5798 7984
rect 5810 7975 5862 7984
rect 5874 7975 5926 7984
rect 5938 7975 5990 7984
rect 6002 7975 6054 7984
rect 6066 7975 6118 7984
rect 6130 8018 6182 8027
rect 6130 7984 6134 8018
rect 6134 7984 6168 8018
rect 6168 7984 6182 8018
rect 6130 7975 6182 7984
rect 6194 8018 6246 8027
rect 6194 7984 6206 8018
rect 6206 7984 6240 8018
rect 6240 7984 6246 8018
rect 6194 7975 6246 7984
rect 6258 8018 6310 8027
rect 6322 8018 6374 8027
rect 6386 8018 6438 8027
rect 6450 8018 6502 8027
rect 6514 8018 6566 8027
rect 6578 8018 6630 8027
rect 6810 8018 6862 8027
rect 6874 8018 6926 8027
rect 6938 8018 6990 8027
rect 7002 8018 7054 8027
rect 6258 7984 6278 8018
rect 6278 7984 6310 8018
rect 6322 7984 6350 8018
rect 6350 7984 6374 8018
rect 6386 7984 6422 8018
rect 6422 7984 6438 8018
rect 6450 7984 6456 8018
rect 6456 7984 6494 8018
rect 6494 7984 6502 8018
rect 6514 7984 6528 8018
rect 6528 7984 6566 8018
rect 6578 7984 6600 8018
rect 6600 7984 6630 8018
rect 6810 7984 6850 8018
rect 6850 7984 6862 8018
rect 6874 7984 6884 8018
rect 6884 7984 6922 8018
rect 6922 7984 6926 8018
rect 6938 7984 6956 8018
rect 6956 7984 6990 8018
rect 7002 7984 7028 8018
rect 7028 7984 7054 8018
rect 6258 7975 6310 7984
rect 6322 7975 6374 7984
rect 6386 7975 6438 7984
rect 6450 7975 6502 7984
rect 6514 7975 6566 7984
rect 6578 7975 6630 7984
rect 6810 7975 6862 7984
rect 6874 7975 6926 7984
rect 6938 7975 6990 7984
rect 7002 7975 7054 7984
rect 7066 8018 7118 8027
rect 7066 7984 7100 8018
rect 7100 7984 7118 8018
rect 7066 7975 7118 7984
rect 7130 8018 7182 8027
rect 7130 7984 7138 8018
rect 7138 7984 7172 8018
rect 7172 7984 7182 8018
rect 7130 7975 7182 7984
rect 7194 8018 7246 8027
rect 7194 7984 7210 8018
rect 7210 7984 7244 8018
rect 7244 7984 7246 8018
rect 7194 7975 7246 7984
rect 7258 8018 7310 8027
rect 7322 8018 7374 8027
rect 7386 8018 7438 8027
rect 7450 8018 7502 8027
rect 7514 8018 7566 8027
rect 7578 8018 7630 8027
rect 7258 7984 7282 8018
rect 7282 7984 7310 8018
rect 7322 7984 7354 8018
rect 7354 7984 7374 8018
rect 7386 7984 7388 8018
rect 7388 7984 7426 8018
rect 7426 7984 7438 8018
rect 7450 7984 7460 8018
rect 7460 7984 7498 8018
rect 7498 7984 7502 8018
rect 7514 7984 7532 8018
rect 7532 7984 7566 8018
rect 7578 7984 7604 8018
rect 7604 7984 7630 8018
rect 7258 7975 7310 7984
rect 7322 7975 7374 7984
rect 7386 7975 7438 7984
rect 7450 7975 7502 7984
rect 7514 7975 7566 7984
rect 7578 7975 7630 7984
rect 7642 8018 7694 8027
rect 7642 7984 7676 8018
rect 7676 7984 7694 8018
rect 7642 7975 7694 7984
rect 7706 8018 7758 8027
rect 7706 7984 7714 8018
rect 7714 7984 7748 8018
rect 7748 7984 7758 8018
rect 7706 7975 7758 7984
rect 7770 8018 7822 8027
rect 7770 7984 7786 8018
rect 7786 7984 7820 8018
rect 7820 7984 7822 8018
rect 7770 7975 7822 7984
rect 7834 8018 7886 8027
rect 7898 8018 7950 8027
rect 7962 8018 8014 8027
rect 8026 8018 8078 8027
rect 8090 8018 8142 8027
rect 8154 8018 8206 8027
rect 7834 7984 7858 8018
rect 7858 7984 7886 8018
rect 7898 7984 7930 8018
rect 7930 7984 7950 8018
rect 7962 7984 7964 8018
rect 7964 7984 8002 8018
rect 8002 7984 8014 8018
rect 8026 7984 8036 8018
rect 8036 7984 8074 8018
rect 8074 7984 8078 8018
rect 8090 7984 8108 8018
rect 8108 7984 8142 8018
rect 8154 7984 8180 8018
rect 8180 7984 8206 8018
rect 7834 7975 7886 7984
rect 7898 7975 7950 7984
rect 7962 7975 8014 7984
rect 8026 7975 8078 7984
rect 8090 7975 8142 7984
rect 8154 7975 8206 7984
rect 8218 8018 8270 8027
rect 8218 7984 8252 8018
rect 8252 7984 8270 8018
rect 8218 7975 8270 7984
rect 8282 8018 8334 8027
rect 8282 7984 8290 8018
rect 8290 7984 8324 8018
rect 8324 7984 8334 8018
rect 8282 7975 8334 7984
rect 8346 8018 8398 8027
rect 8346 7984 8362 8018
rect 8362 7984 8396 8018
rect 8396 7984 8398 8018
rect 8346 7975 8398 7984
rect 8410 8018 8462 8027
rect 8474 8018 8526 8027
rect 8538 8018 8590 8027
rect 8602 8018 8654 8027
rect 8666 8018 8718 8027
rect 8730 8018 8782 8027
rect 8410 7984 8434 8018
rect 8434 7984 8462 8018
rect 8474 7984 8506 8018
rect 8506 7984 8526 8018
rect 8538 7984 8540 8018
rect 8540 7984 8578 8018
rect 8578 7984 8590 8018
rect 8602 7984 8612 8018
rect 8612 7984 8650 8018
rect 8650 7984 8654 8018
rect 8666 7984 8684 8018
rect 8684 7984 8718 8018
rect 8730 7984 8756 8018
rect 8756 7984 8782 8018
rect 8410 7975 8462 7984
rect 8474 7975 8526 7984
rect 8538 7975 8590 7984
rect 8602 7975 8654 7984
rect 8666 7975 8718 7984
rect 8730 7975 8782 7984
rect 8794 8018 8846 8027
rect 8794 7984 8828 8018
rect 8828 7984 8846 8018
rect 8794 7975 8846 7984
rect 8858 8018 8910 8027
rect 8858 7984 8866 8018
rect 8866 7984 8900 8018
rect 8900 7984 8910 8018
rect 8858 7975 8910 7984
rect 8922 8018 8974 8027
rect 8922 7984 8938 8018
rect 8938 7984 8972 8018
rect 8972 7984 8974 8018
rect 8922 7975 8974 7984
rect 8986 8018 9038 8027
rect 9050 8018 9102 8027
rect 9114 8018 9166 8027
rect 9178 8018 9230 8027
rect 9242 8018 9294 8027
rect 9306 8018 9358 8027
rect 8986 7984 9010 8018
rect 9010 7984 9038 8018
rect 9050 7984 9082 8018
rect 9082 7984 9102 8018
rect 9114 7984 9116 8018
rect 9116 7984 9154 8018
rect 9154 7984 9166 8018
rect 9178 7984 9188 8018
rect 9188 7984 9226 8018
rect 9226 7984 9230 8018
rect 9242 7984 9260 8018
rect 9260 7984 9294 8018
rect 9306 7984 9332 8018
rect 9332 7984 9358 8018
rect 8986 7975 9038 7984
rect 9050 7975 9102 7984
rect 9114 7975 9166 7984
rect 9178 7975 9230 7984
rect 9242 7975 9294 7984
rect 9306 7975 9358 7984
rect 9370 8018 9422 8027
rect 9370 7984 9404 8018
rect 9404 7984 9422 8018
rect 9370 7975 9422 7984
rect 9434 8018 9486 8027
rect 9434 7984 9442 8018
rect 9442 7984 9476 8018
rect 9476 7984 9486 8018
rect 9434 7975 9486 7984
rect 9498 8018 9550 8027
rect 9498 7984 9514 8018
rect 9514 7984 9548 8018
rect 9548 7984 9550 8018
rect 9498 7975 9550 7984
rect 9562 8018 9614 8027
rect 9626 8018 9678 8027
rect 9690 8018 9742 8027
rect 9754 8018 9806 8027
rect 9818 8018 9870 8027
rect 9882 8018 9934 8027
rect 9562 7984 9586 8018
rect 9586 7984 9614 8018
rect 9626 7984 9658 8018
rect 9658 7984 9678 8018
rect 9690 7984 9692 8018
rect 9692 7984 9730 8018
rect 9730 7984 9742 8018
rect 9754 7984 9764 8018
rect 9764 7984 9802 8018
rect 9802 7984 9806 8018
rect 9818 7984 9836 8018
rect 9836 7984 9870 8018
rect 9882 7984 9908 8018
rect 9908 7984 9934 8018
rect 9562 7975 9614 7984
rect 9626 7975 9678 7984
rect 9690 7975 9742 7984
rect 9754 7975 9806 7984
rect 9818 7975 9870 7984
rect 9882 7975 9934 7984
rect 9946 8018 9998 8027
rect 9946 7984 9980 8018
rect 9980 7984 9998 8018
rect 9946 7975 9998 7984
rect 10010 8018 10062 8027
rect 10010 7984 10018 8018
rect 10018 7984 10052 8018
rect 10052 7984 10062 8018
rect 10010 7975 10062 7984
rect 10074 8018 10126 8027
rect 10074 7984 10090 8018
rect 10090 7984 10124 8018
rect 10124 7984 10126 8018
rect 10074 7975 10126 7984
rect 10138 8018 10190 8027
rect 10202 8018 10254 8027
rect 10266 8018 10318 8027
rect 10330 8018 10382 8027
rect 10394 8018 10446 8027
rect 10458 8018 10510 8027
rect 10138 7984 10162 8018
rect 10162 7984 10190 8018
rect 10202 7984 10234 8018
rect 10234 7984 10254 8018
rect 10266 7984 10268 8018
rect 10268 7984 10306 8018
rect 10306 7984 10318 8018
rect 10330 7984 10340 8018
rect 10340 7984 10378 8018
rect 10378 7984 10382 8018
rect 10394 7984 10412 8018
rect 10412 7984 10446 8018
rect 10458 7984 10484 8018
rect 10484 7984 10510 8018
rect 10138 7975 10190 7984
rect 10202 7975 10254 7984
rect 10266 7975 10318 7984
rect 10330 7975 10382 7984
rect 10394 7975 10446 7984
rect 10458 7975 10510 7984
rect 10522 8018 10574 8027
rect 10522 7984 10556 8018
rect 10556 7984 10574 8018
rect 10522 7975 10574 7984
rect 10586 8018 10638 8027
rect 10586 7984 10594 8018
rect 10594 7984 10628 8018
rect 10628 7984 10638 8018
rect 10586 7975 10638 7984
rect 10650 8018 10702 8027
rect 10650 7984 10666 8018
rect 10666 7984 10700 8018
rect 10700 7984 10702 8018
rect 10650 7975 10702 7984
rect 10714 8018 10766 8027
rect 10778 8018 10830 8027
rect 10842 8018 10894 8027
rect 10906 8018 10958 8027
rect 10970 8018 11022 8027
rect 11034 8018 11086 8027
rect 10714 7984 10738 8018
rect 10738 7984 10766 8018
rect 10778 7984 10810 8018
rect 10810 7984 10830 8018
rect 10842 7984 10844 8018
rect 10844 7984 10882 8018
rect 10882 7984 10894 8018
rect 10906 7984 10916 8018
rect 10916 7984 10954 8018
rect 10954 7984 10958 8018
rect 10970 7984 10988 8018
rect 10988 7984 11022 8018
rect 11034 7984 11060 8018
rect 11060 7984 11086 8018
rect 10714 7975 10766 7984
rect 10778 7975 10830 7984
rect 10842 7975 10894 7984
rect 10906 7975 10958 7984
rect 10970 7975 11022 7984
rect 11034 7975 11086 7984
rect 11098 8018 11150 8027
rect 11098 7984 11132 8018
rect 11132 7984 11150 8018
rect 11098 7975 11150 7984
rect 11162 8018 11214 8027
rect 11162 7984 11170 8018
rect 11170 7984 11204 8018
rect 11204 7984 11214 8018
rect 11162 7975 11214 7984
rect 11226 8018 11278 8027
rect 11226 7984 11242 8018
rect 11242 7984 11276 8018
rect 11276 7984 11278 8018
rect 11226 7975 11278 7984
rect 11290 8018 11342 8027
rect 11354 8018 11406 8027
rect 11418 8018 11470 8027
rect 11482 8018 11534 8027
rect 11546 8018 11598 8027
rect 11610 8018 11662 8027
rect 11290 7984 11314 8018
rect 11314 7984 11342 8018
rect 11354 7984 11386 8018
rect 11386 7984 11406 8018
rect 11418 7984 11420 8018
rect 11420 7984 11458 8018
rect 11458 7984 11470 8018
rect 11482 7984 11492 8018
rect 11492 7984 11530 8018
rect 11530 7984 11534 8018
rect 11546 7984 11564 8018
rect 11564 7984 11598 8018
rect 11610 7984 11636 8018
rect 11636 7984 11662 8018
rect 11290 7975 11342 7984
rect 11354 7975 11406 7984
rect 11418 7975 11470 7984
rect 11482 7975 11534 7984
rect 11546 7975 11598 7984
rect 11610 7975 11662 7984
rect 11674 8018 11726 8027
rect 11674 7984 11708 8018
rect 11708 7984 11726 8018
rect 11674 7975 11726 7984
rect 11738 8018 11790 8027
rect 11738 7984 11746 8018
rect 11746 7984 11780 8018
rect 11780 7984 11790 8018
rect 11738 7975 11790 7984
rect 11802 8018 11854 8027
rect 11802 7984 11818 8018
rect 11818 7984 11852 8018
rect 11852 7984 11854 8018
rect 11802 7975 11854 7984
rect 11866 8018 11918 8027
rect 11930 8018 11982 8027
rect 11994 8018 12046 8027
rect 12058 8018 12110 8027
rect 12122 8018 12174 8027
rect 12186 8018 12238 8027
rect 11866 7984 11890 8018
rect 11890 7984 11918 8018
rect 11930 7984 11962 8018
rect 11962 7984 11982 8018
rect 11994 7984 11996 8018
rect 11996 7984 12034 8018
rect 12034 7984 12046 8018
rect 12058 7984 12068 8018
rect 12068 7984 12106 8018
rect 12106 7984 12110 8018
rect 12122 7984 12140 8018
rect 12140 7984 12174 8018
rect 12186 7984 12212 8018
rect 12212 7984 12238 8018
rect 11866 7975 11918 7984
rect 11930 7975 11982 7984
rect 11994 7975 12046 7984
rect 12058 7975 12110 7984
rect 12122 7975 12174 7984
rect 12186 7975 12238 7984
rect 12250 8018 12302 8027
rect 12250 7984 12284 8018
rect 12284 7984 12302 8018
rect 12250 7975 12302 7984
rect 12314 8018 12366 8027
rect 12314 7984 12322 8018
rect 12322 7984 12356 8018
rect 12356 7984 12366 8018
rect 12314 7975 12366 7984
rect 12378 8018 12430 8027
rect 12378 7984 12394 8018
rect 12394 7984 12428 8018
rect 12428 7984 12430 8018
rect 12378 7975 12430 7984
rect 12442 8018 12494 8027
rect 12506 8018 12558 8027
rect 12570 8018 12622 8027
rect 12634 8018 12686 8027
rect 12698 8018 12750 8027
rect 12762 8018 12814 8027
rect 12442 7984 12466 8018
rect 12466 7984 12494 8018
rect 12506 7984 12538 8018
rect 12538 7984 12558 8018
rect 12570 7984 12572 8018
rect 12572 7984 12610 8018
rect 12610 7984 12622 8018
rect 12634 7984 12644 8018
rect 12644 7984 12682 8018
rect 12682 7984 12686 8018
rect 12698 7984 12716 8018
rect 12716 7984 12750 8018
rect 12762 7984 12788 8018
rect 12788 7984 12814 8018
rect 12442 7975 12494 7984
rect 12506 7975 12558 7984
rect 12570 7975 12622 7984
rect 12634 7975 12686 7984
rect 12698 7975 12750 7984
rect 12762 7975 12814 7984
rect 12826 8018 12878 8027
rect 12826 7984 12860 8018
rect 12860 7984 12878 8018
rect 12826 7975 12878 7984
rect 12890 8018 12942 8027
rect 12890 7984 12898 8018
rect 12898 7984 12932 8018
rect 12932 7984 12942 8018
rect 12890 7975 12942 7984
rect 12954 8018 13006 8027
rect 12954 7984 12970 8018
rect 12970 7984 13004 8018
rect 13004 7984 13006 8018
rect 12954 7975 13006 7984
rect 13018 8018 13070 8027
rect 13082 8018 13134 8027
rect 13146 8018 13198 8027
rect 13210 8018 13262 8027
rect 13274 8018 13326 8027
rect 13338 8018 13390 8027
rect 13018 7984 13042 8018
rect 13042 7984 13070 8018
rect 13082 7984 13114 8018
rect 13114 7984 13134 8018
rect 13146 7984 13148 8018
rect 13148 7984 13186 8018
rect 13186 7984 13198 8018
rect 13210 7984 13220 8018
rect 13220 7984 13258 8018
rect 13258 7984 13262 8018
rect 13274 7984 13292 8018
rect 13292 7984 13326 8018
rect 13338 7984 13364 8018
rect 13364 7984 13390 8018
rect 13018 7975 13070 7984
rect 13082 7975 13134 7984
rect 13146 7975 13198 7984
rect 13210 7975 13262 7984
rect 13274 7975 13326 7984
rect 13338 7975 13390 7984
rect 13402 8018 13454 8027
rect 13402 7984 13436 8018
rect 13436 7984 13454 8018
rect 13402 7975 13454 7984
rect 13466 8018 13518 8027
rect 13466 7984 13474 8018
rect 13474 7984 13508 8018
rect 13508 7984 13518 8018
rect 13466 7975 13518 7984
rect 13530 8018 13582 8027
rect 13530 7984 13546 8018
rect 13546 7984 13580 8018
rect 13580 7984 13582 8018
rect 13530 7975 13582 7984
rect 13594 7975 13646 8027
rect 473 7873 525 7882
rect 473 7839 478 7873
rect 478 7839 512 7873
rect 512 7839 525 7873
rect 473 7830 525 7839
rect 537 7873 589 7882
rect 537 7839 550 7873
rect 550 7839 584 7873
rect 584 7839 589 7873
rect 537 7830 589 7839
rect 3209 7830 3261 7882
rect 3273 7830 3325 7882
rect 473 7719 525 7728
rect 473 7685 478 7719
rect 478 7685 512 7719
rect 512 7685 525 7719
rect 473 7676 525 7685
rect 537 7719 589 7728
rect 537 7685 550 7719
rect 550 7685 584 7719
rect 584 7685 589 7719
rect 537 7676 589 7685
rect 3213 7676 3265 7728
rect 3277 7676 3329 7728
rect 10285 7676 10337 7728
rect 10349 7676 10401 7728
rect 473 7565 525 7574
rect 473 7531 478 7565
rect 478 7531 512 7565
rect 512 7531 525 7565
rect 473 7522 525 7531
rect 537 7565 589 7574
rect 537 7531 550 7565
rect 550 7531 584 7565
rect 584 7531 589 7565
rect 537 7522 589 7531
rect 3209 7522 3261 7574
rect 3273 7522 3325 7574
rect 473 7411 525 7420
rect 473 7377 478 7411
rect 478 7377 512 7411
rect 512 7377 525 7411
rect 473 7368 525 7377
rect 537 7411 589 7420
rect 537 7377 550 7411
rect 550 7377 584 7411
rect 584 7377 589 7411
rect 537 7368 589 7377
rect 3213 7368 3265 7420
rect 3277 7368 3329 7420
rect 9429 7368 9481 7420
rect 9493 7368 9545 7420
rect 473 7257 525 7266
rect 473 7223 478 7257
rect 478 7223 512 7257
rect 512 7223 525 7257
rect 473 7214 525 7223
rect 537 7257 589 7266
rect 537 7223 550 7257
rect 550 7223 584 7257
rect 584 7223 589 7257
rect 537 7214 589 7223
rect 3209 7214 3261 7266
rect 3273 7214 3325 7266
rect 473 7103 525 7112
rect 473 7069 478 7103
rect 478 7069 512 7103
rect 512 7069 525 7103
rect 473 7060 525 7069
rect 537 7103 589 7112
rect 537 7069 550 7103
rect 550 7069 584 7103
rect 584 7069 589 7103
rect 537 7060 589 7069
rect 3213 7060 3265 7112
rect 3277 7060 3329 7112
rect 8573 7060 8625 7112
rect 8637 7060 8689 7112
rect 473 6949 525 6958
rect 473 6915 478 6949
rect 478 6915 512 6949
rect 512 6915 525 6949
rect 473 6906 525 6915
rect 537 6949 589 6958
rect 537 6915 550 6949
rect 550 6915 584 6949
rect 584 6915 589 6949
rect 537 6906 589 6915
rect 3209 6906 3261 6958
rect 3273 6906 3325 6958
rect 473 6795 525 6804
rect 473 6761 478 6795
rect 478 6761 512 6795
rect 512 6761 525 6795
rect 473 6752 525 6761
rect 537 6795 589 6804
rect 537 6761 550 6795
rect 550 6761 584 6795
rect 584 6761 589 6795
rect 537 6752 589 6761
rect 3213 6752 3265 6804
rect 3277 6752 3329 6804
rect 7717 6752 7769 6804
rect 7781 6752 7833 6804
rect 473 6641 525 6650
rect 473 6607 478 6641
rect 478 6607 512 6641
rect 512 6607 525 6641
rect 473 6598 525 6607
rect 537 6641 589 6650
rect 537 6607 550 6641
rect 550 6607 584 6641
rect 584 6607 589 6641
rect 537 6598 589 6607
rect 3209 6598 3261 6650
rect 3273 6598 3325 6650
rect 473 6487 525 6496
rect 473 6453 478 6487
rect 478 6453 512 6487
rect 512 6453 525 6487
rect 473 6444 525 6453
rect 537 6487 589 6496
rect 537 6453 550 6487
rect 550 6453 584 6487
rect 584 6453 589 6487
rect 537 6444 589 6453
rect 3213 6444 3265 6496
rect 3277 6444 3329 6496
rect 6861 6444 6913 6496
rect 6925 6444 6977 6496
rect 473 6333 525 6342
rect 473 6299 478 6333
rect 478 6299 512 6333
rect 512 6299 525 6333
rect 473 6290 525 6299
rect 537 6333 589 6342
rect 537 6299 550 6333
rect 550 6299 584 6333
rect 584 6299 589 6333
rect 537 6290 589 6299
rect 3209 6290 3261 6342
rect 3273 6290 3325 6342
rect 473 6179 525 6188
rect 473 6145 478 6179
rect 478 6145 512 6179
rect 512 6145 525 6179
rect 473 6136 525 6145
rect 537 6179 589 6188
rect 537 6145 550 6179
rect 550 6145 584 6179
rect 584 6145 589 6179
rect 537 6136 589 6145
rect 3213 6136 3265 6188
rect 3277 6136 3329 6188
rect 6005 6136 6057 6188
rect 6069 6136 6121 6188
rect 354 6033 406 6042
rect 418 6033 470 6042
rect 482 6033 534 6042
rect 546 6033 598 6042
rect 610 6033 662 6042
rect 354 5999 389 6033
rect 389 5999 406 6033
rect 418 5999 423 6033
rect 423 5999 461 6033
rect 461 5999 470 6033
rect 482 5999 495 6033
rect 495 5999 533 6033
rect 533 5999 534 6033
rect 546 5999 567 6033
rect 567 5999 598 6033
rect 610 5999 639 6033
rect 639 5999 662 6033
rect 354 5990 406 5999
rect 418 5990 470 5999
rect 482 5990 534 5999
rect 546 5990 598 5999
rect 610 5990 662 5999
rect 674 6033 726 6042
rect 674 5999 677 6033
rect 677 5999 711 6033
rect 711 5999 726 6033
rect 869 6033 921 6042
rect 933 6033 985 6042
rect 997 6033 1049 6042
rect 1061 6033 1113 6042
rect 869 6032 914 6033
rect 674 5990 726 5999
rect 869 5998 871 6032
rect 871 5999 914 6032
rect 914 5999 921 6033
rect 933 5999 948 6033
rect 948 5999 985 6033
rect 997 5999 1020 6033
rect 1020 5999 1049 6033
rect 1061 5999 1092 6033
rect 1092 5999 1113 6033
rect 871 5998 921 5999
rect 869 5990 921 5998
rect 933 5990 985 5999
rect 997 5990 1049 5999
rect 1061 5990 1113 5999
rect 1125 6033 1177 6042
rect 1125 5999 1130 6033
rect 1130 5999 1164 6033
rect 1164 5999 1177 6033
rect 1125 5990 1177 5999
rect 1189 6033 1241 6042
rect 1189 5999 1202 6033
rect 1202 5999 1236 6033
rect 1236 5999 1241 6033
rect 1189 5990 1241 5999
rect 1253 6033 1305 6042
rect 1317 6033 1369 6042
rect 1381 6033 1433 6042
rect 1445 6033 1497 6042
rect 1509 6033 1561 6042
rect 1573 6033 1625 6042
rect 1637 6033 1689 6042
rect 1253 5999 1274 6033
rect 1274 5999 1305 6033
rect 1317 5999 1346 6033
rect 1346 5999 1369 6033
rect 1381 5999 1418 6033
rect 1418 5999 1433 6033
rect 1445 5999 1452 6033
rect 1452 5999 1490 6033
rect 1490 5999 1497 6033
rect 1509 5999 1524 6033
rect 1524 5999 1561 6033
rect 1573 5999 1596 6033
rect 1596 5999 1625 6033
rect 1637 5999 1668 6033
rect 1668 5999 1689 6033
rect 1253 5990 1305 5999
rect 1317 5990 1369 5999
rect 1381 5990 1433 5999
rect 1445 5990 1497 5999
rect 1509 5990 1561 5999
rect 1573 5990 1625 5999
rect 1637 5990 1689 5999
rect 1701 6033 1753 6042
rect 1701 5999 1706 6033
rect 1706 5999 1740 6033
rect 1740 5999 1753 6033
rect 1701 5990 1753 5999
rect 1765 6033 1817 6042
rect 1765 5999 1778 6033
rect 1778 5999 1812 6033
rect 1812 5999 1817 6033
rect 1765 5990 1817 5999
rect 1829 6033 1881 6042
rect 1893 6033 1945 6042
rect 1957 6033 2009 6042
rect 2021 6033 2073 6042
rect 2085 6033 2137 6042
rect 2149 6033 2201 6042
rect 2213 6033 2265 6042
rect 1829 5999 1850 6033
rect 1850 5999 1881 6033
rect 1893 5999 1922 6033
rect 1922 5999 1945 6033
rect 1957 5999 1994 6033
rect 1994 5999 2009 6033
rect 2021 5999 2028 6033
rect 2028 5999 2066 6033
rect 2066 5999 2073 6033
rect 2085 5999 2100 6033
rect 2100 5999 2137 6033
rect 2149 5999 2172 6033
rect 2172 5999 2201 6033
rect 2213 5999 2244 6033
rect 2244 5999 2265 6033
rect 1829 5990 1881 5999
rect 1893 5990 1945 5999
rect 1957 5990 2009 5999
rect 2021 5990 2073 5999
rect 2085 5990 2137 5999
rect 2149 5990 2201 5999
rect 2213 5990 2265 5999
rect 2277 6033 2329 6042
rect 2277 5999 2282 6033
rect 2282 5999 2316 6033
rect 2316 5999 2329 6033
rect 2277 5990 2329 5999
rect 2341 6033 2393 6042
rect 2341 5999 2354 6033
rect 2354 5999 2388 6033
rect 2388 5999 2393 6033
rect 2341 5990 2393 5999
rect 2405 6033 2457 6042
rect 2469 6033 2521 6042
rect 2533 6033 2585 6042
rect 2597 6033 2649 6042
rect 2661 6033 2713 6042
rect 2725 6033 2777 6042
rect 2789 6033 2841 6042
rect 2405 5999 2426 6033
rect 2426 5999 2457 6033
rect 2469 5999 2498 6033
rect 2498 5999 2521 6033
rect 2533 5999 2570 6033
rect 2570 5999 2585 6033
rect 2597 5999 2604 6033
rect 2604 5999 2642 6033
rect 2642 5999 2649 6033
rect 2661 5999 2676 6033
rect 2676 5999 2713 6033
rect 2725 5999 2748 6033
rect 2748 5999 2777 6033
rect 2789 5999 2820 6033
rect 2820 5999 2841 6033
rect 2405 5990 2457 5999
rect 2469 5990 2521 5999
rect 2533 5990 2585 5999
rect 2597 5990 2649 5999
rect 2661 5990 2713 5999
rect 2725 5990 2777 5999
rect 2789 5990 2841 5999
rect 2853 6033 2905 6042
rect 2853 5999 2858 6033
rect 2858 5999 2892 6033
rect 2892 5999 2905 6033
rect 2853 5990 2905 5999
rect 2917 6033 2969 6042
rect 2917 5999 2930 6033
rect 2930 5999 2964 6033
rect 2964 5999 2969 6033
rect 2917 5990 2969 5999
rect 2981 6033 3033 6042
rect 3045 6033 3097 6042
rect 3109 6033 3161 6042
rect 3173 6033 3225 6042
rect 3237 6033 3289 6042
rect 3301 6033 3353 6042
rect 3365 6033 3417 6042
rect 2981 5999 3002 6033
rect 3002 5999 3033 6033
rect 3045 5999 3074 6033
rect 3074 5999 3097 6033
rect 3109 5999 3146 6033
rect 3146 5999 3161 6033
rect 3173 5999 3180 6033
rect 3180 5999 3218 6033
rect 3218 5999 3225 6033
rect 3237 5999 3252 6033
rect 3252 5999 3289 6033
rect 3301 5999 3324 6033
rect 3324 5999 3353 6033
rect 3365 5999 3396 6033
rect 3396 5999 3417 6033
rect 2981 5990 3033 5999
rect 3045 5990 3097 5999
rect 3109 5990 3161 5999
rect 3173 5990 3225 5999
rect 3237 5990 3289 5999
rect 3301 5990 3353 5999
rect 3365 5990 3417 5999
rect 3429 6033 3481 6042
rect 3429 5999 3434 6033
rect 3434 5999 3468 6033
rect 3468 5999 3481 6033
rect 3429 5990 3481 5999
rect 3493 6033 3545 6042
rect 3493 5999 3506 6033
rect 3506 5999 3540 6033
rect 3540 5999 3545 6033
rect 3493 5990 3545 5999
rect 3557 6033 3609 6042
rect 3621 6033 3673 6042
rect 3685 6033 3737 6042
rect 3749 6033 3801 6042
rect 3813 6033 3865 6042
rect 3877 6033 3929 6042
rect 3941 6033 3993 6042
rect 3557 5999 3578 6033
rect 3578 5999 3609 6033
rect 3621 5999 3650 6033
rect 3650 5999 3673 6033
rect 3685 5999 3722 6033
rect 3722 5999 3737 6033
rect 3749 5999 3756 6033
rect 3756 5999 3794 6033
rect 3794 5999 3801 6033
rect 3813 5999 3828 6033
rect 3828 5999 3865 6033
rect 3877 5999 3900 6033
rect 3900 5999 3929 6033
rect 3941 5999 3972 6033
rect 3972 5999 3993 6033
rect 3557 5990 3609 5999
rect 3621 5990 3673 5999
rect 3685 5990 3737 5999
rect 3749 5990 3801 5999
rect 3813 5990 3865 5999
rect 3877 5990 3929 5999
rect 3941 5990 3993 5999
rect 4005 6033 4057 6042
rect 4005 5999 4010 6033
rect 4010 5999 4044 6033
rect 4044 5999 4057 6033
rect 4005 5990 4057 5999
rect 4069 6033 4121 6042
rect 4069 5999 4082 6033
rect 4082 5999 4116 6033
rect 4116 5999 4121 6033
rect 4069 5990 4121 5999
rect 4133 6033 4185 6042
rect 4197 6033 4249 6042
rect 4261 6033 4313 6042
rect 4325 6033 4377 6042
rect 4389 6033 4441 6042
rect 4453 6033 4505 6042
rect 4517 6033 4569 6042
rect 4133 5999 4154 6033
rect 4154 5999 4185 6033
rect 4197 5999 4226 6033
rect 4226 5999 4249 6033
rect 4261 5999 4298 6033
rect 4298 5999 4313 6033
rect 4325 5999 4332 6033
rect 4332 5999 4370 6033
rect 4370 5999 4377 6033
rect 4389 5999 4404 6033
rect 4404 5999 4441 6033
rect 4453 5999 4476 6033
rect 4476 5999 4505 6033
rect 4517 5999 4548 6033
rect 4548 5999 4569 6033
rect 4757 6033 4809 6042
rect 4133 5990 4185 5999
rect 4197 5990 4249 5999
rect 4261 5990 4313 5999
rect 4325 5990 4377 5999
rect 4389 5990 4441 5999
rect 4453 5990 4505 5999
rect 4517 5990 4569 5999
rect 4757 5999 4773 6033
rect 4773 5999 4807 6033
rect 4807 5999 4809 6033
rect 4757 5990 4809 5999
rect 4821 6033 4873 6042
rect 4885 6033 4937 6042
rect 4949 6033 5001 6042
rect 5013 6033 5065 6042
rect 5077 6033 5129 6042
rect 5141 6033 5193 6042
rect 4821 5999 4845 6033
rect 4845 5999 4873 6033
rect 4885 5999 4917 6033
rect 4917 5999 4937 6033
rect 4949 5999 4951 6033
rect 4951 5999 4989 6033
rect 4989 5999 5001 6033
rect 5013 5999 5023 6033
rect 5023 5999 5061 6033
rect 5061 5999 5065 6033
rect 5077 5999 5095 6033
rect 5095 5999 5129 6033
rect 5141 5999 5167 6033
rect 5167 5999 5193 6033
rect 4821 5990 4873 5999
rect 4885 5990 4937 5999
rect 4949 5990 5001 5999
rect 5013 5990 5065 5999
rect 5077 5990 5129 5999
rect 5141 5990 5193 5999
rect 5205 6033 5257 6042
rect 5205 5999 5239 6033
rect 5239 5999 5257 6033
rect 5205 5990 5257 5999
rect 5269 6033 5321 6042
rect 5269 5999 5277 6033
rect 5277 5999 5311 6033
rect 5311 5999 5321 6033
rect 5269 5990 5321 5999
rect 5333 6033 5385 6042
rect 5333 5999 5349 6033
rect 5349 5999 5383 6033
rect 5383 5999 5385 6033
rect 5333 5990 5385 5999
rect 5397 6033 5449 6042
rect 5461 6033 5513 6042
rect 5525 6033 5577 6042
rect 5589 6033 5641 6042
rect 5653 6033 5705 6042
rect 5717 6033 5769 6042
rect 5397 5999 5421 6033
rect 5421 5999 5449 6033
rect 5461 5999 5493 6033
rect 5493 5999 5513 6033
rect 5525 5999 5527 6033
rect 5527 5999 5565 6033
rect 5565 5999 5577 6033
rect 5589 5999 5599 6033
rect 5599 5999 5637 6033
rect 5637 5999 5641 6033
rect 5653 5999 5671 6033
rect 5671 5999 5705 6033
rect 5717 5999 5743 6033
rect 5743 5999 5769 6033
rect 5397 5990 5449 5999
rect 5461 5990 5513 5999
rect 5525 5990 5577 5999
rect 5589 5990 5641 5999
rect 5653 5990 5705 5999
rect 5717 5990 5769 5999
rect 5781 6033 5833 6042
rect 5781 5999 5815 6033
rect 5815 5999 5833 6033
rect 5781 5990 5833 5999
rect 5845 6033 5897 6042
rect 5845 5999 5853 6033
rect 5853 5999 5887 6033
rect 5887 5999 5897 6033
rect 5845 5990 5897 5999
rect 354 5765 406 5808
rect 354 5756 360 5765
rect 360 5756 394 5765
rect 394 5756 406 5765
rect 418 5799 470 5808
rect 418 5765 434 5799
rect 434 5765 468 5799
rect 468 5765 470 5799
rect 418 5756 470 5765
rect 482 5799 534 5808
rect 546 5799 598 5808
rect 610 5799 662 5808
rect 674 5799 726 5808
rect 738 5799 790 5808
rect 802 5799 854 5808
rect 482 5765 506 5799
rect 506 5765 534 5799
rect 546 5765 578 5799
rect 578 5765 598 5799
rect 610 5765 612 5799
rect 612 5765 650 5799
rect 650 5765 662 5799
rect 674 5765 684 5799
rect 684 5765 722 5799
rect 722 5765 726 5799
rect 738 5765 756 5799
rect 756 5765 790 5799
rect 802 5765 828 5799
rect 828 5765 854 5799
rect 482 5756 534 5765
rect 546 5756 598 5765
rect 610 5756 662 5765
rect 674 5756 726 5765
rect 738 5756 790 5765
rect 802 5756 854 5765
rect 866 5799 918 5808
rect 866 5765 900 5799
rect 900 5765 918 5799
rect 866 5756 918 5765
rect 930 5799 982 5808
rect 930 5765 938 5799
rect 938 5765 972 5799
rect 972 5765 982 5799
rect 930 5756 982 5765
rect 994 5799 1046 5808
rect 994 5765 1010 5799
rect 1010 5765 1044 5799
rect 1044 5765 1046 5799
rect 994 5756 1046 5765
rect 1058 5799 1110 5808
rect 1122 5799 1174 5808
rect 1186 5799 1238 5808
rect 1250 5799 1302 5808
rect 1314 5799 1366 5808
rect 1378 5799 1430 5808
rect 1058 5765 1082 5799
rect 1082 5765 1110 5799
rect 1122 5765 1154 5799
rect 1154 5765 1174 5799
rect 1186 5765 1188 5799
rect 1188 5765 1226 5799
rect 1226 5765 1238 5799
rect 1250 5765 1260 5799
rect 1260 5765 1298 5799
rect 1298 5765 1302 5799
rect 1314 5765 1332 5799
rect 1332 5765 1366 5799
rect 1378 5765 1404 5799
rect 1404 5765 1430 5799
rect 1058 5756 1110 5765
rect 1122 5756 1174 5765
rect 1186 5756 1238 5765
rect 1250 5756 1302 5765
rect 1314 5756 1366 5765
rect 1378 5756 1430 5765
rect 1442 5799 1494 5808
rect 1442 5765 1476 5799
rect 1476 5765 1494 5799
rect 1442 5756 1494 5765
rect 1506 5799 1558 5808
rect 1506 5765 1514 5799
rect 1514 5765 1548 5799
rect 1548 5765 1558 5799
rect 1506 5756 1558 5765
rect 1570 5799 1622 5808
rect 1570 5765 1586 5799
rect 1586 5765 1620 5799
rect 1620 5765 1622 5799
rect 1570 5756 1622 5765
rect 1634 5799 1686 5808
rect 1698 5799 1750 5808
rect 1762 5799 1814 5808
rect 1826 5799 1878 5808
rect 1890 5799 1942 5808
rect 1954 5799 2006 5808
rect 1634 5765 1658 5799
rect 1658 5765 1686 5799
rect 1698 5765 1730 5799
rect 1730 5765 1750 5799
rect 1762 5765 1764 5799
rect 1764 5765 1802 5799
rect 1802 5765 1814 5799
rect 1826 5765 1836 5799
rect 1836 5765 1874 5799
rect 1874 5765 1878 5799
rect 1890 5765 1908 5799
rect 1908 5765 1942 5799
rect 1954 5765 1980 5799
rect 1980 5765 2006 5799
rect 1634 5756 1686 5765
rect 1698 5756 1750 5765
rect 1762 5756 1814 5765
rect 1826 5756 1878 5765
rect 1890 5756 1942 5765
rect 1954 5756 2006 5765
rect 2018 5799 2070 5808
rect 2018 5765 2052 5799
rect 2052 5765 2070 5799
rect 2018 5756 2070 5765
rect 2082 5799 2134 5808
rect 2082 5765 2090 5799
rect 2090 5765 2124 5799
rect 2124 5765 2134 5799
rect 2082 5756 2134 5765
rect 2146 5799 2198 5808
rect 2146 5765 2162 5799
rect 2162 5765 2196 5799
rect 2196 5765 2198 5799
rect 2146 5756 2198 5765
rect 2210 5799 2262 5808
rect 2274 5799 2326 5808
rect 2338 5799 2390 5808
rect 2402 5799 2454 5808
rect 2466 5799 2518 5808
rect 2530 5799 2582 5808
rect 2210 5765 2234 5799
rect 2234 5765 2262 5799
rect 2274 5765 2306 5799
rect 2306 5765 2326 5799
rect 2338 5765 2340 5799
rect 2340 5765 2378 5799
rect 2378 5765 2390 5799
rect 2402 5765 2412 5799
rect 2412 5765 2450 5799
rect 2450 5765 2454 5799
rect 2466 5765 2484 5799
rect 2484 5765 2518 5799
rect 2530 5765 2556 5799
rect 2556 5765 2582 5799
rect 2210 5756 2262 5765
rect 2274 5756 2326 5765
rect 2338 5756 2390 5765
rect 2402 5756 2454 5765
rect 2466 5756 2518 5765
rect 2530 5756 2582 5765
rect 2594 5799 2646 5808
rect 2594 5765 2628 5799
rect 2628 5765 2646 5799
rect 2594 5756 2646 5765
rect 2658 5799 2710 5808
rect 2658 5765 2666 5799
rect 2666 5765 2700 5799
rect 2700 5765 2710 5799
rect 2658 5756 2710 5765
rect 2722 5799 2774 5808
rect 2722 5765 2738 5799
rect 2738 5765 2772 5799
rect 2772 5765 2774 5799
rect 2722 5756 2774 5765
rect 2786 5799 2838 5808
rect 2850 5799 2902 5808
rect 2914 5799 2966 5808
rect 2978 5799 3030 5808
rect 3042 5799 3094 5808
rect 3106 5799 3158 5808
rect 2786 5765 2810 5799
rect 2810 5765 2838 5799
rect 2850 5765 2882 5799
rect 2882 5765 2902 5799
rect 2914 5765 2916 5799
rect 2916 5765 2954 5799
rect 2954 5765 2966 5799
rect 2978 5765 2988 5799
rect 2988 5765 3026 5799
rect 3026 5765 3030 5799
rect 3042 5765 3060 5799
rect 3060 5765 3094 5799
rect 3106 5765 3132 5799
rect 3132 5765 3158 5799
rect 2786 5756 2838 5765
rect 2850 5756 2902 5765
rect 2914 5756 2966 5765
rect 2978 5756 3030 5765
rect 3042 5756 3094 5765
rect 3106 5756 3158 5765
rect 3170 5799 3222 5808
rect 3170 5765 3204 5799
rect 3204 5765 3222 5799
rect 3170 5756 3222 5765
rect 3234 5799 3286 5808
rect 3234 5765 3242 5799
rect 3242 5765 3276 5799
rect 3276 5765 3286 5799
rect 3234 5756 3286 5765
rect 3298 5799 3350 5808
rect 3298 5765 3314 5799
rect 3314 5765 3348 5799
rect 3348 5765 3350 5799
rect 3298 5756 3350 5765
rect 3362 5799 3414 5808
rect 3427 5799 3479 5808
rect 3492 5799 3544 5808
rect 3557 5799 3609 5808
rect 3622 5799 3674 5808
rect 3687 5799 3739 5808
rect 3752 5799 3804 5808
rect 3362 5765 3386 5799
rect 3386 5765 3414 5799
rect 3427 5765 3458 5799
rect 3458 5765 3479 5799
rect 3492 5765 3530 5799
rect 3530 5765 3544 5799
rect 3557 5765 3564 5799
rect 3564 5765 3602 5799
rect 3602 5765 3609 5799
rect 3622 5765 3636 5799
rect 3636 5765 3674 5799
rect 3687 5765 3708 5799
rect 3708 5765 3739 5799
rect 3752 5765 3780 5799
rect 3780 5765 3804 5799
rect 3362 5756 3414 5765
rect 3427 5756 3479 5765
rect 3492 5756 3544 5765
rect 3557 5756 3609 5765
rect 3622 5756 3674 5765
rect 3687 5756 3739 5765
rect 3752 5756 3804 5765
rect 3817 5799 3869 5808
rect 3817 5765 3818 5799
rect 3818 5765 3852 5799
rect 3852 5765 3869 5799
rect 3817 5756 3869 5765
rect 3882 5799 3934 5808
rect 3882 5765 3890 5799
rect 3890 5765 3924 5799
rect 3924 5765 3934 5799
rect 3882 5756 3934 5765
rect 3947 5799 3999 5808
rect 3947 5765 3962 5799
rect 3962 5765 3996 5799
rect 3996 5765 3999 5799
rect 3947 5756 3999 5765
rect 4012 5799 4064 5808
rect 4077 5799 4129 5808
rect 4142 5799 4194 5808
rect 4207 5799 4259 5808
rect 4272 5799 4324 5808
rect 4337 5799 4389 5808
rect 4402 5799 4454 5808
rect 4467 5799 4519 5808
rect 4012 5765 4034 5799
rect 4034 5765 4064 5799
rect 4077 5765 4106 5799
rect 4106 5765 4129 5799
rect 4142 5765 4178 5799
rect 4178 5765 4194 5799
rect 4207 5765 4212 5799
rect 4212 5765 4250 5799
rect 4250 5765 4259 5799
rect 4272 5765 4284 5799
rect 4284 5765 4322 5799
rect 4322 5765 4324 5799
rect 4337 5765 4356 5799
rect 4356 5765 4389 5799
rect 4402 5765 4428 5799
rect 4428 5765 4454 5799
rect 4467 5765 4500 5799
rect 4500 5765 4519 5799
rect 4012 5756 4064 5765
rect 4077 5756 4129 5765
rect 4142 5756 4194 5765
rect 4207 5756 4259 5765
rect 4272 5756 4324 5765
rect 4337 5756 4389 5765
rect 4402 5756 4454 5765
rect 4467 5756 4519 5765
rect 4532 5799 4584 5808
rect 4532 5765 4538 5799
rect 4538 5765 4572 5799
rect 4572 5765 4584 5799
rect 4532 5756 4584 5765
rect 4597 5799 4649 5808
rect 4597 5765 4610 5799
rect 4610 5765 4644 5799
rect 4644 5765 4649 5799
rect 4597 5756 4649 5765
rect 4662 5799 4714 5808
rect 4727 5799 4779 5808
rect 4792 5799 4844 5808
rect 4857 5799 4909 5808
rect 4922 5799 4974 5808
rect 4987 5799 5039 5808
rect 5052 5799 5104 5808
rect 5117 5799 5169 5808
rect 4662 5765 4682 5799
rect 4682 5765 4714 5799
rect 4727 5765 4754 5799
rect 4754 5765 4779 5799
rect 4792 5765 4826 5799
rect 4826 5765 4844 5799
rect 4857 5765 4860 5799
rect 4860 5765 4898 5799
rect 4898 5765 4909 5799
rect 4922 5765 4932 5799
rect 4932 5765 4970 5799
rect 4970 5765 4974 5799
rect 4987 5765 5004 5799
rect 5004 5765 5039 5799
rect 5052 5765 5076 5799
rect 5076 5765 5104 5799
rect 5117 5765 5148 5799
rect 5148 5765 5169 5799
rect 4662 5756 4714 5765
rect 4727 5756 4779 5765
rect 4792 5756 4844 5765
rect 4857 5756 4909 5765
rect 4922 5756 4974 5765
rect 4987 5756 5039 5765
rect 5052 5756 5104 5765
rect 5117 5756 5169 5765
rect 5182 5799 5234 5808
rect 5182 5765 5186 5799
rect 5186 5765 5220 5799
rect 5220 5765 5234 5799
rect 5182 5756 5234 5765
rect 5247 5799 5299 5808
rect 5247 5765 5258 5799
rect 5258 5765 5292 5799
rect 5292 5765 5299 5799
rect 5247 5756 5299 5765
rect 5312 5799 5364 5808
rect 5312 5765 5330 5799
rect 5330 5765 5364 5799
rect 5312 5756 5364 5765
rect 5377 5799 5429 5808
rect 5442 5799 5494 5808
rect 5507 5799 5559 5808
rect 5572 5799 5624 5808
rect 5637 5799 5689 5808
rect 5702 5799 5754 5808
rect 5767 5799 5819 5808
rect 5377 5765 5402 5799
rect 5402 5765 5429 5799
rect 5442 5765 5474 5799
rect 5474 5765 5494 5799
rect 5507 5765 5508 5799
rect 5508 5765 5546 5799
rect 5546 5765 5559 5799
rect 5572 5765 5580 5799
rect 5580 5765 5618 5799
rect 5618 5765 5624 5799
rect 5637 5765 5652 5799
rect 5652 5765 5689 5799
rect 5702 5765 5724 5799
rect 5724 5765 5754 5799
rect 5767 5765 5797 5799
rect 5797 5765 5819 5799
rect 5377 5756 5429 5765
rect 5442 5756 5494 5765
rect 5507 5756 5559 5765
rect 5572 5756 5624 5765
rect 5637 5756 5689 5765
rect 5702 5756 5754 5765
rect 5767 5756 5819 5765
rect 5832 5799 5884 5808
rect 5832 5765 5836 5799
rect 5836 5765 5870 5799
rect 5870 5765 5884 5799
rect 5832 5756 5884 5765
rect 5897 5799 5949 5808
rect 5897 5765 5909 5799
rect 5909 5765 5943 5799
rect 5943 5765 5949 5799
rect 5897 5756 5949 5765
rect 351 5371 360 5402
rect 360 5371 394 5402
rect 394 5371 403 5402
rect 351 5350 403 5371
rect 351 5333 403 5338
rect 351 5299 360 5333
rect 360 5299 394 5333
rect 394 5299 403 5333
rect 351 5286 403 5299
rect 351 5261 403 5274
rect 351 5227 360 5261
rect 360 5227 394 5261
rect 394 5227 403 5261
rect 351 5222 403 5227
rect 351 5189 403 5210
rect 351 5158 360 5189
rect 360 5158 394 5189
rect 394 5158 403 5189
rect 351 5117 403 5146
rect 351 5094 360 5117
rect 360 5094 394 5117
rect 394 5094 403 5117
rect 351 5045 403 5082
rect 351 5030 360 5045
rect 360 5030 394 5045
rect 394 5030 403 5045
rect 351 5011 360 5018
rect 360 5011 394 5018
rect 394 5011 403 5018
rect 351 4973 403 5011
rect 351 4966 360 4973
rect 360 4966 394 4973
rect 394 4966 403 4973
rect 351 4939 360 4954
rect 360 4939 394 4954
rect 394 4939 403 4954
rect 351 4902 403 4939
rect 351 4867 360 4890
rect 360 4867 394 4890
rect 394 4867 403 4890
rect 351 4838 403 4867
rect 351 4795 360 4826
rect 360 4795 394 4826
rect 394 4795 403 4826
rect 351 4774 403 4795
rect 351 4757 403 4762
rect 351 4723 360 4757
rect 360 4723 394 4757
rect 394 4723 403 4757
rect 351 4710 403 4723
rect 351 4685 403 4698
rect 351 4651 360 4685
rect 360 4651 394 4685
rect 394 4651 403 4685
rect 351 4646 403 4651
rect 351 4613 403 4634
rect 351 4582 360 4613
rect 360 4582 394 4613
rect 394 4582 403 4613
rect 351 4541 403 4570
rect 351 4518 360 4541
rect 360 4518 394 4541
rect 394 4518 403 4541
rect 471 5377 480 5402
rect 480 5377 514 5402
rect 514 5377 523 5402
rect 471 5350 523 5377
rect 471 5305 480 5338
rect 480 5305 514 5338
rect 514 5305 523 5338
rect 471 5286 523 5305
rect 471 5267 523 5274
rect 471 5233 480 5267
rect 480 5233 514 5267
rect 514 5233 523 5267
rect 471 5222 523 5233
rect 471 5195 523 5210
rect 471 5161 480 5195
rect 480 5161 514 5195
rect 514 5161 523 5195
rect 471 5158 523 5161
rect 471 5123 523 5146
rect 471 5094 480 5123
rect 480 5094 514 5123
rect 514 5094 523 5123
rect 471 5051 523 5082
rect 471 5030 480 5051
rect 480 5030 514 5051
rect 514 5030 523 5051
rect 471 5017 480 5018
rect 480 5017 514 5018
rect 514 5017 523 5018
rect 471 4979 523 5017
rect 471 4966 480 4979
rect 480 4966 514 4979
rect 514 4966 523 4979
rect 471 4945 480 4954
rect 480 4945 514 4954
rect 514 4945 523 4954
rect 471 4907 523 4945
rect 471 4902 480 4907
rect 480 4902 514 4907
rect 514 4902 523 4907
rect 471 4873 480 4890
rect 480 4873 514 4890
rect 514 4873 523 4890
rect 471 4838 523 4873
rect 471 4801 480 4826
rect 480 4801 514 4826
rect 514 4801 523 4826
rect 471 4774 523 4801
rect 471 4729 480 4762
rect 480 4729 514 4762
rect 514 4729 523 4762
rect 471 4710 523 4729
rect 471 4691 523 4698
rect 471 4657 480 4691
rect 480 4657 514 4691
rect 514 4657 523 4691
rect 471 4646 523 4657
rect 471 4619 523 4634
rect 471 4585 480 4619
rect 480 4585 514 4619
rect 514 4585 523 4619
rect 471 4582 523 4585
rect 471 4547 523 4570
rect 471 4518 480 4547
rect 480 4518 514 4547
rect 514 4518 523 4547
rect 1327 5377 1336 5402
rect 1336 5377 1370 5402
rect 1370 5377 1379 5402
rect 1327 5350 1379 5377
rect 1327 5305 1336 5338
rect 1336 5305 1370 5338
rect 1370 5305 1379 5338
rect 1327 5286 1379 5305
rect 1327 5267 1379 5274
rect 1327 5233 1336 5267
rect 1336 5233 1370 5267
rect 1370 5233 1379 5267
rect 1327 5222 1379 5233
rect 1327 5195 1379 5210
rect 1327 5161 1336 5195
rect 1336 5161 1370 5195
rect 1370 5161 1379 5195
rect 1327 5158 1379 5161
rect 1327 5123 1379 5146
rect 1327 5094 1336 5123
rect 1336 5094 1370 5123
rect 1370 5094 1379 5123
rect 1327 5051 1379 5082
rect 1327 5030 1336 5051
rect 1336 5030 1370 5051
rect 1370 5030 1379 5051
rect 1327 5017 1336 5018
rect 1336 5017 1370 5018
rect 1370 5017 1379 5018
rect 1327 4979 1379 5017
rect 1327 4966 1336 4979
rect 1336 4966 1370 4979
rect 1370 4966 1379 4979
rect 1327 4945 1336 4954
rect 1336 4945 1370 4954
rect 1370 4945 1379 4954
rect 1327 4907 1379 4945
rect 1327 4902 1336 4907
rect 1336 4902 1370 4907
rect 1370 4902 1379 4907
rect 1327 4873 1336 4890
rect 1336 4873 1370 4890
rect 1370 4873 1379 4890
rect 1327 4838 1379 4873
rect 1327 4801 1336 4826
rect 1336 4801 1370 4826
rect 1370 4801 1379 4826
rect 1327 4774 1379 4801
rect 1327 4729 1336 4762
rect 1336 4729 1370 4762
rect 1370 4729 1379 4762
rect 1327 4710 1379 4729
rect 1327 4691 1379 4698
rect 1327 4657 1336 4691
rect 1336 4657 1370 4691
rect 1370 4657 1379 4691
rect 1327 4646 1379 4657
rect 1327 4619 1379 4634
rect 1327 4585 1336 4619
rect 1336 4585 1370 4619
rect 1370 4585 1379 4619
rect 1327 4582 1379 4585
rect 1327 4547 1379 4570
rect 1327 4518 1336 4547
rect 1336 4518 1370 4547
rect 1370 4518 1379 4547
rect 2183 5377 2192 5402
rect 2192 5377 2226 5402
rect 2226 5377 2235 5402
rect 2183 5350 2235 5377
rect 2183 5305 2192 5338
rect 2192 5305 2226 5338
rect 2226 5305 2235 5338
rect 2183 5286 2235 5305
rect 2183 5267 2235 5274
rect 2183 5233 2192 5267
rect 2192 5233 2226 5267
rect 2226 5233 2235 5267
rect 2183 5222 2235 5233
rect 2183 5195 2235 5210
rect 2183 5161 2192 5195
rect 2192 5161 2226 5195
rect 2226 5161 2235 5195
rect 2183 5158 2235 5161
rect 2183 5123 2235 5146
rect 2183 5094 2192 5123
rect 2192 5094 2226 5123
rect 2226 5094 2235 5123
rect 2183 5051 2235 5082
rect 2183 5030 2192 5051
rect 2192 5030 2226 5051
rect 2226 5030 2235 5051
rect 2183 5017 2192 5018
rect 2192 5017 2226 5018
rect 2226 5017 2235 5018
rect 2183 4979 2235 5017
rect 2183 4966 2192 4979
rect 2192 4966 2226 4979
rect 2226 4966 2235 4979
rect 2183 4945 2192 4954
rect 2192 4945 2226 4954
rect 2226 4945 2235 4954
rect 2183 4907 2235 4945
rect 2183 4902 2192 4907
rect 2192 4902 2226 4907
rect 2226 4902 2235 4907
rect 2183 4873 2192 4890
rect 2192 4873 2226 4890
rect 2226 4873 2235 4890
rect 2183 4838 2235 4873
rect 2183 4801 2192 4826
rect 2192 4801 2226 4826
rect 2226 4801 2235 4826
rect 2183 4774 2235 4801
rect 2183 4729 2192 4762
rect 2192 4729 2226 4762
rect 2226 4729 2235 4762
rect 2183 4710 2235 4729
rect 2183 4691 2235 4698
rect 2183 4657 2192 4691
rect 2192 4657 2226 4691
rect 2226 4657 2235 4691
rect 2183 4646 2235 4657
rect 2183 4619 2235 4634
rect 2183 4585 2192 4619
rect 2192 4585 2226 4619
rect 2226 4585 2235 4619
rect 2183 4582 2235 4585
rect 2183 4547 2235 4570
rect 2183 4518 2192 4547
rect 2192 4518 2226 4547
rect 2226 4518 2235 4547
rect 3039 5377 3048 5402
rect 3048 5377 3082 5402
rect 3082 5377 3091 5402
rect 3039 5350 3091 5377
rect 3039 5305 3048 5338
rect 3048 5305 3082 5338
rect 3082 5305 3091 5338
rect 3039 5286 3091 5305
rect 3039 5267 3091 5274
rect 3039 5233 3048 5267
rect 3048 5233 3082 5267
rect 3082 5233 3091 5267
rect 3039 5222 3091 5233
rect 3039 5195 3091 5210
rect 3039 5161 3048 5195
rect 3048 5161 3082 5195
rect 3082 5161 3091 5195
rect 3039 5158 3091 5161
rect 3039 5123 3091 5146
rect 3039 5094 3048 5123
rect 3048 5094 3082 5123
rect 3082 5094 3091 5123
rect 3039 5051 3091 5082
rect 3039 5030 3048 5051
rect 3048 5030 3082 5051
rect 3082 5030 3091 5051
rect 3039 5017 3048 5018
rect 3048 5017 3082 5018
rect 3082 5017 3091 5018
rect 3039 4979 3091 5017
rect 3039 4966 3048 4979
rect 3048 4966 3082 4979
rect 3082 4966 3091 4979
rect 3039 4945 3048 4954
rect 3048 4945 3082 4954
rect 3082 4945 3091 4954
rect 3039 4907 3091 4945
rect 3039 4902 3048 4907
rect 3048 4902 3082 4907
rect 3082 4902 3091 4907
rect 3039 4873 3048 4890
rect 3048 4873 3082 4890
rect 3082 4873 3091 4890
rect 3039 4838 3091 4873
rect 3039 4801 3048 4826
rect 3048 4801 3082 4826
rect 3082 4801 3091 4826
rect 3039 4774 3091 4801
rect 3039 4729 3048 4762
rect 3048 4729 3082 4762
rect 3082 4729 3091 4762
rect 3039 4710 3091 4729
rect 3039 4691 3091 4698
rect 3039 4657 3048 4691
rect 3048 4657 3082 4691
rect 3082 4657 3091 4691
rect 3039 4646 3091 4657
rect 3039 4619 3091 4634
rect 3039 4585 3048 4619
rect 3048 4585 3082 4619
rect 3082 4585 3091 4619
rect 3039 4582 3091 4585
rect 3039 4547 3091 4570
rect 3039 4518 3048 4547
rect 3048 4518 3082 4547
rect 3082 4518 3091 4547
rect 3895 5377 3904 5402
rect 3904 5377 3938 5402
rect 3938 5377 3947 5402
rect 3895 5350 3947 5377
rect 3895 5305 3904 5338
rect 3904 5305 3938 5338
rect 3938 5305 3947 5338
rect 3895 5286 3947 5305
rect 3895 5267 3947 5274
rect 3895 5233 3904 5267
rect 3904 5233 3938 5267
rect 3938 5233 3947 5267
rect 3895 5222 3947 5233
rect 3895 5195 3947 5210
rect 3895 5161 3904 5195
rect 3904 5161 3938 5195
rect 3938 5161 3947 5195
rect 3895 5158 3947 5161
rect 3895 5123 3947 5146
rect 3895 5094 3904 5123
rect 3904 5094 3938 5123
rect 3938 5094 3947 5123
rect 3895 5051 3947 5082
rect 3895 5030 3904 5051
rect 3904 5030 3938 5051
rect 3938 5030 3947 5051
rect 3895 5017 3904 5018
rect 3904 5017 3938 5018
rect 3938 5017 3947 5018
rect 3895 4979 3947 5017
rect 3895 4966 3904 4979
rect 3904 4966 3938 4979
rect 3938 4966 3947 4979
rect 3895 4945 3904 4954
rect 3904 4945 3938 4954
rect 3938 4945 3947 4954
rect 3895 4907 3947 4945
rect 3895 4902 3904 4907
rect 3904 4902 3938 4907
rect 3938 4902 3947 4907
rect 3895 4873 3904 4890
rect 3904 4873 3938 4890
rect 3938 4873 3947 4890
rect 3895 4838 3947 4873
rect 3895 4801 3904 4826
rect 3904 4801 3938 4826
rect 3938 4801 3947 4826
rect 3895 4774 3947 4801
rect 3895 4729 3904 4762
rect 3904 4729 3938 4762
rect 3938 4729 3947 4762
rect 3895 4710 3947 4729
rect 3895 4691 3947 4698
rect 3895 4657 3904 4691
rect 3904 4657 3938 4691
rect 3938 4657 3947 4691
rect 3895 4646 3947 4657
rect 3895 4619 3947 4634
rect 3895 4585 3904 4619
rect 3904 4585 3938 4619
rect 3938 4585 3947 4619
rect 3895 4582 3947 4585
rect 3895 4547 3947 4570
rect 3895 4518 3904 4547
rect 3904 4518 3938 4547
rect 3938 4518 3947 4547
rect 4751 5377 4760 5402
rect 4760 5377 4794 5402
rect 4794 5377 4803 5402
rect 4751 5350 4803 5377
rect 4751 5305 4760 5338
rect 4760 5305 4794 5338
rect 4794 5305 4803 5338
rect 4751 5286 4803 5305
rect 4751 5267 4803 5274
rect 4751 5233 4760 5267
rect 4760 5233 4794 5267
rect 4794 5233 4803 5267
rect 4751 5222 4803 5233
rect 4751 5195 4803 5210
rect 4751 5161 4760 5195
rect 4760 5161 4794 5195
rect 4794 5161 4803 5195
rect 4751 5158 4803 5161
rect 4751 5123 4803 5146
rect 4751 5094 4760 5123
rect 4760 5094 4794 5123
rect 4794 5094 4803 5123
rect 4751 5051 4803 5082
rect 4751 5030 4760 5051
rect 4760 5030 4794 5051
rect 4794 5030 4803 5051
rect 4751 5017 4760 5018
rect 4760 5017 4794 5018
rect 4794 5017 4803 5018
rect 4751 4979 4803 5017
rect 4751 4966 4760 4979
rect 4760 4966 4794 4979
rect 4794 4966 4803 4979
rect 4751 4945 4760 4954
rect 4760 4945 4794 4954
rect 4794 4945 4803 4954
rect 4751 4907 4803 4945
rect 4751 4902 4760 4907
rect 4760 4902 4794 4907
rect 4794 4902 4803 4907
rect 4751 4873 4760 4890
rect 4760 4873 4794 4890
rect 4794 4873 4803 4890
rect 4751 4838 4803 4873
rect 4751 4801 4760 4826
rect 4760 4801 4794 4826
rect 4794 4801 4803 4826
rect 4751 4774 4803 4801
rect 4751 4729 4760 4762
rect 4760 4729 4794 4762
rect 4794 4729 4803 4762
rect 4751 4710 4803 4729
rect 4751 4691 4803 4698
rect 4751 4657 4760 4691
rect 4760 4657 4794 4691
rect 4794 4657 4803 4691
rect 4751 4646 4803 4657
rect 4751 4619 4803 4634
rect 4751 4585 4760 4619
rect 4760 4585 4794 4619
rect 4794 4585 4803 4619
rect 4751 4582 4803 4585
rect 4751 4547 4803 4570
rect 4751 4518 4760 4547
rect 4760 4518 4794 4547
rect 4794 4518 4803 4547
rect 5607 5377 5616 5402
rect 5616 5377 5650 5402
rect 5650 5377 5659 5402
rect 5607 5350 5659 5377
rect 5607 5305 5616 5338
rect 5616 5305 5650 5338
rect 5650 5305 5659 5338
rect 5607 5286 5659 5305
rect 5607 5267 5659 5274
rect 5607 5233 5616 5267
rect 5616 5233 5650 5267
rect 5650 5233 5659 5267
rect 5607 5222 5659 5233
rect 5607 5195 5659 5210
rect 5607 5161 5616 5195
rect 5616 5161 5650 5195
rect 5650 5161 5659 5195
rect 5607 5158 5659 5161
rect 5607 5123 5659 5146
rect 5607 5094 5616 5123
rect 5616 5094 5650 5123
rect 5650 5094 5659 5123
rect 5607 5051 5659 5082
rect 5607 5030 5616 5051
rect 5616 5030 5650 5051
rect 5650 5030 5659 5051
rect 5607 5017 5616 5018
rect 5616 5017 5650 5018
rect 5650 5017 5659 5018
rect 5607 4979 5659 5017
rect 5607 4966 5616 4979
rect 5616 4966 5650 4979
rect 5650 4966 5659 4979
rect 5607 4945 5616 4954
rect 5616 4945 5650 4954
rect 5650 4945 5659 4954
rect 5607 4907 5659 4945
rect 5607 4902 5616 4907
rect 5616 4902 5650 4907
rect 5650 4902 5659 4907
rect 5607 4873 5616 4890
rect 5616 4873 5650 4890
rect 5650 4873 5659 4890
rect 5607 4838 5659 4873
rect 5607 4801 5616 4826
rect 5616 4801 5650 4826
rect 5650 4801 5659 4826
rect 5607 4774 5659 4801
rect 5607 4729 5616 4762
rect 5616 4729 5650 4762
rect 5650 4729 5659 4762
rect 5607 4710 5659 4729
rect 5607 4691 5659 4698
rect 5607 4657 5616 4691
rect 5616 4657 5650 4691
rect 5650 4657 5659 4691
rect 5607 4646 5659 4657
rect 5607 4619 5659 4634
rect 5607 4585 5616 4619
rect 5616 4585 5650 4619
rect 5650 4585 5659 4619
rect 5607 4582 5659 4585
rect 5607 4547 5659 4570
rect 5607 4518 5616 4547
rect 5616 4518 5650 4547
rect 5650 4518 5659 4547
rect 6189 6033 6241 6042
rect 6189 5999 6195 6033
rect 6195 5999 6229 6033
rect 6229 5999 6241 6033
rect 6189 5990 6241 5999
rect 6254 6033 6306 6042
rect 6254 5999 6269 6033
rect 6269 5999 6303 6033
rect 6303 5999 6306 6033
rect 6254 5990 6306 5999
rect 6319 6033 6371 6042
rect 6384 6033 6436 6042
rect 6448 6033 6500 6042
rect 6512 6033 6564 6042
rect 6576 6033 6628 6042
rect 6640 6033 6692 6042
rect 6319 5999 6342 6033
rect 6342 5999 6371 6033
rect 6384 5999 6415 6033
rect 6415 5999 6436 6033
rect 6448 5999 6449 6033
rect 6449 5999 6488 6033
rect 6488 5999 6500 6033
rect 6512 5999 6522 6033
rect 6522 5999 6561 6033
rect 6561 5999 6564 6033
rect 6576 5999 6595 6033
rect 6595 5999 6628 6033
rect 6640 5999 6668 6033
rect 6668 5999 6692 6033
rect 6319 5990 6371 5999
rect 6384 5990 6436 5999
rect 6448 5990 6500 5999
rect 6512 5990 6564 5999
rect 6576 5990 6628 5999
rect 6640 5990 6692 5999
rect 6704 6033 6756 6042
rect 6704 5999 6707 6033
rect 6707 5999 6741 6033
rect 6741 5999 6756 6033
rect 6704 5990 6756 5999
rect 6768 6033 6820 6042
rect 6768 5999 6780 6033
rect 6780 5999 6814 6033
rect 6814 5999 6820 6033
rect 6768 5990 6820 5999
rect 6189 5799 6241 5808
rect 6189 5765 6195 5799
rect 6195 5765 6229 5799
rect 6229 5765 6241 5799
rect 6189 5756 6241 5765
rect 6254 5799 6306 5808
rect 6254 5765 6269 5799
rect 6269 5765 6303 5799
rect 6303 5765 6306 5799
rect 6254 5756 6306 5765
rect 6319 5799 6371 5808
rect 6384 5799 6436 5808
rect 6448 5799 6500 5808
rect 6512 5799 6564 5808
rect 6576 5799 6628 5808
rect 6640 5799 6692 5808
rect 6319 5765 6342 5799
rect 6342 5765 6371 5799
rect 6384 5765 6415 5799
rect 6415 5765 6436 5799
rect 6448 5765 6449 5799
rect 6449 5765 6488 5799
rect 6488 5765 6500 5799
rect 6512 5765 6522 5799
rect 6522 5765 6561 5799
rect 6561 5765 6564 5799
rect 6576 5765 6595 5799
rect 6595 5765 6628 5799
rect 6640 5765 6668 5799
rect 6668 5765 6692 5799
rect 6319 5756 6371 5765
rect 6384 5756 6436 5765
rect 6448 5756 6500 5765
rect 6512 5756 6564 5765
rect 6576 5756 6628 5765
rect 6640 5756 6692 5765
rect 6704 5799 6756 5808
rect 6704 5765 6707 5799
rect 6707 5765 6741 5799
rect 6741 5765 6756 5799
rect 6704 5756 6756 5765
rect 6768 5799 6820 5808
rect 6768 5765 6780 5799
rect 6780 5765 6814 5799
rect 6814 5765 6820 5799
rect 6768 5756 6820 5765
rect 6463 5377 6472 5402
rect 6472 5377 6506 5402
rect 6506 5377 6515 5402
rect 6463 5350 6515 5377
rect 6463 5305 6472 5338
rect 6472 5305 6506 5338
rect 6506 5305 6515 5338
rect 6463 5286 6515 5305
rect 6463 5267 6515 5274
rect 6463 5233 6472 5267
rect 6472 5233 6506 5267
rect 6506 5233 6515 5267
rect 6463 5222 6515 5233
rect 6463 5195 6515 5210
rect 6463 5161 6472 5195
rect 6472 5161 6506 5195
rect 6506 5161 6515 5195
rect 6463 5158 6515 5161
rect 6463 5123 6515 5146
rect 6463 5094 6472 5123
rect 6472 5094 6506 5123
rect 6506 5094 6515 5123
rect 6463 5051 6515 5082
rect 6463 5030 6472 5051
rect 6472 5030 6506 5051
rect 6506 5030 6515 5051
rect 6463 5017 6472 5018
rect 6472 5017 6506 5018
rect 6506 5017 6515 5018
rect 6463 4979 6515 5017
rect 6463 4966 6472 4979
rect 6472 4966 6506 4979
rect 6506 4966 6515 4979
rect 6463 4945 6472 4954
rect 6472 4945 6506 4954
rect 6506 4945 6515 4954
rect 6463 4907 6515 4945
rect 6463 4902 6472 4907
rect 6472 4902 6506 4907
rect 6506 4902 6515 4907
rect 6463 4873 6472 4890
rect 6472 4873 6506 4890
rect 6506 4873 6515 4890
rect 6463 4838 6515 4873
rect 6463 4801 6472 4826
rect 6472 4801 6506 4826
rect 6506 4801 6515 4826
rect 6463 4774 6515 4801
rect 6463 4729 6472 4762
rect 6472 4729 6506 4762
rect 6506 4729 6515 4762
rect 6463 4710 6515 4729
rect 6463 4691 6515 4698
rect 6463 4657 6472 4691
rect 6472 4657 6506 4691
rect 6506 4657 6515 4691
rect 6463 4646 6515 4657
rect 6463 4619 6515 4634
rect 6463 4585 6472 4619
rect 6472 4585 6506 4619
rect 6506 4585 6515 4619
rect 6463 4582 6515 4585
rect 6463 4547 6515 4570
rect 6463 4518 6472 4547
rect 6472 4518 6506 4547
rect 6506 4518 6515 4547
rect 7060 6033 7112 6042
rect 7060 5999 7069 6033
rect 7069 5999 7103 6033
rect 7103 5999 7112 6033
rect 7060 5990 7112 5999
rect 7124 6033 7176 6042
rect 7124 5999 7141 6033
rect 7141 5999 7175 6033
rect 7175 5999 7176 6033
rect 7124 5990 7176 5999
rect 7188 6033 7240 6042
rect 7252 6033 7304 6042
rect 7316 6033 7368 6042
rect 7380 6033 7432 6042
rect 7444 6033 7496 6042
rect 7508 6033 7560 6042
rect 7188 5999 7213 6033
rect 7213 5999 7240 6033
rect 7252 5999 7285 6033
rect 7285 5999 7304 6033
rect 7316 5999 7319 6033
rect 7319 5999 7357 6033
rect 7357 5999 7368 6033
rect 7380 5999 7391 6033
rect 7391 5999 7429 6033
rect 7429 5999 7432 6033
rect 7444 5999 7463 6033
rect 7463 5999 7496 6033
rect 7508 5999 7535 6033
rect 7535 5999 7560 6033
rect 7188 5990 7240 5999
rect 7252 5990 7304 5999
rect 7316 5990 7368 5999
rect 7380 5990 7432 5999
rect 7444 5990 7496 5999
rect 7508 5990 7560 5999
rect 7572 6033 7624 6042
rect 7572 5999 7573 6033
rect 7573 5999 7607 6033
rect 7607 5999 7624 6033
rect 7572 5990 7624 5999
rect 7060 5799 7112 5808
rect 7060 5765 7069 5799
rect 7069 5765 7103 5799
rect 7103 5765 7112 5799
rect 7060 5756 7112 5765
rect 7124 5799 7176 5808
rect 7124 5765 7141 5799
rect 7141 5765 7175 5799
rect 7175 5765 7176 5799
rect 7124 5756 7176 5765
rect 7188 5799 7240 5808
rect 7252 5799 7304 5808
rect 7316 5799 7368 5808
rect 7380 5799 7432 5808
rect 7444 5799 7496 5808
rect 7508 5799 7560 5808
rect 7188 5765 7213 5799
rect 7213 5765 7240 5799
rect 7252 5765 7285 5799
rect 7285 5765 7304 5799
rect 7316 5765 7319 5799
rect 7319 5765 7357 5799
rect 7357 5765 7368 5799
rect 7380 5765 7391 5799
rect 7391 5765 7429 5799
rect 7429 5765 7432 5799
rect 7444 5765 7463 5799
rect 7463 5765 7496 5799
rect 7508 5765 7535 5799
rect 7535 5765 7560 5799
rect 7188 5756 7240 5765
rect 7252 5756 7304 5765
rect 7316 5756 7368 5765
rect 7380 5756 7432 5765
rect 7444 5756 7496 5765
rect 7508 5756 7560 5765
rect 7572 5799 7624 5808
rect 7572 5765 7573 5799
rect 7573 5765 7607 5799
rect 7607 5765 7624 5799
rect 7572 5756 7624 5765
rect 7319 5377 7328 5402
rect 7328 5377 7362 5402
rect 7362 5377 7371 5402
rect 7319 5350 7371 5377
rect 7319 5305 7328 5338
rect 7328 5305 7362 5338
rect 7362 5305 7371 5338
rect 7319 5286 7371 5305
rect 7319 5267 7371 5274
rect 7319 5233 7328 5267
rect 7328 5233 7362 5267
rect 7362 5233 7371 5267
rect 7319 5222 7371 5233
rect 7319 5195 7371 5210
rect 7319 5161 7328 5195
rect 7328 5161 7362 5195
rect 7362 5161 7371 5195
rect 7319 5158 7371 5161
rect 7319 5123 7371 5146
rect 7319 5094 7328 5123
rect 7328 5094 7362 5123
rect 7362 5094 7371 5123
rect 7319 5051 7371 5082
rect 7319 5030 7328 5051
rect 7328 5030 7362 5051
rect 7362 5030 7371 5051
rect 7319 5017 7328 5018
rect 7328 5017 7362 5018
rect 7362 5017 7371 5018
rect 7319 4979 7371 5017
rect 7319 4966 7328 4979
rect 7328 4966 7362 4979
rect 7362 4966 7371 4979
rect 7319 4945 7328 4954
rect 7328 4945 7362 4954
rect 7362 4945 7371 4954
rect 7319 4907 7371 4945
rect 7319 4902 7328 4907
rect 7328 4902 7362 4907
rect 7362 4902 7371 4907
rect 7319 4873 7328 4890
rect 7328 4873 7362 4890
rect 7362 4873 7371 4890
rect 7319 4838 7371 4873
rect 7319 4801 7328 4826
rect 7328 4801 7362 4826
rect 7362 4801 7371 4826
rect 7319 4774 7371 4801
rect 7319 4729 7328 4762
rect 7328 4729 7362 4762
rect 7362 4729 7371 4762
rect 7319 4710 7371 4729
rect 7319 4691 7371 4698
rect 7319 4657 7328 4691
rect 7328 4657 7362 4691
rect 7362 4657 7371 4691
rect 7319 4646 7371 4657
rect 7319 4619 7371 4634
rect 7319 4585 7328 4619
rect 7328 4585 7362 4619
rect 7362 4585 7371 4619
rect 7319 4582 7371 4585
rect 7319 4547 7371 4570
rect 7319 4518 7328 4547
rect 7328 4518 7362 4547
rect 7362 4518 7371 4547
rect 7923 6033 7975 6042
rect 7923 5999 7932 6033
rect 7932 5999 7966 6033
rect 7966 5999 7975 6033
rect 7923 5990 7975 5999
rect 7987 6033 8039 6042
rect 7987 5999 8004 6033
rect 8004 5999 8038 6033
rect 8038 5999 8039 6033
rect 7987 5990 8039 5999
rect 8051 6033 8103 6042
rect 8115 6033 8167 6042
rect 8179 6033 8231 6042
rect 8243 6033 8295 6042
rect 8307 6033 8359 6042
rect 8371 6033 8423 6042
rect 8051 5999 8076 6033
rect 8076 5999 8103 6033
rect 8115 5999 8148 6033
rect 8148 5999 8167 6033
rect 8179 5999 8182 6033
rect 8182 5999 8220 6033
rect 8220 5999 8231 6033
rect 8243 5999 8254 6033
rect 8254 5999 8292 6033
rect 8292 5999 8295 6033
rect 8307 5999 8326 6033
rect 8326 5999 8359 6033
rect 8371 5999 8398 6033
rect 8398 5999 8423 6033
rect 8051 5990 8103 5999
rect 8115 5990 8167 5999
rect 8179 5990 8231 5999
rect 8243 5990 8295 5999
rect 8307 5990 8359 5999
rect 8371 5990 8423 5999
rect 8435 6033 8487 6042
rect 8435 5999 8436 6033
rect 8436 5999 8470 6033
rect 8470 5999 8487 6033
rect 8435 5990 8487 5999
rect 7923 5799 7975 5808
rect 7923 5765 7932 5799
rect 7932 5765 7966 5799
rect 7966 5765 7975 5799
rect 7923 5756 7975 5765
rect 7987 5799 8039 5808
rect 7987 5765 8004 5799
rect 8004 5765 8038 5799
rect 8038 5765 8039 5799
rect 7987 5756 8039 5765
rect 8051 5799 8103 5808
rect 8115 5799 8167 5808
rect 8179 5799 8231 5808
rect 8243 5799 8295 5808
rect 8307 5799 8359 5808
rect 8371 5799 8423 5808
rect 8051 5765 8076 5799
rect 8076 5765 8103 5799
rect 8115 5765 8148 5799
rect 8148 5765 8167 5799
rect 8179 5765 8182 5799
rect 8182 5765 8220 5799
rect 8220 5765 8231 5799
rect 8243 5765 8254 5799
rect 8254 5765 8292 5799
rect 8292 5765 8295 5799
rect 8307 5765 8326 5799
rect 8326 5765 8359 5799
rect 8371 5765 8398 5799
rect 8398 5765 8423 5799
rect 8051 5756 8103 5765
rect 8115 5756 8167 5765
rect 8179 5756 8231 5765
rect 8243 5756 8295 5765
rect 8307 5756 8359 5765
rect 8371 5756 8423 5765
rect 8435 5799 8487 5808
rect 8435 5765 8436 5799
rect 8436 5765 8470 5799
rect 8470 5765 8487 5799
rect 8435 5756 8487 5765
rect 8175 5377 8184 5402
rect 8184 5377 8218 5402
rect 8218 5377 8227 5402
rect 8175 5350 8227 5377
rect 8175 5305 8184 5338
rect 8184 5305 8218 5338
rect 8218 5305 8227 5338
rect 8175 5286 8227 5305
rect 8175 5267 8227 5274
rect 8175 5233 8184 5267
rect 8184 5233 8218 5267
rect 8218 5233 8227 5267
rect 8175 5222 8227 5233
rect 8175 5195 8227 5210
rect 8175 5161 8184 5195
rect 8184 5161 8218 5195
rect 8218 5161 8227 5195
rect 8175 5158 8227 5161
rect 8175 5123 8227 5146
rect 8175 5094 8184 5123
rect 8184 5094 8218 5123
rect 8218 5094 8227 5123
rect 8175 5051 8227 5082
rect 8175 5030 8184 5051
rect 8184 5030 8218 5051
rect 8218 5030 8227 5051
rect 8175 5017 8184 5018
rect 8184 5017 8218 5018
rect 8218 5017 8227 5018
rect 8175 4979 8227 5017
rect 8175 4966 8184 4979
rect 8184 4966 8218 4979
rect 8218 4966 8227 4979
rect 8175 4945 8184 4954
rect 8184 4945 8218 4954
rect 8218 4945 8227 4954
rect 8175 4907 8227 4945
rect 8175 4902 8184 4907
rect 8184 4902 8218 4907
rect 8218 4902 8227 4907
rect 8175 4873 8184 4890
rect 8184 4873 8218 4890
rect 8218 4873 8227 4890
rect 8175 4838 8227 4873
rect 8175 4801 8184 4826
rect 8184 4801 8218 4826
rect 8218 4801 8227 4826
rect 8175 4774 8227 4801
rect 8175 4729 8184 4762
rect 8184 4729 8218 4762
rect 8218 4729 8227 4762
rect 8175 4710 8227 4729
rect 8175 4691 8227 4698
rect 8175 4657 8184 4691
rect 8184 4657 8218 4691
rect 8218 4657 8227 4691
rect 8175 4646 8227 4657
rect 8175 4619 8227 4634
rect 8175 4585 8184 4619
rect 8184 4585 8218 4619
rect 8218 4585 8227 4619
rect 8175 4582 8227 4585
rect 8175 4547 8227 4570
rect 8175 4518 8184 4547
rect 8184 4518 8218 4547
rect 8218 4518 8227 4547
rect 8781 6033 8833 6042
rect 8781 5999 8790 6033
rect 8790 5999 8824 6033
rect 8824 5999 8833 6033
rect 8781 5990 8833 5999
rect 8845 6033 8897 6042
rect 8845 5999 8862 6033
rect 8862 5999 8896 6033
rect 8896 5999 8897 6033
rect 8845 5990 8897 5999
rect 8909 6033 8961 6042
rect 8973 6033 9025 6042
rect 9037 6033 9089 6042
rect 9101 6033 9153 6042
rect 9165 6033 9217 6042
rect 9229 6033 9281 6042
rect 8909 5999 8934 6033
rect 8934 5999 8961 6033
rect 8973 5999 9006 6033
rect 9006 5999 9025 6033
rect 9037 5999 9040 6033
rect 9040 5999 9078 6033
rect 9078 5999 9089 6033
rect 9101 5999 9112 6033
rect 9112 5999 9150 6033
rect 9150 5999 9153 6033
rect 9165 5999 9184 6033
rect 9184 5999 9217 6033
rect 9229 5999 9256 6033
rect 9256 5999 9281 6033
rect 8909 5990 8961 5999
rect 8973 5990 9025 5999
rect 9037 5990 9089 5999
rect 9101 5990 9153 5999
rect 9165 5990 9217 5999
rect 9229 5990 9281 5999
rect 9293 6033 9345 6042
rect 9293 5999 9294 6033
rect 9294 5999 9328 6033
rect 9328 5999 9345 6033
rect 9293 5990 9345 5999
rect 8781 5799 8833 5808
rect 8781 5765 8790 5799
rect 8790 5765 8824 5799
rect 8824 5765 8833 5799
rect 8781 5756 8833 5765
rect 8845 5799 8897 5808
rect 8845 5765 8862 5799
rect 8862 5765 8896 5799
rect 8896 5765 8897 5799
rect 8845 5756 8897 5765
rect 8909 5799 8961 5808
rect 8973 5799 9025 5808
rect 9037 5799 9089 5808
rect 9101 5799 9153 5808
rect 9165 5799 9217 5808
rect 9229 5799 9281 5808
rect 8909 5765 8934 5799
rect 8934 5765 8961 5799
rect 8973 5765 9006 5799
rect 9006 5765 9025 5799
rect 9037 5765 9040 5799
rect 9040 5765 9078 5799
rect 9078 5765 9089 5799
rect 9101 5765 9112 5799
rect 9112 5765 9150 5799
rect 9150 5765 9153 5799
rect 9165 5765 9184 5799
rect 9184 5765 9217 5799
rect 9229 5765 9256 5799
rect 9256 5765 9281 5799
rect 8909 5756 8961 5765
rect 8973 5756 9025 5765
rect 9037 5756 9089 5765
rect 9101 5756 9153 5765
rect 9165 5756 9217 5765
rect 9229 5756 9281 5765
rect 9293 5799 9345 5808
rect 9293 5765 9294 5799
rect 9294 5765 9328 5799
rect 9328 5765 9345 5799
rect 9293 5756 9345 5765
rect 9031 5377 9040 5402
rect 9040 5377 9074 5402
rect 9074 5377 9083 5402
rect 9031 5350 9083 5377
rect 9031 5305 9040 5338
rect 9040 5305 9074 5338
rect 9074 5305 9083 5338
rect 9031 5286 9083 5305
rect 9031 5267 9083 5274
rect 9031 5233 9040 5267
rect 9040 5233 9074 5267
rect 9074 5233 9083 5267
rect 9031 5222 9083 5233
rect 9031 5195 9083 5210
rect 9031 5161 9040 5195
rect 9040 5161 9074 5195
rect 9074 5161 9083 5195
rect 9031 5158 9083 5161
rect 9031 5123 9083 5146
rect 9031 5094 9040 5123
rect 9040 5094 9074 5123
rect 9074 5094 9083 5123
rect 9031 5051 9083 5082
rect 9031 5030 9040 5051
rect 9040 5030 9074 5051
rect 9074 5030 9083 5051
rect 9031 5017 9040 5018
rect 9040 5017 9074 5018
rect 9074 5017 9083 5018
rect 9031 4979 9083 5017
rect 9031 4966 9040 4979
rect 9040 4966 9074 4979
rect 9074 4966 9083 4979
rect 9031 4945 9040 4954
rect 9040 4945 9074 4954
rect 9074 4945 9083 4954
rect 9031 4907 9083 4945
rect 9031 4902 9040 4907
rect 9040 4902 9074 4907
rect 9074 4902 9083 4907
rect 9031 4873 9040 4890
rect 9040 4873 9074 4890
rect 9074 4873 9083 4890
rect 9031 4838 9083 4873
rect 9031 4801 9040 4826
rect 9040 4801 9074 4826
rect 9074 4801 9083 4826
rect 9031 4774 9083 4801
rect 9031 4729 9040 4762
rect 9040 4729 9074 4762
rect 9074 4729 9083 4762
rect 9031 4710 9083 4729
rect 9031 4691 9083 4698
rect 9031 4657 9040 4691
rect 9040 4657 9074 4691
rect 9074 4657 9083 4691
rect 9031 4646 9083 4657
rect 9031 4619 9083 4634
rect 9031 4585 9040 4619
rect 9040 4585 9074 4619
rect 9074 4585 9083 4619
rect 9031 4582 9083 4585
rect 9031 4547 9083 4570
rect 9031 4518 9040 4547
rect 9040 4518 9074 4547
rect 9074 4518 9083 4547
rect 9619 6033 9671 6042
rect 9619 5999 9628 6033
rect 9628 5999 9662 6033
rect 9662 5999 9671 6033
rect 9619 5990 9671 5999
rect 9683 6033 9735 6042
rect 9683 5999 9700 6033
rect 9700 5999 9734 6033
rect 9734 5999 9735 6033
rect 9683 5990 9735 5999
rect 9747 6033 9799 6042
rect 9811 6033 9863 6042
rect 9875 6033 9927 6042
rect 9939 6033 9991 6042
rect 10003 6033 10055 6042
rect 10067 6033 10119 6042
rect 9747 5999 9772 6033
rect 9772 5999 9799 6033
rect 9811 5999 9844 6033
rect 9844 5999 9863 6033
rect 9875 5999 9878 6033
rect 9878 5999 9916 6033
rect 9916 5999 9927 6033
rect 9939 5999 9950 6033
rect 9950 5999 9988 6033
rect 9988 5999 9991 6033
rect 10003 5999 10022 6033
rect 10022 5999 10055 6033
rect 10067 5999 10094 6033
rect 10094 5999 10119 6033
rect 9747 5990 9799 5999
rect 9811 5990 9863 5999
rect 9875 5990 9927 5999
rect 9939 5990 9991 5999
rect 10003 5990 10055 5999
rect 10067 5990 10119 5999
rect 10131 6033 10183 6042
rect 10131 5999 10132 6033
rect 10132 5999 10166 6033
rect 10166 5999 10183 6033
rect 10131 5990 10183 5999
rect 9619 5799 9671 5808
rect 9619 5765 9628 5799
rect 9628 5765 9662 5799
rect 9662 5765 9671 5799
rect 9619 5756 9671 5765
rect 9683 5799 9735 5808
rect 9683 5765 9700 5799
rect 9700 5765 9734 5799
rect 9734 5765 9735 5799
rect 9683 5756 9735 5765
rect 9747 5799 9799 5808
rect 9811 5799 9863 5808
rect 9875 5799 9927 5808
rect 9939 5799 9991 5808
rect 10003 5799 10055 5808
rect 10067 5799 10119 5808
rect 9747 5765 9772 5799
rect 9772 5765 9799 5799
rect 9811 5765 9844 5799
rect 9844 5765 9863 5799
rect 9875 5765 9878 5799
rect 9878 5765 9916 5799
rect 9916 5765 9927 5799
rect 9939 5765 9950 5799
rect 9950 5765 9988 5799
rect 9988 5765 9991 5799
rect 10003 5765 10022 5799
rect 10022 5765 10055 5799
rect 10067 5765 10094 5799
rect 10094 5765 10119 5799
rect 9747 5756 9799 5765
rect 9811 5756 9863 5765
rect 9875 5756 9927 5765
rect 9939 5756 9991 5765
rect 10003 5756 10055 5765
rect 10067 5756 10119 5765
rect 10131 5799 10183 5808
rect 10131 5765 10132 5799
rect 10132 5765 10166 5799
rect 10166 5765 10183 5799
rect 10131 5756 10183 5765
rect 9887 5377 9896 5402
rect 9896 5377 9930 5402
rect 9930 5377 9939 5402
rect 9887 5350 9939 5377
rect 9887 5305 9896 5338
rect 9896 5305 9930 5338
rect 9930 5305 9939 5338
rect 9887 5286 9939 5305
rect 9887 5267 9939 5274
rect 9887 5233 9896 5267
rect 9896 5233 9930 5267
rect 9930 5233 9939 5267
rect 9887 5222 9939 5233
rect 9887 5195 9939 5210
rect 9887 5161 9896 5195
rect 9896 5161 9930 5195
rect 9930 5161 9939 5195
rect 9887 5158 9939 5161
rect 9887 5123 9939 5146
rect 9887 5094 9896 5123
rect 9896 5094 9930 5123
rect 9930 5094 9939 5123
rect 9887 5051 9939 5082
rect 9887 5030 9896 5051
rect 9896 5030 9930 5051
rect 9930 5030 9939 5051
rect 9887 5017 9896 5018
rect 9896 5017 9930 5018
rect 9930 5017 9939 5018
rect 9887 4979 9939 5017
rect 9887 4966 9896 4979
rect 9896 4966 9930 4979
rect 9930 4966 9939 4979
rect 9887 4945 9896 4954
rect 9896 4945 9930 4954
rect 9930 4945 9939 4954
rect 9887 4907 9939 4945
rect 9887 4902 9896 4907
rect 9896 4902 9930 4907
rect 9930 4902 9939 4907
rect 9887 4873 9896 4890
rect 9896 4873 9930 4890
rect 9930 4873 9939 4890
rect 9887 4838 9939 4873
rect 9887 4801 9896 4826
rect 9896 4801 9930 4826
rect 9930 4801 9939 4826
rect 9887 4774 9939 4801
rect 9887 4729 9896 4762
rect 9896 4729 9930 4762
rect 9930 4729 9939 4762
rect 9887 4710 9939 4729
rect 9887 4691 9939 4698
rect 9887 4657 9896 4691
rect 9896 4657 9930 4691
rect 9930 4657 9939 4691
rect 9887 4646 9939 4657
rect 9887 4619 9939 4634
rect 9887 4585 9896 4619
rect 9896 4585 9930 4619
rect 9930 4585 9939 4619
rect 9887 4582 9939 4585
rect 9887 4547 9939 4570
rect 9887 4518 9896 4547
rect 9896 4518 9930 4547
rect 9930 4518 9939 4547
rect 10465 5990 10517 6042
rect 10529 6033 10581 6042
rect 10529 5999 10538 6033
rect 10538 5999 10572 6033
rect 10572 5999 10581 6033
rect 10529 5990 10581 5999
rect 10593 6033 10645 6042
rect 10593 5999 10610 6033
rect 10610 5999 10644 6033
rect 10644 5999 10645 6033
rect 10593 5990 10645 5999
rect 10657 6033 10709 6042
rect 10721 6033 10773 6042
rect 10785 6033 10837 6042
rect 10849 6033 10901 6042
rect 10913 6033 10965 6042
rect 10977 6033 11029 6042
rect 10657 5999 10682 6033
rect 10682 5999 10709 6033
rect 10721 5999 10754 6033
rect 10754 5999 10773 6033
rect 10785 5999 10788 6033
rect 10788 5999 10826 6033
rect 10826 5999 10837 6033
rect 10849 5999 10860 6033
rect 10860 5999 10898 6033
rect 10898 5999 10901 6033
rect 10913 5999 10932 6033
rect 10932 5999 10965 6033
rect 10977 5999 11004 6033
rect 11004 5999 11029 6033
rect 10657 5990 10709 5999
rect 10721 5990 10773 5999
rect 10785 5990 10837 5999
rect 10849 5990 10901 5999
rect 10913 5990 10965 5999
rect 10977 5990 11029 5999
rect 11041 6033 11093 6042
rect 11041 5999 11042 6033
rect 11042 5999 11076 6033
rect 11076 5999 11093 6033
rect 11041 5990 11093 5999
rect 11105 6033 11157 6042
rect 11105 5999 11114 6033
rect 11114 5999 11148 6033
rect 11148 5999 11157 6033
rect 11105 5990 11157 5999
rect 11169 6033 11221 6042
rect 11169 5999 11186 6033
rect 11186 5999 11220 6033
rect 11220 5999 11221 6033
rect 11169 5990 11221 5999
rect 11233 6033 11285 6042
rect 11297 6033 11349 6042
rect 11361 6033 11413 6042
rect 11425 6033 11477 6042
rect 11489 6033 11541 6042
rect 11553 6033 11605 6042
rect 11233 5999 11258 6033
rect 11258 5999 11285 6033
rect 11297 5999 11330 6033
rect 11330 5999 11349 6033
rect 11361 5999 11364 6033
rect 11364 5999 11402 6033
rect 11402 5999 11413 6033
rect 11425 5999 11436 6033
rect 11436 5999 11474 6033
rect 11474 5999 11477 6033
rect 11489 5999 11508 6033
rect 11508 5999 11541 6033
rect 11553 5999 11580 6033
rect 11580 5999 11605 6033
rect 11233 5990 11285 5999
rect 11297 5990 11349 5999
rect 11361 5990 11413 5999
rect 11425 5990 11477 5999
rect 11489 5990 11541 5999
rect 11553 5990 11605 5999
rect 11617 6033 11669 6042
rect 11617 5999 11618 6033
rect 11618 5999 11652 6033
rect 11652 5999 11669 6033
rect 11617 5990 11669 5999
rect 11681 6033 11733 6042
rect 11681 5999 11690 6033
rect 11690 5999 11724 6033
rect 11724 5999 11733 6033
rect 11681 5990 11733 5999
rect 11745 6033 11797 6042
rect 11745 5999 11762 6033
rect 11762 5999 11796 6033
rect 11796 5999 11797 6033
rect 11745 5990 11797 5999
rect 11809 6033 11861 6042
rect 11873 6033 11925 6042
rect 11937 6033 11989 6042
rect 12001 6033 12053 6042
rect 12065 6033 12117 6042
rect 12129 6033 12181 6042
rect 11809 5999 11834 6033
rect 11834 5999 11861 6033
rect 11873 5999 11906 6033
rect 11906 5999 11925 6033
rect 11937 5999 11940 6033
rect 11940 5999 11978 6033
rect 11978 5999 11989 6033
rect 12001 5999 12012 6033
rect 12012 5999 12050 6033
rect 12050 5999 12053 6033
rect 12065 5999 12084 6033
rect 12084 5999 12117 6033
rect 12129 5999 12156 6033
rect 12156 5999 12181 6033
rect 11809 5990 11861 5999
rect 11873 5990 11925 5999
rect 11937 5990 11989 5999
rect 12001 5990 12053 5999
rect 12065 5990 12117 5999
rect 12129 5990 12181 5999
rect 12193 6033 12245 6042
rect 12193 5999 12194 6033
rect 12194 5999 12228 6033
rect 12228 5999 12245 6033
rect 12193 5990 12245 5999
rect 12257 6033 12309 6042
rect 12257 5999 12266 6033
rect 12266 5999 12300 6033
rect 12300 5999 12309 6033
rect 12257 5990 12309 5999
rect 12321 6033 12373 6042
rect 12321 5999 12338 6033
rect 12338 5999 12372 6033
rect 12372 5999 12373 6033
rect 12321 5990 12373 5999
rect 12385 6033 12437 6042
rect 12449 6033 12501 6042
rect 12513 6033 12565 6042
rect 12577 6033 12629 6042
rect 12641 6033 12693 6042
rect 12705 6033 12757 6042
rect 12385 5999 12410 6033
rect 12410 5999 12437 6033
rect 12449 5999 12482 6033
rect 12482 5999 12501 6033
rect 12513 5999 12516 6033
rect 12516 5999 12554 6033
rect 12554 5999 12565 6033
rect 12577 5999 12588 6033
rect 12588 5999 12626 6033
rect 12626 5999 12629 6033
rect 12641 5999 12660 6033
rect 12660 5999 12693 6033
rect 12705 5999 12732 6033
rect 12732 5999 12757 6033
rect 12385 5990 12437 5999
rect 12449 5990 12501 5999
rect 12513 5990 12565 5999
rect 12577 5990 12629 5999
rect 12641 5990 12693 5999
rect 12705 5990 12757 5999
rect 12769 6033 12821 6042
rect 12769 5999 12770 6033
rect 12770 5999 12804 6033
rect 12804 5999 12821 6033
rect 12769 5990 12821 5999
rect 12833 6033 12885 6042
rect 12833 5999 12842 6033
rect 12842 5999 12876 6033
rect 12876 5999 12885 6033
rect 12833 5990 12885 5999
rect 12897 6033 12949 6042
rect 12897 5999 12914 6033
rect 12914 5999 12948 6033
rect 12948 5999 12949 6033
rect 12897 5990 12949 5999
rect 12961 6033 13013 6042
rect 13025 6033 13077 6042
rect 13089 6033 13141 6042
rect 12961 5999 12986 6033
rect 12986 5999 13013 6033
rect 13025 5999 13058 6033
rect 13058 5999 13077 6033
rect 13089 5999 13092 6033
rect 13092 5999 13141 6033
rect 12961 5990 13013 5999
rect 13025 5990 13077 5999
rect 13089 5990 13141 5999
rect 13153 6033 13205 6042
rect 13153 5999 13165 6033
rect 13165 5999 13199 6033
rect 13199 5999 13205 6033
rect 13153 5990 13205 5999
rect 13217 6033 13269 6042
rect 13281 6033 13333 6042
rect 13345 6033 13397 6042
rect 13409 6033 13461 6042
rect 13473 6033 13525 6042
rect 13217 5999 13240 6033
rect 13240 5999 13269 6033
rect 13281 5999 13315 6033
rect 13315 5999 13333 6033
rect 13345 5999 13349 6033
rect 13349 5999 13390 6033
rect 13390 5999 13397 6033
rect 13409 5999 13424 6033
rect 13424 5999 13461 6033
rect 13473 5999 13499 6033
rect 13499 5999 13525 6033
rect 13217 5990 13269 5999
rect 13281 5990 13333 5999
rect 13345 5990 13397 5999
rect 13409 5990 13461 5999
rect 13473 5990 13525 5999
rect 13537 6033 13589 6042
rect 13537 5999 13540 6033
rect 13540 5999 13574 6033
rect 13574 5999 13589 6033
rect 13537 5990 13589 5999
rect 13601 6033 13653 6042
rect 13601 5999 13615 6033
rect 13615 5999 13649 6033
rect 13649 5999 13653 6033
rect 13601 5990 13653 5999
rect 13665 6033 13717 6042
rect 13729 6033 13781 6042
rect 13793 6033 13845 6042
rect 13857 6033 13909 6042
rect 13921 6033 13973 6042
rect 13665 5999 13690 6033
rect 13690 5999 13717 6033
rect 13729 5999 13765 6033
rect 13765 5999 13781 6033
rect 13793 5999 13799 6033
rect 13799 5999 13840 6033
rect 13840 5999 13845 6033
rect 13857 5999 13874 6033
rect 13874 5999 13909 6033
rect 13921 5999 13949 6033
rect 13949 5999 13973 6033
rect 13665 5990 13717 5999
rect 13729 5990 13781 5999
rect 13793 5990 13845 5999
rect 13857 5990 13909 5999
rect 13921 5990 13973 5999
rect 13985 6033 14037 6042
rect 13985 5999 13990 6033
rect 13990 5999 14024 6033
rect 14024 5999 14037 6033
rect 13985 5990 14037 5999
rect 14049 6033 14101 6042
rect 14049 5999 14065 6033
rect 14065 5999 14099 6033
rect 14099 5999 14101 6033
rect 14049 5990 14101 5999
rect 14114 6033 14166 6042
rect 14179 6033 14231 6042
rect 14244 6033 14296 6042
rect 14309 6033 14361 6042
rect 14374 6033 14426 6042
rect 14114 5999 14140 6033
rect 14140 5999 14166 6033
rect 14179 5999 14215 6033
rect 14215 5999 14231 6033
rect 14244 5999 14249 6033
rect 14249 5999 14290 6033
rect 14290 5999 14296 6033
rect 14309 5999 14324 6033
rect 14324 5999 14361 6033
rect 14374 5999 14399 6033
rect 14399 5999 14426 6033
rect 14114 5990 14166 5999
rect 14179 5990 14231 5999
rect 14244 5990 14296 5999
rect 14309 5990 14361 5999
rect 14374 5990 14426 5999
rect 14439 6033 14491 6042
rect 14439 5999 14440 6033
rect 14440 5999 14474 6033
rect 14474 5999 14491 6033
rect 14439 5990 14491 5999
rect 14504 6033 14556 6042
rect 14504 5999 14515 6033
rect 14515 5999 14549 6033
rect 14549 5999 14556 6033
rect 14504 5990 14556 5999
rect 10992 5910 11044 5962
rect 11056 5910 11108 5962
rect 11390 5910 11442 5962
rect 11454 5910 11506 5962
rect 10476 5799 10528 5808
rect 10476 5765 10487 5799
rect 10487 5765 10521 5799
rect 10521 5765 10528 5799
rect 10476 5756 10528 5765
rect 10540 5799 10592 5808
rect 10604 5799 10656 5808
rect 10668 5799 10720 5808
rect 10732 5799 10784 5808
rect 10796 5799 10848 5808
rect 10860 5799 10912 5808
rect 10540 5765 10559 5799
rect 10559 5765 10592 5799
rect 10604 5765 10631 5799
rect 10631 5765 10656 5799
rect 10668 5765 10703 5799
rect 10703 5765 10720 5799
rect 10732 5765 10737 5799
rect 10737 5765 10775 5799
rect 10775 5765 10784 5799
rect 10796 5765 10809 5799
rect 10809 5765 10847 5799
rect 10847 5765 10848 5799
rect 10860 5765 10881 5799
rect 10881 5765 10912 5799
rect 10540 5756 10592 5765
rect 10604 5756 10656 5765
rect 10668 5756 10720 5765
rect 10732 5756 10784 5765
rect 10796 5756 10848 5765
rect 10860 5756 10912 5765
rect 10743 5377 10752 5402
rect 10752 5377 10786 5402
rect 10786 5377 10795 5402
rect 10743 5350 10795 5377
rect 10743 5305 10752 5338
rect 10752 5305 10786 5338
rect 10786 5305 10795 5338
rect 10743 5286 10795 5305
rect 10743 5267 10795 5274
rect 10743 5233 10752 5267
rect 10752 5233 10786 5267
rect 10786 5233 10795 5267
rect 10743 5222 10795 5233
rect 10743 5195 10795 5210
rect 10743 5161 10752 5195
rect 10752 5161 10786 5195
rect 10786 5161 10795 5195
rect 10743 5158 10795 5161
rect 10743 5123 10795 5146
rect 10743 5094 10752 5123
rect 10752 5094 10786 5123
rect 10786 5094 10795 5123
rect 10743 5051 10795 5082
rect 10743 5030 10752 5051
rect 10752 5030 10786 5051
rect 10786 5030 10795 5051
rect 10743 5017 10752 5018
rect 10752 5017 10786 5018
rect 10786 5017 10795 5018
rect 10743 4979 10795 5017
rect 10743 4966 10752 4979
rect 10752 4966 10786 4979
rect 10786 4966 10795 4979
rect 10743 4945 10752 4954
rect 10752 4945 10786 4954
rect 10786 4945 10795 4954
rect 10743 4907 10795 4945
rect 10743 4902 10752 4907
rect 10752 4902 10786 4907
rect 10786 4902 10795 4907
rect 10743 4873 10752 4890
rect 10752 4873 10786 4890
rect 10786 4873 10795 4890
rect 10743 4838 10795 4873
rect 10743 4801 10752 4826
rect 10752 4801 10786 4826
rect 10786 4801 10795 4826
rect 10743 4774 10795 4801
rect 10743 4729 10752 4762
rect 10752 4729 10786 4762
rect 10786 4729 10795 4762
rect 10743 4710 10795 4729
rect 10743 4691 10795 4698
rect 10743 4657 10752 4691
rect 10752 4657 10786 4691
rect 10786 4657 10795 4691
rect 10743 4646 10795 4657
rect 10743 4619 10795 4634
rect 10743 4585 10752 4619
rect 10752 4585 10786 4619
rect 10786 4585 10795 4619
rect 10743 4582 10795 4585
rect 10743 4547 10795 4570
rect 10743 4518 10752 4547
rect 10752 4518 10786 4547
rect 10786 4518 10795 4547
rect 10863 5388 10872 5402
rect 10872 5388 10906 5402
rect 10906 5388 10915 5402
rect 10863 5350 10915 5388
rect 10863 5316 10872 5338
rect 10872 5316 10906 5338
rect 10906 5316 10915 5338
rect 10863 5286 10915 5316
rect 10863 5244 10872 5274
rect 10872 5244 10906 5274
rect 10906 5244 10915 5274
rect 10863 5222 10915 5244
rect 10863 5206 10915 5210
rect 10863 5172 10872 5206
rect 10872 5172 10906 5206
rect 10906 5172 10915 5206
rect 10863 5158 10915 5172
rect 10863 5134 10915 5146
rect 10863 5100 10872 5134
rect 10872 5100 10906 5134
rect 10906 5100 10915 5134
rect 10863 5094 10915 5100
rect 10863 5062 10915 5082
rect 10863 5030 10872 5062
rect 10872 5030 10906 5062
rect 10906 5030 10915 5062
rect 10863 4990 10915 5018
rect 10863 4966 10872 4990
rect 10872 4966 10906 4990
rect 10906 4966 10915 4990
rect 10863 4918 10915 4954
rect 10863 4902 10872 4918
rect 10872 4902 10906 4918
rect 10906 4902 10915 4918
rect 10863 4884 10872 4890
rect 10872 4884 10906 4890
rect 10906 4884 10915 4890
rect 10863 4846 10915 4884
rect 10863 4838 10872 4846
rect 10872 4838 10906 4846
rect 10906 4838 10915 4846
rect 10863 4812 10872 4826
rect 10872 4812 10906 4826
rect 10906 4812 10915 4826
rect 10863 4774 10915 4812
rect 10863 4740 10872 4762
rect 10872 4740 10906 4762
rect 10906 4740 10915 4762
rect 10863 4710 10915 4740
rect 10863 4668 10872 4698
rect 10872 4668 10906 4698
rect 10906 4668 10915 4698
rect 10863 4646 10915 4668
rect 10863 4630 10915 4634
rect 10863 4596 10872 4630
rect 10872 4596 10906 4630
rect 10906 4596 10915 4630
rect 10863 4582 10915 4596
rect 10863 4558 10915 4570
rect 10863 4524 10872 4558
rect 10872 4524 10906 4558
rect 10906 4524 10915 4558
rect 10863 4518 10915 4524
rect 491 3612 500 3637
rect 500 3612 534 3637
rect 534 3612 543 3637
rect 491 3585 543 3612
rect 491 3540 500 3573
rect 500 3540 534 3573
rect 534 3540 543 3573
rect 491 3521 543 3540
rect 491 3502 543 3509
rect 491 3468 500 3502
rect 500 3468 534 3502
rect 534 3468 543 3502
rect 491 3457 543 3468
rect 491 3430 543 3445
rect 491 3396 500 3430
rect 500 3396 534 3430
rect 534 3396 543 3430
rect 491 3393 543 3396
rect 491 3358 543 3381
rect 491 3329 500 3358
rect 500 3329 534 3358
rect 534 3329 543 3358
rect 491 3286 543 3317
rect 491 3265 500 3286
rect 500 3265 534 3286
rect 534 3265 543 3286
rect 491 3252 500 3253
rect 500 3252 534 3253
rect 534 3252 543 3253
rect 491 3214 543 3252
rect 491 3201 500 3214
rect 500 3201 534 3214
rect 534 3201 543 3214
rect 491 3180 500 3189
rect 500 3180 534 3189
rect 534 3180 543 3189
rect 491 3142 543 3180
rect 491 3137 500 3142
rect 500 3137 534 3142
rect 534 3137 543 3142
rect 491 3108 500 3125
rect 500 3108 534 3125
rect 534 3108 543 3125
rect 491 3073 543 3108
rect 491 3036 500 3061
rect 500 3036 534 3061
rect 534 3036 543 3061
rect 491 3009 543 3036
rect 491 2964 500 2997
rect 500 2964 534 2997
rect 534 2964 543 2997
rect 491 2945 543 2964
rect 491 2926 543 2933
rect 491 2892 500 2926
rect 500 2892 534 2926
rect 534 2892 543 2926
rect 491 2881 543 2892
rect 491 2854 543 2869
rect 491 2820 500 2854
rect 500 2820 534 2854
rect 534 2820 543 2854
rect 491 2817 543 2820
rect 491 2782 543 2805
rect 491 2753 500 2782
rect 500 2753 534 2782
rect 534 2753 543 2782
rect 351 2676 360 2685
rect 360 2676 394 2685
rect 394 2676 403 2685
rect 351 2638 403 2676
rect 351 2633 360 2638
rect 360 2633 394 2638
rect 394 2633 403 2638
rect 351 2604 360 2621
rect 360 2604 394 2621
rect 394 2604 403 2621
rect 351 2569 403 2604
rect 351 2532 360 2557
rect 360 2532 394 2557
rect 394 2532 403 2557
rect 351 2505 403 2532
rect 351 2460 360 2493
rect 360 2460 394 2493
rect 394 2460 403 2493
rect 351 2441 403 2460
rect 351 2422 403 2429
rect 351 2388 360 2422
rect 360 2388 394 2422
rect 394 2388 403 2422
rect 351 2377 403 2388
rect 351 2350 403 2365
rect 351 2316 360 2350
rect 360 2316 394 2350
rect 394 2316 403 2350
rect 351 2313 403 2316
rect 351 2278 403 2301
rect 351 2249 360 2278
rect 360 2249 394 2278
rect 394 2249 403 2278
rect 381 2180 433 2232
rect 445 2223 497 2232
rect 445 2189 456 2223
rect 456 2189 490 2223
rect 490 2189 497 2223
rect 445 2180 497 2189
rect 509 2223 561 2232
rect 573 2223 625 2232
rect 509 2189 528 2223
rect 528 2189 561 2223
rect 573 2189 600 2223
rect 600 2189 625 2223
rect 509 2180 561 2189
rect 573 2180 625 2189
rect 637 2180 689 2232
rect 354 2102 406 2154
rect 418 2102 470 2154
rect 482 2102 534 2154
rect 546 2102 598 2154
rect 610 2102 662 2154
rect 674 2102 726 2154
rect 354 2060 406 2075
rect 354 2026 360 2060
rect 360 2026 394 2060
rect 394 2026 406 2060
rect 354 2023 406 2026
rect 418 2069 470 2075
rect 482 2069 534 2075
rect 546 2069 598 2075
rect 610 2069 662 2075
rect 674 2069 726 2075
rect 418 2035 449 2069
rect 449 2035 470 2069
rect 482 2035 483 2069
rect 483 2035 521 2069
rect 521 2035 534 2069
rect 546 2035 555 2069
rect 555 2035 593 2069
rect 593 2035 598 2069
rect 610 2035 627 2069
rect 627 2035 662 2069
rect 674 2035 699 2069
rect 699 2035 726 2069
rect 418 2023 470 2035
rect 482 2023 534 2035
rect 546 2023 598 2035
rect 610 2023 662 2035
rect 674 2023 726 2035
rect 473 1924 525 1933
rect 473 1890 478 1924
rect 478 1890 512 1924
rect 512 1890 525 1924
rect 473 1881 525 1890
rect 537 1924 589 1933
rect 537 1890 550 1924
rect 550 1890 584 1924
rect 584 1890 589 1924
rect 537 1881 589 1890
rect 1347 3630 1356 3637
rect 1356 3630 1390 3637
rect 1390 3630 1399 3637
rect 1347 3592 1399 3630
rect 1347 3585 1356 3592
rect 1356 3585 1390 3592
rect 1390 3585 1399 3592
rect 1347 3558 1356 3573
rect 1356 3558 1390 3573
rect 1390 3558 1399 3573
rect 1347 3521 1399 3558
rect 1347 3486 1356 3509
rect 1356 3486 1390 3509
rect 1390 3486 1399 3509
rect 1347 3457 1399 3486
rect 1347 3414 1356 3445
rect 1356 3414 1390 3445
rect 1390 3414 1399 3445
rect 1347 3393 1399 3414
rect 1347 3376 1399 3381
rect 1347 3342 1356 3376
rect 1356 3342 1390 3376
rect 1390 3342 1399 3376
rect 1347 3329 1399 3342
rect 1347 3304 1399 3317
rect 1347 3270 1356 3304
rect 1356 3270 1390 3304
rect 1390 3270 1399 3304
rect 1347 3265 1399 3270
rect 1347 3232 1399 3253
rect 1347 3201 1356 3232
rect 1356 3201 1390 3232
rect 1390 3201 1399 3232
rect 1347 3160 1399 3189
rect 1347 3137 1356 3160
rect 1356 3137 1390 3160
rect 1390 3137 1399 3160
rect 1347 3088 1399 3125
rect 1347 3073 1356 3088
rect 1356 3073 1390 3088
rect 1390 3073 1399 3088
rect 1347 3054 1356 3061
rect 1356 3054 1390 3061
rect 1390 3054 1399 3061
rect 1347 3016 1399 3054
rect 1347 3009 1356 3016
rect 1356 3009 1390 3016
rect 1390 3009 1399 3016
rect 1347 2982 1356 2997
rect 1356 2982 1390 2997
rect 1390 2982 1399 2997
rect 1347 2945 1399 2982
rect 1347 2910 1356 2933
rect 1356 2910 1390 2933
rect 1390 2910 1399 2933
rect 1347 2881 1399 2910
rect 1347 2838 1356 2869
rect 1356 2838 1390 2869
rect 1390 2838 1399 2869
rect 1347 2817 1399 2838
rect 1347 2800 1399 2805
rect 1347 2766 1356 2800
rect 1356 2766 1390 2800
rect 1390 2766 1399 2800
rect 1347 2753 1399 2766
rect 1047 2223 1099 2229
rect 1111 2223 1163 2229
rect 1175 2223 1227 2229
rect 1239 2223 1291 2229
rect 1047 2189 1069 2223
rect 1069 2189 1099 2223
rect 1111 2189 1141 2223
rect 1141 2189 1163 2223
rect 1175 2189 1213 2223
rect 1213 2189 1227 2223
rect 1239 2189 1247 2223
rect 1247 2189 1291 2223
rect 1047 2177 1099 2189
rect 1111 2177 1163 2189
rect 1175 2177 1227 2189
rect 1239 2177 1291 2189
rect 1047 2102 1099 2154
rect 1111 2102 1163 2154
rect 1175 2102 1227 2154
rect 1239 2102 1291 2154
rect 1047 2069 1099 2075
rect 1111 2069 1163 2075
rect 1175 2069 1227 2075
rect 1239 2069 1291 2075
rect 1047 2035 1069 2069
rect 1069 2035 1099 2069
rect 1111 2035 1141 2069
rect 1141 2035 1163 2069
rect 1175 2035 1213 2069
rect 1213 2035 1227 2069
rect 1239 2035 1247 2069
rect 1247 2035 1291 2069
rect 1047 2023 1099 2035
rect 1111 2023 1163 2035
rect 1175 2023 1227 2035
rect 1239 2023 1291 2035
rect 1436 2223 1488 2229
rect 1500 2223 1552 2229
rect 1564 2223 1616 2229
rect 1628 2223 1680 2229
rect 1436 2189 1458 2223
rect 1458 2189 1488 2223
rect 1500 2189 1530 2223
rect 1530 2189 1552 2223
rect 1564 2189 1602 2223
rect 1602 2189 1616 2223
rect 1628 2189 1636 2223
rect 1636 2189 1680 2223
rect 1436 2177 1488 2189
rect 1500 2177 1552 2189
rect 1564 2177 1616 2189
rect 1628 2177 1680 2189
rect 1436 2102 1488 2154
rect 1500 2102 1552 2154
rect 1564 2102 1616 2154
rect 1628 2102 1680 2154
rect 1436 2069 1488 2075
rect 1500 2069 1552 2075
rect 1564 2069 1616 2075
rect 1628 2069 1680 2075
rect 1436 2035 1458 2069
rect 1458 2035 1488 2069
rect 1500 2035 1530 2069
rect 1530 2035 1552 2069
rect 1564 2035 1602 2069
rect 1602 2035 1616 2069
rect 1628 2035 1636 2069
rect 1636 2035 1680 2069
rect 1436 2023 1488 2035
rect 1500 2023 1552 2035
rect 1564 2023 1616 2035
rect 1628 2023 1680 2035
rect 1315 1881 1367 1933
rect 1379 1881 1431 1933
rect 473 1770 525 1779
rect 473 1736 478 1770
rect 478 1736 512 1770
rect 512 1736 525 1770
rect 473 1727 525 1736
rect 537 1770 589 1779
rect 537 1736 550 1770
rect 550 1736 584 1770
rect 584 1736 589 1770
rect 537 1727 589 1736
rect 869 1727 921 1779
rect 933 1727 985 1779
rect 473 1616 525 1625
rect 473 1582 478 1616
rect 478 1582 512 1616
rect 512 1582 525 1616
rect 473 1573 525 1582
rect 537 1616 589 1625
rect 537 1582 550 1616
rect 550 1582 584 1616
rect 584 1582 589 1616
rect 537 1573 589 1582
rect 2203 3630 2212 3637
rect 2212 3630 2246 3637
rect 2246 3630 2255 3637
rect 2203 3592 2255 3630
rect 2203 3585 2212 3592
rect 2212 3585 2246 3592
rect 2246 3585 2255 3592
rect 2203 3558 2212 3573
rect 2212 3558 2246 3573
rect 2246 3558 2255 3573
rect 2203 3521 2255 3558
rect 2203 3486 2212 3509
rect 2212 3486 2246 3509
rect 2246 3486 2255 3509
rect 2203 3457 2255 3486
rect 2203 3414 2212 3445
rect 2212 3414 2246 3445
rect 2246 3414 2255 3445
rect 2203 3393 2255 3414
rect 2203 3376 2255 3381
rect 2203 3342 2212 3376
rect 2212 3342 2246 3376
rect 2246 3342 2255 3376
rect 2203 3329 2255 3342
rect 2203 3304 2255 3317
rect 2203 3270 2212 3304
rect 2212 3270 2246 3304
rect 2246 3270 2255 3304
rect 2203 3265 2255 3270
rect 2203 3232 2255 3253
rect 2203 3201 2212 3232
rect 2212 3201 2246 3232
rect 2246 3201 2255 3232
rect 2203 3160 2255 3189
rect 2203 3137 2212 3160
rect 2212 3137 2246 3160
rect 2246 3137 2255 3160
rect 2203 3088 2255 3125
rect 2203 3073 2212 3088
rect 2212 3073 2246 3088
rect 2246 3073 2255 3088
rect 2203 3054 2212 3061
rect 2212 3054 2246 3061
rect 2246 3054 2255 3061
rect 2203 3016 2255 3054
rect 2203 3009 2212 3016
rect 2212 3009 2246 3016
rect 2246 3009 2255 3016
rect 2203 2982 2212 2997
rect 2212 2982 2246 2997
rect 2246 2982 2255 2997
rect 2203 2945 2255 2982
rect 2203 2910 2212 2933
rect 2212 2910 2246 2933
rect 2246 2910 2255 2933
rect 2203 2881 2255 2910
rect 2203 2838 2212 2869
rect 2212 2838 2246 2869
rect 2246 2838 2255 2869
rect 2203 2817 2255 2838
rect 2203 2800 2255 2805
rect 2203 2766 2212 2800
rect 2212 2766 2246 2800
rect 2246 2766 2255 2800
rect 2203 2753 2255 2766
rect 1890 2223 1942 2229
rect 1954 2223 2006 2229
rect 2018 2223 2070 2229
rect 2082 2223 2134 2229
rect 1890 2189 1912 2223
rect 1912 2189 1942 2223
rect 1954 2189 1984 2223
rect 1984 2189 2006 2223
rect 2018 2189 2056 2223
rect 2056 2189 2070 2223
rect 2082 2189 2090 2223
rect 2090 2189 2134 2223
rect 1890 2177 1942 2189
rect 1954 2177 2006 2189
rect 2018 2177 2070 2189
rect 2082 2177 2134 2189
rect 1890 2102 1942 2154
rect 1954 2102 2006 2154
rect 2018 2102 2070 2154
rect 2082 2102 2134 2154
rect 1890 2069 1942 2075
rect 1954 2069 2006 2075
rect 2018 2069 2070 2075
rect 2082 2069 2134 2075
rect 1890 2035 1912 2069
rect 1912 2035 1942 2069
rect 1954 2035 1984 2069
rect 1984 2035 2006 2069
rect 2018 2035 2056 2069
rect 2056 2035 2070 2069
rect 2082 2035 2090 2069
rect 2090 2035 2134 2069
rect 1890 2023 1942 2035
rect 1954 2023 2006 2035
rect 2018 2023 2070 2035
rect 2082 2023 2134 2035
rect 2295 2223 2347 2229
rect 2359 2223 2411 2229
rect 2423 2223 2475 2229
rect 2487 2223 2539 2229
rect 2295 2189 2317 2223
rect 2317 2189 2347 2223
rect 2359 2189 2389 2223
rect 2389 2189 2411 2223
rect 2423 2189 2461 2223
rect 2461 2189 2475 2223
rect 2487 2189 2495 2223
rect 2495 2189 2539 2223
rect 2295 2177 2347 2189
rect 2359 2177 2411 2189
rect 2423 2177 2475 2189
rect 2487 2177 2539 2189
rect 2295 2102 2347 2154
rect 2359 2102 2411 2154
rect 2423 2102 2475 2154
rect 2487 2102 2539 2154
rect 2295 2069 2347 2075
rect 2359 2069 2411 2075
rect 2423 2069 2475 2075
rect 2487 2069 2539 2075
rect 2295 2035 2317 2069
rect 2317 2035 2347 2069
rect 2359 2035 2389 2069
rect 2389 2035 2411 2069
rect 2423 2035 2461 2069
rect 2461 2035 2475 2069
rect 2487 2035 2495 2069
rect 2495 2035 2539 2069
rect 2295 2023 2347 2035
rect 2359 2023 2411 2035
rect 2423 2023 2475 2035
rect 2487 2023 2539 2035
rect 2171 1573 2223 1625
rect 2235 1573 2287 1625
rect 473 1462 525 1471
rect 473 1428 478 1462
rect 478 1428 512 1462
rect 512 1428 525 1462
rect 473 1419 525 1428
rect 537 1462 589 1471
rect 537 1428 550 1462
rect 550 1428 584 1462
rect 584 1428 589 1462
rect 537 1419 589 1428
rect 1725 1419 1777 1471
rect 1789 1419 1841 1471
rect 473 1308 525 1317
rect 473 1274 478 1308
rect 478 1274 512 1308
rect 512 1274 525 1308
rect 473 1265 525 1274
rect 537 1308 589 1317
rect 537 1274 550 1308
rect 550 1274 584 1308
rect 584 1274 589 1308
rect 537 1265 589 1274
rect 3059 3630 3068 3637
rect 3068 3630 3102 3637
rect 3102 3630 3111 3637
rect 3059 3592 3111 3630
rect 3059 3585 3068 3592
rect 3068 3585 3102 3592
rect 3102 3585 3111 3592
rect 3059 3558 3068 3573
rect 3068 3558 3102 3573
rect 3102 3558 3111 3573
rect 3059 3521 3111 3558
rect 3059 3486 3068 3509
rect 3068 3486 3102 3509
rect 3102 3486 3111 3509
rect 3059 3457 3111 3486
rect 3059 3414 3068 3445
rect 3068 3414 3102 3445
rect 3102 3414 3111 3445
rect 3059 3393 3111 3414
rect 3059 3376 3111 3381
rect 3059 3342 3068 3376
rect 3068 3342 3102 3376
rect 3102 3342 3111 3376
rect 3059 3329 3111 3342
rect 3059 3304 3111 3317
rect 3059 3270 3068 3304
rect 3068 3270 3102 3304
rect 3102 3270 3111 3304
rect 3059 3265 3111 3270
rect 3059 3232 3111 3253
rect 3059 3201 3068 3232
rect 3068 3201 3102 3232
rect 3102 3201 3111 3232
rect 3059 3160 3111 3189
rect 3059 3137 3068 3160
rect 3068 3137 3102 3160
rect 3102 3137 3111 3160
rect 3059 3088 3111 3125
rect 3059 3073 3068 3088
rect 3068 3073 3102 3088
rect 3102 3073 3111 3088
rect 3059 3054 3068 3061
rect 3068 3054 3102 3061
rect 3102 3054 3111 3061
rect 3059 3016 3111 3054
rect 3059 3009 3068 3016
rect 3068 3009 3102 3016
rect 3102 3009 3111 3016
rect 3059 2982 3068 2997
rect 3068 2982 3102 2997
rect 3102 2982 3111 2997
rect 3059 2945 3111 2982
rect 3059 2910 3068 2933
rect 3068 2910 3102 2933
rect 3102 2910 3111 2933
rect 3059 2881 3111 2910
rect 3059 2838 3068 2869
rect 3068 2838 3102 2869
rect 3102 2838 3111 2869
rect 3059 2817 3111 2838
rect 3059 2800 3111 2805
rect 3059 2766 3068 2800
rect 3068 2766 3102 2800
rect 3102 2766 3111 2800
rect 3059 2753 3111 2766
rect 3915 3630 3924 3637
rect 3924 3630 3958 3637
rect 3958 3630 3967 3637
rect 3915 3592 3967 3630
rect 3915 3585 3924 3592
rect 3924 3585 3958 3592
rect 3958 3585 3967 3592
rect 3915 3558 3924 3573
rect 3924 3558 3958 3573
rect 3958 3558 3967 3573
rect 3915 3521 3967 3558
rect 3915 3486 3924 3509
rect 3924 3486 3958 3509
rect 3958 3486 3967 3509
rect 3915 3457 3967 3486
rect 3915 3414 3924 3445
rect 3924 3414 3958 3445
rect 3958 3414 3967 3445
rect 3915 3393 3967 3414
rect 3915 3376 3967 3381
rect 3915 3342 3924 3376
rect 3924 3342 3958 3376
rect 3958 3342 3967 3376
rect 3915 3329 3967 3342
rect 3915 3304 3967 3317
rect 3915 3270 3924 3304
rect 3924 3270 3958 3304
rect 3958 3270 3967 3304
rect 3915 3265 3967 3270
rect 3915 3232 3967 3253
rect 3915 3201 3924 3232
rect 3924 3201 3958 3232
rect 3958 3201 3967 3232
rect 3915 3160 3967 3189
rect 3915 3137 3924 3160
rect 3924 3137 3958 3160
rect 3958 3137 3967 3160
rect 3915 3088 3967 3125
rect 3915 3073 3924 3088
rect 3924 3073 3958 3088
rect 3958 3073 3967 3088
rect 3915 3054 3924 3061
rect 3924 3054 3958 3061
rect 3958 3054 3967 3061
rect 3915 3016 3967 3054
rect 3915 3009 3924 3016
rect 3924 3009 3958 3016
rect 3958 3009 3967 3016
rect 3915 2982 3924 2997
rect 3924 2982 3958 2997
rect 3958 2982 3967 2997
rect 3915 2945 3967 2982
rect 3915 2910 3924 2933
rect 3924 2910 3958 2933
rect 3958 2910 3967 2933
rect 3915 2881 3967 2910
rect 3915 2838 3924 2869
rect 3924 2838 3958 2869
rect 3958 2838 3967 2869
rect 3915 2817 3967 2838
rect 3915 2800 3967 2805
rect 3915 2766 3924 2800
rect 3924 2766 3958 2800
rect 3958 2766 3967 2800
rect 3915 2753 3967 2766
rect 2759 2223 2811 2229
rect 2823 2223 2875 2229
rect 2887 2223 2939 2229
rect 2951 2223 3003 2229
rect 2759 2189 2781 2223
rect 2781 2189 2811 2223
rect 2823 2189 2853 2223
rect 2853 2189 2875 2223
rect 2887 2189 2925 2223
rect 2925 2189 2939 2223
rect 2951 2189 2959 2223
rect 2959 2189 3003 2223
rect 2759 2177 2811 2189
rect 2823 2177 2875 2189
rect 2887 2177 2939 2189
rect 2951 2177 3003 2189
rect 2759 2102 2811 2154
rect 2823 2102 2875 2154
rect 2887 2102 2939 2154
rect 2951 2102 3003 2154
rect 2759 2069 2811 2075
rect 2823 2069 2875 2075
rect 2887 2069 2939 2075
rect 2951 2069 3003 2075
rect 2759 2035 2781 2069
rect 2781 2035 2811 2069
rect 2823 2035 2853 2069
rect 2853 2035 2875 2069
rect 2887 2035 2925 2069
rect 2925 2035 2939 2069
rect 2951 2035 2959 2069
rect 2959 2035 3003 2069
rect 2759 2023 2811 2035
rect 2823 2023 2875 2035
rect 2887 2023 2939 2035
rect 2951 2023 3003 2035
rect 3209 2223 3261 2232
rect 3209 2189 3219 2223
rect 3219 2189 3253 2223
rect 3253 2189 3261 2223
rect 3209 2180 3261 2189
rect 3273 2223 3325 2232
rect 3273 2189 3291 2223
rect 3291 2189 3325 2223
rect 3273 2180 3325 2189
rect 3337 2223 3389 2232
rect 3401 2223 3453 2232
rect 3465 2223 3517 2232
rect 3529 2223 3581 2232
rect 3593 2223 3645 2232
rect 3337 2189 3363 2223
rect 3363 2189 3389 2223
rect 3401 2189 3435 2223
rect 3435 2189 3453 2223
rect 3465 2189 3469 2223
rect 3469 2189 3507 2223
rect 3507 2189 3517 2223
rect 3529 2189 3541 2223
rect 3541 2189 3579 2223
rect 3579 2189 3581 2223
rect 3593 2189 3613 2223
rect 3613 2189 3645 2223
rect 3337 2180 3389 2189
rect 3401 2180 3453 2189
rect 3465 2180 3517 2189
rect 3529 2180 3581 2189
rect 3593 2180 3645 2189
rect 3209 2102 3261 2154
rect 3273 2102 3325 2154
rect 3337 2102 3389 2154
rect 3401 2102 3453 2154
rect 3465 2102 3517 2154
rect 3529 2102 3581 2154
rect 3593 2102 3645 2154
rect 3209 2069 3261 2078
rect 3209 2035 3219 2069
rect 3219 2035 3253 2069
rect 3253 2035 3261 2069
rect 3209 2026 3261 2035
rect 3273 2069 3325 2078
rect 3273 2035 3291 2069
rect 3291 2035 3325 2069
rect 3273 2026 3325 2035
rect 3337 2069 3389 2078
rect 3401 2069 3453 2078
rect 3465 2069 3517 2078
rect 3529 2069 3581 2078
rect 3593 2069 3645 2078
rect 3337 2035 3363 2069
rect 3363 2035 3389 2069
rect 3401 2035 3435 2069
rect 3435 2035 3453 2069
rect 3465 2035 3469 2069
rect 3469 2035 3507 2069
rect 3507 2035 3517 2069
rect 3529 2035 3541 2069
rect 3541 2035 3579 2069
rect 3579 2035 3581 2069
rect 3593 2035 3613 2069
rect 3613 2035 3645 2069
rect 3337 2026 3389 2035
rect 3401 2026 3453 2035
rect 3465 2026 3517 2035
rect 3529 2026 3581 2035
rect 3593 2026 3645 2035
rect 3213 1881 3265 1933
rect 3277 1881 3329 1933
rect 3209 1727 3261 1779
rect 3273 1727 3325 1779
rect 3213 1573 3265 1625
rect 3277 1573 3329 1625
rect 3209 1419 3261 1471
rect 3273 1419 3325 1471
rect 3213 1265 3265 1317
rect 3277 1265 3329 1317
rect 473 1154 525 1163
rect 473 1120 478 1154
rect 478 1120 512 1154
rect 512 1120 525 1154
rect 473 1111 525 1120
rect 537 1154 589 1163
rect 537 1120 550 1154
rect 550 1120 584 1154
rect 584 1120 589 1154
rect 537 1111 589 1120
rect 2581 1111 2633 1163
rect 2645 1111 2697 1163
rect 3209 1111 3261 1163
rect 3273 1111 3325 1163
rect 473 1000 525 1009
rect 473 966 478 1000
rect 478 966 512 1000
rect 512 966 525 1000
rect 473 957 525 966
rect 537 1000 589 1009
rect 537 966 550 1000
rect 550 966 584 1000
rect 584 966 589 1000
rect 537 957 589 966
rect 3213 957 3265 1009
rect 3277 957 3329 1009
rect 3971 2223 4023 2229
rect 4035 2223 4087 2229
rect 4099 2223 4151 2229
rect 4163 2223 4215 2229
rect 3971 2189 3993 2223
rect 3993 2189 4023 2223
rect 4035 2189 4065 2223
rect 4065 2189 4087 2223
rect 4099 2189 4137 2223
rect 4137 2189 4151 2223
rect 4163 2189 4171 2223
rect 4171 2189 4215 2223
rect 3971 2177 4023 2189
rect 4035 2177 4087 2189
rect 4099 2177 4151 2189
rect 4163 2177 4215 2189
rect 3971 2102 4023 2154
rect 4035 2102 4087 2154
rect 4099 2102 4151 2154
rect 4163 2102 4215 2154
rect 3971 2069 4023 2075
rect 4035 2069 4087 2075
rect 4099 2069 4151 2075
rect 4163 2069 4215 2075
rect 3971 2035 3993 2069
rect 3993 2035 4023 2069
rect 4035 2035 4065 2069
rect 4065 2035 4087 2069
rect 4099 2035 4137 2069
rect 4137 2035 4151 2069
rect 4163 2035 4171 2069
rect 4171 2035 4215 2069
rect 3971 2023 4023 2035
rect 4035 2023 4087 2035
rect 4099 2023 4151 2035
rect 4163 2023 4215 2035
rect 473 846 525 855
rect 473 812 478 846
rect 478 812 512 846
rect 512 812 525 846
rect 473 803 525 812
rect 537 846 589 855
rect 537 812 550 846
rect 550 812 584 846
rect 584 812 589 846
rect 537 803 589 812
rect 3209 803 3261 855
rect 3273 803 3325 855
rect 3762 803 3814 855
rect 3826 803 3878 855
rect 473 692 525 701
rect 473 658 478 692
rect 478 658 512 692
rect 512 658 525 692
rect 473 649 525 658
rect 537 692 589 701
rect 537 658 550 692
rect 550 658 584 692
rect 584 658 589 692
rect 537 649 589 658
rect 3213 649 3265 701
rect 3277 649 3329 701
rect 4771 3630 4780 3637
rect 4780 3630 4814 3637
rect 4814 3630 4823 3637
rect 4771 3592 4823 3630
rect 4771 3585 4780 3592
rect 4780 3585 4814 3592
rect 4814 3585 4823 3592
rect 4771 3558 4780 3573
rect 4780 3558 4814 3573
rect 4814 3558 4823 3573
rect 4771 3521 4823 3558
rect 4771 3486 4780 3509
rect 4780 3486 4814 3509
rect 4814 3486 4823 3509
rect 4771 3457 4823 3486
rect 4771 3414 4780 3445
rect 4780 3414 4814 3445
rect 4814 3414 4823 3445
rect 4771 3393 4823 3414
rect 4771 3376 4823 3381
rect 4771 3342 4780 3376
rect 4780 3342 4814 3376
rect 4814 3342 4823 3376
rect 4771 3329 4823 3342
rect 4771 3304 4823 3317
rect 4771 3270 4780 3304
rect 4780 3270 4814 3304
rect 4814 3270 4823 3304
rect 4771 3265 4823 3270
rect 4771 3232 4823 3253
rect 4771 3201 4780 3232
rect 4780 3201 4814 3232
rect 4814 3201 4823 3232
rect 4771 3160 4823 3189
rect 4771 3137 4780 3160
rect 4780 3137 4814 3160
rect 4814 3137 4823 3160
rect 4771 3088 4823 3125
rect 4771 3073 4780 3088
rect 4780 3073 4814 3088
rect 4814 3073 4823 3088
rect 4771 3054 4780 3061
rect 4780 3054 4814 3061
rect 4814 3054 4823 3061
rect 4771 3016 4823 3054
rect 4771 3009 4780 3016
rect 4780 3009 4814 3016
rect 4814 3009 4823 3016
rect 4771 2982 4780 2997
rect 4780 2982 4814 2997
rect 4814 2982 4823 2997
rect 4771 2945 4823 2982
rect 4771 2910 4780 2933
rect 4780 2910 4814 2933
rect 4814 2910 4823 2933
rect 4771 2881 4823 2910
rect 4771 2838 4780 2869
rect 4780 2838 4814 2869
rect 4814 2838 4823 2869
rect 4771 2817 4823 2838
rect 4771 2800 4823 2805
rect 4771 2766 4780 2800
rect 4780 2766 4814 2800
rect 4814 2766 4823 2800
rect 4771 2753 4823 2766
rect 4466 2223 4518 2229
rect 4530 2223 4582 2229
rect 4594 2223 4646 2229
rect 4658 2223 4710 2229
rect 4466 2189 4488 2223
rect 4488 2189 4518 2223
rect 4530 2189 4560 2223
rect 4560 2189 4582 2223
rect 4594 2189 4632 2223
rect 4632 2189 4646 2223
rect 4658 2189 4666 2223
rect 4666 2189 4710 2223
rect 4466 2177 4518 2189
rect 4530 2177 4582 2189
rect 4594 2177 4646 2189
rect 4658 2177 4710 2189
rect 4466 2102 4518 2154
rect 4530 2102 4582 2154
rect 4594 2102 4646 2154
rect 4658 2102 4710 2154
rect 4466 2069 4518 2075
rect 4530 2069 4582 2075
rect 4594 2069 4646 2075
rect 4658 2069 4710 2075
rect 4466 2035 4488 2069
rect 4488 2035 4518 2069
rect 4530 2035 4560 2069
rect 4560 2035 4582 2069
rect 4594 2035 4632 2069
rect 4632 2035 4646 2069
rect 4658 2035 4666 2069
rect 4666 2035 4710 2069
rect 4466 2023 4518 2035
rect 4530 2023 4582 2035
rect 4594 2023 4646 2035
rect 4658 2023 4710 2035
rect 4860 2223 4912 2229
rect 4924 2223 4976 2229
rect 4988 2223 5040 2229
rect 5052 2223 5104 2229
rect 4860 2189 4882 2223
rect 4882 2189 4912 2223
rect 4924 2189 4954 2223
rect 4954 2189 4976 2223
rect 4988 2189 5026 2223
rect 5026 2189 5040 2223
rect 5052 2189 5060 2223
rect 5060 2189 5104 2223
rect 4860 2177 4912 2189
rect 4924 2177 4976 2189
rect 4988 2177 5040 2189
rect 5052 2177 5104 2189
rect 4860 2102 4912 2154
rect 4924 2102 4976 2154
rect 4988 2102 5040 2154
rect 5052 2102 5104 2154
rect 4860 2069 4912 2075
rect 4924 2069 4976 2075
rect 4988 2069 5040 2075
rect 5052 2069 5104 2075
rect 4860 2035 4882 2069
rect 4882 2035 4912 2069
rect 4924 2035 4954 2069
rect 4954 2035 4976 2069
rect 4988 2035 5026 2069
rect 5026 2035 5040 2069
rect 5052 2035 5060 2069
rect 5060 2035 5104 2069
rect 4860 2023 4912 2035
rect 4924 2023 4976 2035
rect 4988 2023 5040 2035
rect 5052 2023 5104 2035
rect 4739 957 4791 1009
rect 4803 957 4855 1009
rect 473 538 525 547
rect 473 504 478 538
rect 478 504 512 538
rect 512 504 525 538
rect 473 495 525 504
rect 537 538 589 547
rect 537 504 550 538
rect 550 504 584 538
rect 584 504 589 538
rect 537 495 589 504
rect 3209 495 3261 547
rect 3273 495 3325 547
rect 4293 495 4345 547
rect 4357 495 4409 547
rect 473 384 525 393
rect 473 350 478 384
rect 478 350 512 384
rect 512 350 525 384
rect 473 341 525 350
rect 537 384 589 393
rect 537 350 550 384
rect 550 350 584 384
rect 584 350 589 384
rect 537 341 589 350
rect 3213 341 3265 393
rect 3277 341 3329 393
rect 5627 3630 5636 3637
rect 5636 3630 5670 3637
rect 5670 3630 5679 3637
rect 5627 3592 5679 3630
rect 5627 3585 5636 3592
rect 5636 3585 5670 3592
rect 5670 3585 5679 3592
rect 5627 3558 5636 3573
rect 5636 3558 5670 3573
rect 5670 3558 5679 3573
rect 5627 3521 5679 3558
rect 5627 3486 5636 3509
rect 5636 3486 5670 3509
rect 5670 3486 5679 3509
rect 5627 3457 5679 3486
rect 5627 3414 5636 3445
rect 5636 3414 5670 3445
rect 5670 3414 5679 3445
rect 5627 3393 5679 3414
rect 5627 3376 5679 3381
rect 5627 3342 5636 3376
rect 5636 3342 5670 3376
rect 5670 3342 5679 3376
rect 5627 3329 5679 3342
rect 5627 3304 5679 3317
rect 5627 3270 5636 3304
rect 5636 3270 5670 3304
rect 5670 3270 5679 3304
rect 5627 3265 5679 3270
rect 5627 3232 5679 3253
rect 5627 3201 5636 3232
rect 5636 3201 5670 3232
rect 5670 3201 5679 3232
rect 5627 3160 5679 3189
rect 5627 3137 5636 3160
rect 5636 3137 5670 3160
rect 5670 3137 5679 3160
rect 5627 3088 5679 3125
rect 5627 3073 5636 3088
rect 5636 3073 5670 3088
rect 5670 3073 5679 3088
rect 5627 3054 5636 3061
rect 5636 3054 5670 3061
rect 5670 3054 5679 3061
rect 5627 3016 5679 3054
rect 5627 3009 5636 3016
rect 5636 3009 5670 3016
rect 5670 3009 5679 3016
rect 5627 2982 5636 2997
rect 5636 2982 5670 2997
rect 5670 2982 5679 2997
rect 5627 2945 5679 2982
rect 5627 2910 5636 2933
rect 5636 2910 5670 2933
rect 5670 2910 5679 2933
rect 5627 2881 5679 2910
rect 5627 2838 5636 2869
rect 5636 2838 5670 2869
rect 5670 2838 5679 2869
rect 5627 2817 5679 2838
rect 5627 2800 5679 2805
rect 5627 2766 5636 2800
rect 5636 2766 5670 2800
rect 5670 2766 5679 2800
rect 5627 2753 5679 2766
rect 5325 2223 5377 2229
rect 5389 2223 5441 2229
rect 5453 2223 5505 2229
rect 5517 2223 5569 2229
rect 5325 2189 5347 2223
rect 5347 2189 5377 2223
rect 5389 2189 5419 2223
rect 5419 2189 5441 2223
rect 5453 2189 5491 2223
rect 5491 2189 5505 2223
rect 5517 2189 5525 2223
rect 5525 2189 5569 2223
rect 5325 2177 5377 2189
rect 5389 2177 5441 2189
rect 5453 2177 5505 2189
rect 5517 2177 5569 2189
rect 5325 2102 5377 2154
rect 5389 2102 5441 2154
rect 5453 2102 5505 2154
rect 5517 2102 5569 2154
rect 5325 2069 5377 2075
rect 5389 2069 5441 2075
rect 5453 2069 5505 2075
rect 5517 2069 5569 2075
rect 5325 2035 5347 2069
rect 5347 2035 5377 2069
rect 5389 2035 5419 2069
rect 5419 2035 5441 2069
rect 5453 2035 5491 2069
rect 5491 2035 5505 2069
rect 5517 2035 5525 2069
rect 5525 2035 5569 2069
rect 5325 2023 5377 2035
rect 5389 2023 5441 2035
rect 5453 2023 5505 2035
rect 5517 2023 5569 2035
rect 5719 2223 5771 2229
rect 5783 2223 5835 2229
rect 5847 2223 5899 2229
rect 5911 2223 5963 2229
rect 5719 2189 5741 2223
rect 5741 2189 5771 2223
rect 5783 2189 5813 2223
rect 5813 2189 5835 2223
rect 5847 2189 5885 2223
rect 5885 2189 5899 2223
rect 5911 2189 5919 2223
rect 5919 2189 5963 2223
rect 5719 2177 5771 2189
rect 5783 2177 5835 2189
rect 5847 2177 5899 2189
rect 5911 2177 5963 2189
rect 5719 2102 5771 2154
rect 5783 2102 5835 2154
rect 5847 2102 5899 2154
rect 5911 2102 5963 2154
rect 5719 2069 5771 2075
rect 5783 2069 5835 2075
rect 5847 2069 5899 2075
rect 5911 2069 5963 2075
rect 5719 2035 5741 2069
rect 5741 2035 5771 2069
rect 5783 2035 5813 2069
rect 5813 2035 5835 2069
rect 5847 2035 5885 2069
rect 5885 2035 5899 2069
rect 5911 2035 5919 2069
rect 5919 2035 5963 2069
rect 5719 2023 5771 2035
rect 5783 2023 5835 2035
rect 5847 2023 5899 2035
rect 5911 2023 5963 2035
rect 6483 3630 6492 3637
rect 6492 3630 6526 3637
rect 6526 3630 6535 3637
rect 6483 3592 6535 3630
rect 6483 3585 6492 3592
rect 6492 3585 6526 3592
rect 6526 3585 6535 3592
rect 6483 3558 6492 3573
rect 6492 3558 6526 3573
rect 6526 3558 6535 3573
rect 6483 3521 6535 3558
rect 6483 3486 6492 3509
rect 6492 3486 6526 3509
rect 6526 3486 6535 3509
rect 6483 3457 6535 3486
rect 6483 3414 6492 3445
rect 6492 3414 6526 3445
rect 6526 3414 6535 3445
rect 6483 3393 6535 3414
rect 6483 3376 6535 3381
rect 6483 3342 6492 3376
rect 6492 3342 6526 3376
rect 6526 3342 6535 3376
rect 6483 3329 6535 3342
rect 6483 3304 6535 3317
rect 6483 3270 6492 3304
rect 6492 3270 6526 3304
rect 6526 3270 6535 3304
rect 6483 3265 6535 3270
rect 6483 3232 6535 3253
rect 6483 3201 6492 3232
rect 6492 3201 6526 3232
rect 6526 3201 6535 3232
rect 6483 3160 6535 3189
rect 6483 3137 6492 3160
rect 6492 3137 6526 3160
rect 6526 3137 6535 3160
rect 6483 3088 6535 3125
rect 6483 3073 6492 3088
rect 6492 3073 6526 3088
rect 6526 3073 6535 3088
rect 6483 3054 6492 3061
rect 6492 3054 6526 3061
rect 6526 3054 6535 3061
rect 6483 3016 6535 3054
rect 6483 3009 6492 3016
rect 6492 3009 6526 3016
rect 6526 3009 6535 3016
rect 6483 2982 6492 2997
rect 6492 2982 6526 2997
rect 6526 2982 6535 2997
rect 6483 2945 6535 2982
rect 6483 2910 6492 2933
rect 6492 2910 6526 2933
rect 6526 2910 6535 2933
rect 6483 2881 6535 2910
rect 6483 2838 6492 2869
rect 6492 2838 6526 2869
rect 6526 2838 6535 2869
rect 6483 2817 6535 2838
rect 6483 2800 6535 2805
rect 6483 2766 6492 2800
rect 6492 2766 6526 2800
rect 6526 2766 6535 2800
rect 6483 2753 6535 2766
rect 6189 2223 6241 2229
rect 6253 2223 6305 2229
rect 6317 2223 6369 2229
rect 6381 2223 6433 2229
rect 6189 2189 6211 2223
rect 6211 2189 6241 2223
rect 6253 2189 6283 2223
rect 6283 2189 6305 2223
rect 6317 2189 6355 2223
rect 6355 2189 6369 2223
rect 6381 2189 6389 2223
rect 6389 2189 6433 2223
rect 6189 2177 6241 2189
rect 6253 2177 6305 2189
rect 6317 2177 6369 2189
rect 6381 2177 6433 2189
rect 6189 2102 6241 2154
rect 6253 2102 6305 2154
rect 6317 2102 6369 2154
rect 6381 2102 6433 2154
rect 6189 2069 6241 2075
rect 6253 2069 6305 2075
rect 6317 2069 6369 2075
rect 6381 2069 6433 2075
rect 6189 2035 6211 2069
rect 6211 2035 6241 2069
rect 6253 2035 6283 2069
rect 6283 2035 6305 2069
rect 6317 2035 6355 2069
rect 6355 2035 6369 2069
rect 6381 2035 6389 2069
rect 6389 2035 6433 2069
rect 6189 2023 6241 2035
rect 6253 2023 6305 2035
rect 6317 2023 6369 2035
rect 6381 2023 6433 2035
rect 5807 1881 5859 1933
rect 5871 1881 5923 1933
rect 5595 649 5647 701
rect 5659 649 5711 701
rect 7339 3630 7348 3637
rect 7348 3630 7382 3637
rect 7382 3630 7391 3637
rect 7339 3592 7391 3630
rect 7339 3585 7348 3592
rect 7348 3585 7382 3592
rect 7382 3585 7391 3592
rect 7339 3558 7348 3573
rect 7348 3558 7382 3573
rect 7382 3558 7391 3573
rect 7339 3521 7391 3558
rect 7339 3486 7348 3509
rect 7348 3486 7382 3509
rect 7382 3486 7391 3509
rect 7339 3457 7391 3486
rect 7339 3414 7348 3445
rect 7348 3414 7382 3445
rect 7382 3414 7391 3445
rect 7339 3393 7391 3414
rect 7339 3376 7391 3381
rect 7339 3342 7348 3376
rect 7348 3342 7382 3376
rect 7382 3342 7391 3376
rect 7339 3329 7391 3342
rect 7339 3304 7391 3317
rect 7339 3270 7348 3304
rect 7348 3270 7382 3304
rect 7382 3270 7391 3304
rect 7339 3265 7391 3270
rect 7339 3232 7391 3253
rect 7339 3201 7348 3232
rect 7348 3201 7382 3232
rect 7382 3201 7391 3232
rect 7339 3160 7391 3189
rect 7339 3137 7348 3160
rect 7348 3137 7382 3160
rect 7382 3137 7391 3160
rect 7339 3088 7391 3125
rect 7339 3073 7348 3088
rect 7348 3073 7382 3088
rect 7382 3073 7391 3088
rect 7339 3054 7348 3061
rect 7348 3054 7382 3061
rect 7382 3054 7391 3061
rect 7339 3016 7391 3054
rect 7339 3009 7348 3016
rect 7348 3009 7382 3016
rect 7382 3009 7391 3016
rect 7339 2982 7348 2997
rect 7348 2982 7382 2997
rect 7382 2982 7391 2997
rect 7339 2945 7391 2982
rect 7339 2910 7348 2933
rect 7348 2910 7382 2933
rect 7382 2910 7391 2933
rect 7339 2881 7391 2910
rect 7339 2838 7348 2869
rect 7348 2838 7382 2869
rect 7382 2838 7391 2869
rect 7339 2817 7391 2838
rect 7339 2800 7391 2805
rect 7339 2766 7348 2800
rect 7348 2766 7382 2800
rect 7382 2766 7391 2800
rect 7339 2753 7391 2766
rect 8195 3630 8204 3637
rect 8204 3630 8238 3637
rect 8238 3630 8247 3637
rect 8195 3592 8247 3630
rect 8195 3585 8204 3592
rect 8204 3585 8238 3592
rect 8238 3585 8247 3592
rect 8195 3558 8204 3573
rect 8204 3558 8238 3573
rect 8238 3558 8247 3573
rect 8195 3521 8247 3558
rect 8195 3486 8204 3509
rect 8204 3486 8238 3509
rect 8238 3486 8247 3509
rect 8195 3457 8247 3486
rect 8195 3414 8204 3445
rect 8204 3414 8238 3445
rect 8238 3414 8247 3445
rect 8195 3393 8247 3414
rect 8195 3376 8247 3381
rect 8195 3342 8204 3376
rect 8204 3342 8238 3376
rect 8238 3342 8247 3376
rect 8195 3329 8247 3342
rect 8195 3304 8247 3317
rect 8195 3270 8204 3304
rect 8204 3270 8238 3304
rect 8238 3270 8247 3304
rect 8195 3265 8247 3270
rect 8195 3232 8247 3253
rect 8195 3201 8204 3232
rect 8204 3201 8238 3232
rect 8238 3201 8247 3232
rect 8195 3160 8247 3189
rect 8195 3137 8204 3160
rect 8204 3137 8238 3160
rect 8238 3137 8247 3160
rect 8195 3088 8247 3125
rect 8195 3073 8204 3088
rect 8204 3073 8238 3088
rect 8238 3073 8247 3088
rect 8195 3054 8204 3061
rect 8204 3054 8238 3061
rect 8238 3054 8247 3061
rect 8195 3016 8247 3054
rect 8195 3009 8204 3016
rect 8204 3009 8238 3016
rect 8238 3009 8247 3016
rect 8195 2982 8204 2997
rect 8204 2982 8238 2997
rect 8238 2982 8247 2997
rect 8195 2945 8247 2982
rect 8195 2910 8204 2933
rect 8204 2910 8238 2933
rect 8238 2910 8247 2933
rect 8195 2881 8247 2910
rect 8195 2838 8204 2869
rect 8204 2838 8238 2869
rect 8238 2838 8247 2869
rect 8195 2817 8247 2838
rect 8195 2800 8247 2805
rect 8195 2766 8204 2800
rect 8204 2766 8238 2800
rect 8238 2766 8247 2800
rect 8195 2753 8247 2766
rect 9051 3630 9060 3637
rect 9060 3630 9094 3637
rect 9094 3630 9103 3637
rect 9051 3592 9103 3630
rect 9051 3585 9060 3592
rect 9060 3585 9094 3592
rect 9094 3585 9103 3592
rect 9051 3558 9060 3573
rect 9060 3558 9094 3573
rect 9094 3558 9103 3573
rect 9051 3521 9103 3558
rect 9051 3486 9060 3509
rect 9060 3486 9094 3509
rect 9094 3486 9103 3509
rect 9051 3457 9103 3486
rect 9051 3414 9060 3445
rect 9060 3414 9094 3445
rect 9094 3414 9103 3445
rect 9051 3393 9103 3414
rect 9051 3376 9103 3381
rect 9051 3342 9060 3376
rect 9060 3342 9094 3376
rect 9094 3342 9103 3376
rect 9051 3329 9103 3342
rect 9051 3304 9103 3317
rect 9051 3270 9060 3304
rect 9060 3270 9094 3304
rect 9094 3270 9103 3304
rect 9051 3265 9103 3270
rect 9051 3232 9103 3253
rect 9051 3201 9060 3232
rect 9060 3201 9094 3232
rect 9094 3201 9103 3232
rect 9051 3160 9103 3189
rect 9051 3137 9060 3160
rect 9060 3137 9094 3160
rect 9094 3137 9103 3160
rect 9051 3088 9103 3125
rect 9051 3073 9060 3088
rect 9060 3073 9094 3088
rect 9094 3073 9103 3088
rect 9051 3054 9060 3061
rect 9060 3054 9094 3061
rect 9094 3054 9103 3061
rect 9051 3016 9103 3054
rect 9051 3009 9060 3016
rect 9060 3009 9094 3016
rect 9094 3009 9103 3016
rect 9051 2982 9060 2997
rect 9060 2982 9094 2997
rect 9094 2982 9103 2997
rect 9051 2945 9103 2982
rect 9051 2910 9060 2933
rect 9060 2910 9094 2933
rect 9094 2910 9103 2933
rect 9051 2881 9103 2910
rect 9051 2838 9060 2869
rect 9060 2838 9094 2869
rect 9094 2838 9103 2869
rect 9051 2817 9103 2838
rect 9051 2800 9103 2805
rect 9051 2766 9060 2800
rect 9060 2766 9094 2800
rect 9094 2766 9103 2800
rect 9051 2753 9103 2766
rect 9907 3630 9916 3637
rect 9916 3630 9950 3637
rect 9950 3630 9959 3637
rect 9907 3592 9959 3630
rect 9907 3585 9916 3592
rect 9916 3585 9950 3592
rect 9950 3585 9959 3592
rect 9907 3558 9916 3573
rect 9916 3558 9950 3573
rect 9950 3558 9959 3573
rect 9907 3521 9959 3558
rect 9907 3486 9916 3509
rect 9916 3486 9950 3509
rect 9950 3486 9959 3509
rect 9907 3457 9959 3486
rect 9907 3414 9916 3445
rect 9916 3414 9950 3445
rect 9950 3414 9959 3445
rect 9907 3393 9959 3414
rect 9907 3376 9959 3381
rect 9907 3342 9916 3376
rect 9916 3342 9950 3376
rect 9950 3342 9959 3376
rect 9907 3329 9959 3342
rect 9907 3304 9959 3317
rect 9907 3270 9916 3304
rect 9916 3270 9950 3304
rect 9950 3270 9959 3304
rect 9907 3265 9959 3270
rect 9907 3232 9959 3253
rect 9907 3201 9916 3232
rect 9916 3201 9950 3232
rect 9950 3201 9959 3232
rect 9907 3160 9959 3189
rect 9907 3137 9916 3160
rect 9916 3137 9950 3160
rect 9950 3137 9959 3160
rect 9907 3088 9959 3125
rect 9907 3073 9916 3088
rect 9916 3073 9950 3088
rect 9950 3073 9959 3088
rect 9907 3054 9916 3061
rect 9916 3054 9950 3061
rect 9950 3054 9959 3061
rect 9907 3016 9959 3054
rect 9907 3009 9916 3016
rect 9916 3009 9950 3016
rect 9950 3009 9959 3016
rect 9907 2982 9916 2997
rect 9916 2982 9950 2997
rect 9950 2982 9959 2997
rect 9907 2945 9959 2982
rect 9907 2910 9916 2933
rect 9916 2910 9950 2933
rect 9950 2910 9959 2933
rect 9907 2881 9959 2910
rect 9907 2838 9916 2869
rect 9916 2838 9950 2869
rect 9950 2838 9959 2869
rect 9907 2817 9959 2838
rect 9907 2800 9959 2805
rect 9907 2766 9916 2800
rect 9916 2766 9950 2800
rect 9950 2766 9959 2800
rect 9907 2753 9959 2766
rect 10763 3630 10772 3637
rect 10772 3630 10806 3637
rect 10806 3630 10815 3637
rect 10763 3592 10815 3630
rect 10763 3585 10772 3592
rect 10772 3585 10806 3592
rect 10806 3585 10815 3592
rect 10763 3558 10772 3573
rect 10772 3558 10806 3573
rect 10806 3558 10815 3573
rect 10763 3521 10815 3558
rect 10763 3486 10772 3509
rect 10772 3486 10806 3509
rect 10806 3486 10815 3509
rect 10763 3457 10815 3486
rect 10763 3414 10772 3445
rect 10772 3414 10806 3445
rect 10806 3414 10815 3445
rect 10763 3393 10815 3414
rect 10763 3376 10815 3381
rect 10763 3342 10772 3376
rect 10772 3342 10806 3376
rect 10806 3342 10815 3376
rect 10763 3329 10815 3342
rect 10763 3304 10815 3317
rect 10763 3270 10772 3304
rect 10772 3270 10806 3304
rect 10806 3270 10815 3304
rect 10763 3265 10815 3270
rect 10763 3232 10815 3253
rect 10763 3201 10772 3232
rect 10772 3201 10806 3232
rect 10806 3201 10815 3232
rect 10763 3160 10815 3189
rect 10763 3137 10772 3160
rect 10772 3137 10806 3160
rect 10806 3137 10815 3160
rect 10763 3088 10815 3125
rect 10763 3073 10772 3088
rect 10772 3073 10806 3088
rect 10806 3073 10815 3088
rect 10763 3054 10772 3061
rect 10772 3054 10806 3061
rect 10806 3054 10815 3061
rect 10763 3016 10815 3054
rect 10763 3009 10772 3016
rect 10772 3009 10806 3016
rect 10806 3009 10815 3016
rect 10763 2982 10772 2997
rect 10772 2982 10806 2997
rect 10806 2982 10815 2997
rect 10763 2945 10815 2982
rect 10763 2910 10772 2933
rect 10772 2910 10806 2933
rect 10806 2910 10815 2933
rect 10763 2881 10815 2910
rect 10763 2838 10772 2869
rect 10772 2838 10806 2869
rect 10806 2838 10815 2869
rect 10763 2817 10815 2838
rect 10763 2800 10815 2805
rect 10763 2766 10772 2800
rect 10772 2766 10806 2800
rect 10806 2766 10815 2800
rect 10763 2753 10815 2766
rect 10904 2676 10912 2679
rect 10912 2676 10946 2679
rect 10946 2676 10956 2679
rect 10904 2638 10956 2676
rect 10904 2627 10912 2638
rect 10912 2627 10946 2638
rect 10946 2627 10956 2638
rect 10904 2604 10912 2615
rect 10912 2604 10946 2615
rect 10946 2604 10956 2615
rect 10904 2566 10956 2604
rect 10904 2563 10912 2566
rect 10912 2563 10946 2566
rect 10946 2563 10956 2566
rect 10904 2532 10912 2550
rect 10912 2532 10946 2550
rect 10946 2532 10956 2550
rect 10904 2498 10956 2532
rect 10904 2460 10912 2485
rect 10912 2460 10946 2485
rect 10946 2460 10956 2485
rect 10904 2433 10956 2460
rect 10904 2388 10912 2420
rect 10912 2388 10946 2420
rect 10946 2388 10956 2420
rect 10904 2368 10956 2388
rect 10904 2350 10956 2355
rect 10904 2316 10912 2350
rect 10912 2316 10946 2350
rect 10946 2316 10956 2350
rect 10904 2303 10956 2316
rect 6576 2177 6628 2229
rect 6640 2223 6692 2229
rect 6704 2223 6756 2229
rect 6640 2189 6663 2223
rect 6663 2189 6692 2223
rect 6704 2189 6735 2223
rect 6735 2189 6756 2223
rect 6640 2177 6692 2189
rect 6704 2177 6756 2189
rect 6768 2223 6820 2229
rect 6768 2189 6773 2223
rect 6773 2189 6807 2223
rect 6807 2189 6820 2223
rect 6768 2177 6820 2189
rect 6832 2223 6884 2229
rect 6832 2189 6845 2223
rect 6845 2189 6879 2223
rect 6879 2189 6884 2223
rect 6832 2177 6884 2189
rect 6896 2223 6948 2229
rect 6960 2223 7012 2229
rect 7024 2223 7076 2229
rect 7088 2223 7140 2229
rect 7152 2223 7204 2229
rect 7216 2223 7268 2229
rect 7280 2223 7332 2229
rect 6896 2189 6917 2223
rect 6917 2189 6948 2223
rect 6960 2189 6989 2223
rect 6989 2189 7012 2223
rect 7024 2189 7061 2223
rect 7061 2189 7076 2223
rect 7088 2189 7095 2223
rect 7095 2189 7133 2223
rect 7133 2189 7140 2223
rect 7152 2189 7167 2223
rect 7167 2189 7204 2223
rect 7216 2189 7239 2223
rect 7239 2189 7268 2223
rect 7280 2189 7311 2223
rect 7311 2189 7332 2223
rect 6896 2177 6948 2189
rect 6960 2177 7012 2189
rect 7024 2177 7076 2189
rect 7088 2177 7140 2189
rect 7152 2177 7204 2189
rect 7216 2177 7268 2189
rect 7280 2177 7332 2189
rect 7344 2223 7396 2229
rect 7344 2189 7349 2223
rect 7349 2189 7383 2223
rect 7383 2189 7396 2223
rect 7344 2177 7396 2189
rect 7408 2223 7460 2229
rect 7408 2189 7421 2223
rect 7421 2189 7455 2223
rect 7455 2189 7460 2223
rect 7408 2177 7460 2189
rect 7472 2223 7524 2229
rect 7536 2223 7588 2229
rect 7600 2223 7652 2229
rect 7664 2223 7716 2229
rect 7728 2223 7780 2229
rect 7792 2223 7844 2229
rect 7856 2223 7908 2229
rect 7472 2189 7493 2223
rect 7493 2189 7524 2223
rect 7536 2189 7565 2223
rect 7565 2189 7588 2223
rect 7600 2189 7637 2223
rect 7637 2189 7652 2223
rect 7664 2189 7671 2223
rect 7671 2189 7709 2223
rect 7709 2189 7716 2223
rect 7728 2189 7743 2223
rect 7743 2189 7780 2223
rect 7792 2189 7815 2223
rect 7815 2189 7844 2223
rect 7856 2189 7887 2223
rect 7887 2189 7908 2223
rect 7472 2177 7524 2189
rect 7536 2177 7588 2189
rect 7600 2177 7652 2189
rect 7664 2177 7716 2189
rect 7728 2177 7780 2189
rect 7792 2177 7844 2189
rect 7856 2177 7908 2189
rect 7920 2223 7972 2229
rect 7920 2189 7925 2223
rect 7925 2189 7959 2223
rect 7959 2189 7972 2223
rect 7920 2177 7972 2189
rect 7984 2223 8036 2229
rect 7984 2189 7997 2223
rect 7997 2189 8031 2223
rect 8031 2189 8036 2223
rect 7984 2177 8036 2189
rect 8048 2223 8100 2229
rect 8112 2223 8164 2229
rect 8176 2223 8228 2229
rect 8240 2223 8292 2229
rect 8304 2223 8356 2229
rect 8368 2223 8420 2229
rect 8432 2223 8484 2229
rect 8048 2189 8069 2223
rect 8069 2189 8100 2223
rect 8112 2189 8141 2223
rect 8141 2189 8164 2223
rect 8176 2189 8213 2223
rect 8213 2189 8228 2223
rect 8240 2189 8247 2223
rect 8247 2189 8285 2223
rect 8285 2189 8292 2223
rect 8304 2189 8319 2223
rect 8319 2189 8356 2223
rect 8368 2189 8391 2223
rect 8391 2189 8420 2223
rect 8432 2189 8463 2223
rect 8463 2189 8484 2223
rect 8048 2177 8100 2189
rect 8112 2177 8164 2189
rect 8176 2177 8228 2189
rect 8240 2177 8292 2189
rect 8304 2177 8356 2189
rect 8368 2177 8420 2189
rect 8432 2177 8484 2189
rect 8496 2223 8548 2229
rect 8496 2189 8501 2223
rect 8501 2189 8535 2223
rect 8535 2189 8548 2223
rect 8496 2177 8548 2189
rect 8560 2223 8612 2229
rect 8560 2189 8573 2223
rect 8573 2189 8607 2223
rect 8607 2189 8612 2223
rect 8560 2177 8612 2189
rect 8624 2223 8676 2229
rect 8688 2223 8740 2229
rect 8752 2223 8804 2229
rect 8816 2223 8868 2229
rect 8880 2223 8932 2229
rect 8944 2223 8996 2229
rect 9008 2223 9060 2229
rect 8624 2189 8645 2223
rect 8645 2189 8676 2223
rect 8688 2189 8717 2223
rect 8717 2189 8740 2223
rect 8752 2189 8789 2223
rect 8789 2189 8804 2223
rect 8816 2189 8823 2223
rect 8823 2189 8861 2223
rect 8861 2189 8868 2223
rect 8880 2189 8895 2223
rect 8895 2189 8932 2223
rect 8944 2189 8967 2223
rect 8967 2189 8996 2223
rect 9008 2189 9039 2223
rect 9039 2189 9060 2223
rect 8624 2177 8676 2189
rect 8688 2177 8740 2189
rect 8752 2177 8804 2189
rect 8816 2177 8868 2189
rect 8880 2177 8932 2189
rect 8944 2177 8996 2189
rect 9008 2177 9060 2189
rect 9072 2223 9124 2229
rect 9072 2189 9077 2223
rect 9077 2189 9111 2223
rect 9111 2189 9124 2223
rect 9072 2177 9124 2189
rect 9136 2223 9188 2229
rect 9136 2189 9149 2223
rect 9149 2189 9183 2223
rect 9183 2189 9188 2223
rect 9136 2177 9188 2189
rect 9200 2223 9252 2229
rect 9264 2223 9316 2229
rect 9328 2223 9380 2229
rect 9392 2223 9444 2229
rect 9456 2223 9508 2229
rect 9520 2223 9572 2229
rect 9584 2223 9636 2229
rect 9200 2189 9221 2223
rect 9221 2189 9252 2223
rect 9264 2189 9293 2223
rect 9293 2189 9316 2223
rect 9328 2189 9365 2223
rect 9365 2189 9380 2223
rect 9392 2189 9399 2223
rect 9399 2189 9437 2223
rect 9437 2189 9444 2223
rect 9456 2189 9471 2223
rect 9471 2189 9508 2223
rect 9520 2189 9543 2223
rect 9543 2189 9572 2223
rect 9584 2189 9615 2223
rect 9615 2189 9636 2223
rect 9200 2177 9252 2189
rect 9264 2177 9316 2189
rect 9328 2177 9380 2189
rect 9392 2177 9444 2189
rect 9456 2177 9508 2189
rect 9520 2177 9572 2189
rect 9584 2177 9636 2189
rect 9648 2223 9700 2229
rect 9648 2189 9653 2223
rect 9653 2189 9687 2223
rect 9687 2189 9700 2223
rect 9648 2177 9700 2189
rect 9712 2223 9764 2229
rect 9712 2189 9725 2223
rect 9725 2189 9759 2223
rect 9759 2189 9764 2223
rect 9712 2177 9764 2189
rect 9776 2223 9828 2229
rect 9840 2223 9892 2229
rect 9904 2223 9956 2229
rect 9968 2223 10020 2229
rect 10032 2223 10084 2229
rect 10096 2223 10148 2229
rect 10160 2223 10212 2229
rect 9776 2189 9797 2223
rect 9797 2189 9828 2223
rect 9840 2189 9869 2223
rect 9869 2189 9892 2223
rect 9904 2189 9941 2223
rect 9941 2189 9956 2223
rect 9968 2189 9975 2223
rect 9975 2189 10013 2223
rect 10013 2189 10020 2223
rect 10032 2189 10047 2223
rect 10047 2189 10084 2223
rect 10096 2189 10119 2223
rect 10119 2189 10148 2223
rect 10160 2189 10191 2223
rect 10191 2189 10212 2223
rect 9776 2177 9828 2189
rect 9840 2177 9892 2189
rect 9904 2177 9956 2189
rect 9968 2177 10020 2189
rect 10032 2177 10084 2189
rect 10096 2177 10148 2189
rect 10160 2177 10212 2189
rect 10224 2223 10276 2229
rect 10224 2189 10229 2223
rect 10229 2189 10263 2223
rect 10263 2189 10276 2223
rect 10224 2177 10276 2189
rect 10288 2223 10340 2229
rect 10288 2189 10301 2223
rect 10301 2189 10335 2223
rect 10335 2189 10340 2223
rect 10288 2177 10340 2189
rect 10352 2223 10404 2229
rect 10416 2223 10468 2229
rect 10480 2223 10532 2229
rect 10544 2223 10596 2229
rect 10608 2223 10660 2229
rect 10672 2223 10724 2229
rect 10736 2223 10788 2229
rect 10352 2189 10373 2223
rect 10373 2189 10404 2223
rect 10416 2189 10445 2223
rect 10445 2189 10468 2223
rect 10480 2189 10517 2223
rect 10517 2189 10532 2223
rect 10544 2189 10551 2223
rect 10551 2189 10589 2223
rect 10589 2189 10596 2223
rect 10608 2189 10623 2223
rect 10623 2189 10660 2223
rect 10672 2189 10695 2223
rect 10695 2189 10724 2223
rect 10736 2189 10767 2223
rect 10767 2189 10788 2223
rect 10352 2177 10404 2189
rect 10416 2177 10468 2189
rect 10480 2177 10532 2189
rect 10544 2177 10596 2189
rect 10608 2177 10660 2189
rect 10672 2177 10724 2189
rect 10736 2177 10788 2189
rect 10800 2223 10852 2229
rect 10800 2189 10805 2223
rect 10805 2189 10839 2223
rect 10839 2189 10852 2223
rect 10800 2177 10852 2189
rect 10864 2223 10916 2229
rect 10864 2189 10877 2223
rect 10877 2189 10911 2223
rect 10911 2189 10916 2223
rect 10864 2177 10916 2189
rect 6576 2144 6628 2154
rect 6641 2144 6693 2154
rect 6706 2144 6758 2154
rect 6576 2110 6625 2144
rect 6625 2110 6628 2144
rect 6641 2110 6659 2144
rect 6659 2110 6693 2144
rect 6706 2110 6732 2144
rect 6732 2110 6758 2144
rect 6576 2102 6628 2110
rect 6641 2102 6693 2110
rect 6706 2102 6758 2110
rect 6771 2144 6823 2154
rect 6771 2110 6805 2144
rect 6805 2110 6823 2144
rect 6771 2102 6823 2110
rect 6836 2144 6888 2154
rect 6836 2110 6844 2144
rect 6844 2110 6878 2144
rect 6878 2110 6888 2144
rect 6836 2102 6888 2110
rect 6901 2144 6953 2154
rect 6901 2110 6917 2144
rect 6917 2110 6951 2144
rect 6951 2110 6953 2144
rect 6901 2102 6953 2110
rect 6966 2144 7018 2154
rect 7031 2144 7083 2154
rect 7096 2144 7148 2154
rect 7161 2144 7213 2154
rect 7226 2144 7278 2154
rect 7291 2144 7343 2154
rect 6966 2110 6990 2144
rect 6990 2110 7018 2144
rect 7031 2110 7063 2144
rect 7063 2110 7083 2144
rect 7096 2110 7097 2144
rect 7097 2110 7136 2144
rect 7136 2110 7148 2144
rect 7161 2110 7170 2144
rect 7170 2110 7209 2144
rect 7209 2110 7213 2144
rect 7226 2110 7243 2144
rect 7243 2110 7278 2144
rect 7291 2110 7316 2144
rect 7316 2110 7343 2144
rect 6966 2102 7018 2110
rect 7031 2102 7083 2110
rect 7096 2102 7148 2110
rect 7161 2102 7213 2110
rect 7226 2102 7278 2110
rect 7291 2102 7343 2110
rect 7355 2144 7407 2154
rect 7355 2110 7389 2144
rect 7389 2110 7407 2144
rect 7355 2102 7407 2110
rect 7419 2144 7471 2154
rect 7419 2110 7428 2144
rect 7428 2110 7462 2144
rect 7462 2110 7471 2144
rect 7419 2102 7471 2110
rect 7483 2144 7535 2154
rect 7483 2110 7501 2144
rect 7501 2110 7535 2144
rect 7483 2102 7535 2110
rect 7547 2144 7599 2154
rect 7611 2144 7663 2154
rect 7675 2144 7727 2154
rect 7739 2144 7791 2154
rect 7803 2144 7855 2154
rect 7867 2144 7919 2154
rect 7547 2110 7574 2144
rect 7574 2110 7599 2144
rect 7611 2110 7647 2144
rect 7647 2110 7663 2144
rect 7675 2110 7681 2144
rect 7681 2110 7720 2144
rect 7720 2110 7727 2144
rect 7739 2110 7754 2144
rect 7754 2110 7791 2144
rect 7803 2110 7826 2144
rect 7826 2110 7855 2144
rect 7867 2110 7898 2144
rect 7898 2110 7919 2144
rect 7547 2102 7599 2110
rect 7611 2102 7663 2110
rect 7675 2102 7727 2110
rect 7739 2102 7791 2110
rect 7803 2102 7855 2110
rect 7867 2102 7919 2110
rect 7931 2144 7983 2154
rect 7931 2110 7936 2144
rect 7936 2110 7970 2144
rect 7970 2110 7983 2144
rect 7931 2102 7983 2110
rect 7995 2144 8047 2154
rect 7995 2110 8008 2144
rect 8008 2110 8042 2144
rect 8042 2110 8047 2144
rect 7995 2102 8047 2110
rect 8059 2144 8111 2154
rect 8123 2144 8175 2154
rect 8187 2144 8239 2154
rect 8251 2144 8303 2154
rect 8315 2144 8367 2154
rect 8379 2144 8431 2154
rect 8443 2144 8495 2154
rect 8059 2110 8080 2144
rect 8080 2110 8111 2144
rect 8123 2110 8152 2144
rect 8152 2110 8175 2144
rect 8187 2110 8224 2144
rect 8224 2110 8239 2144
rect 8251 2110 8258 2144
rect 8258 2110 8296 2144
rect 8296 2110 8303 2144
rect 8315 2110 8330 2144
rect 8330 2110 8367 2144
rect 8379 2110 8402 2144
rect 8402 2110 8431 2144
rect 8443 2110 8474 2144
rect 8474 2110 8495 2144
rect 8059 2102 8111 2110
rect 8123 2102 8175 2110
rect 8187 2102 8239 2110
rect 8251 2102 8303 2110
rect 8315 2102 8367 2110
rect 8379 2102 8431 2110
rect 8443 2102 8495 2110
rect 8507 2144 8559 2154
rect 8507 2110 8512 2144
rect 8512 2110 8546 2144
rect 8546 2110 8559 2144
rect 8507 2102 8559 2110
rect 8571 2144 8623 2154
rect 8571 2110 8584 2144
rect 8584 2110 8618 2144
rect 8618 2110 8623 2144
rect 8571 2102 8623 2110
rect 8635 2144 8687 2154
rect 8699 2144 8751 2154
rect 8763 2144 8815 2154
rect 8827 2144 8879 2154
rect 8891 2144 8943 2154
rect 8955 2144 9007 2154
rect 9019 2144 9071 2154
rect 8635 2110 8656 2144
rect 8656 2110 8687 2144
rect 8699 2110 8728 2144
rect 8728 2110 8751 2144
rect 8763 2110 8800 2144
rect 8800 2110 8815 2144
rect 8827 2110 8834 2144
rect 8834 2110 8872 2144
rect 8872 2110 8879 2144
rect 8891 2110 8906 2144
rect 8906 2110 8943 2144
rect 8955 2110 8978 2144
rect 8978 2110 9007 2144
rect 9019 2110 9050 2144
rect 9050 2110 9071 2144
rect 8635 2102 8687 2110
rect 8699 2102 8751 2110
rect 8763 2102 8815 2110
rect 8827 2102 8879 2110
rect 8891 2102 8943 2110
rect 8955 2102 9007 2110
rect 9019 2102 9071 2110
rect 9083 2144 9135 2154
rect 9083 2110 9088 2144
rect 9088 2110 9122 2144
rect 9122 2110 9135 2144
rect 9083 2102 9135 2110
rect 9147 2144 9199 2154
rect 9147 2110 9160 2144
rect 9160 2110 9194 2144
rect 9194 2110 9199 2144
rect 9147 2102 9199 2110
rect 9211 2144 9263 2154
rect 9275 2144 9327 2154
rect 9339 2144 9391 2154
rect 9403 2144 9455 2154
rect 9467 2144 9519 2154
rect 9531 2144 9583 2154
rect 9595 2144 9647 2154
rect 9211 2110 9232 2144
rect 9232 2110 9263 2144
rect 9275 2110 9304 2144
rect 9304 2110 9327 2144
rect 9339 2110 9376 2144
rect 9376 2110 9391 2144
rect 9403 2110 9410 2144
rect 9410 2110 9448 2144
rect 9448 2110 9455 2144
rect 9467 2110 9482 2144
rect 9482 2110 9519 2144
rect 9531 2110 9554 2144
rect 9554 2110 9583 2144
rect 9595 2110 9626 2144
rect 9626 2110 9647 2144
rect 9211 2102 9263 2110
rect 9275 2102 9327 2110
rect 9339 2102 9391 2110
rect 9403 2102 9455 2110
rect 9467 2102 9519 2110
rect 9531 2102 9583 2110
rect 9595 2102 9647 2110
rect 9659 2144 9711 2154
rect 9659 2110 9664 2144
rect 9664 2110 9698 2144
rect 9698 2110 9711 2144
rect 9659 2102 9711 2110
rect 9723 2144 9775 2154
rect 9723 2110 9736 2144
rect 9736 2110 9770 2144
rect 9770 2110 9775 2144
rect 9723 2102 9775 2110
rect 9787 2144 9839 2154
rect 9851 2144 9903 2154
rect 9915 2144 9967 2154
rect 9979 2144 10031 2154
rect 10043 2144 10095 2154
rect 10107 2144 10159 2154
rect 10171 2144 10223 2154
rect 9787 2110 9808 2144
rect 9808 2110 9839 2144
rect 9851 2110 9880 2144
rect 9880 2110 9903 2144
rect 9915 2110 9952 2144
rect 9952 2110 9967 2144
rect 9979 2110 9986 2144
rect 9986 2110 10024 2144
rect 10024 2110 10031 2144
rect 10043 2110 10058 2144
rect 10058 2110 10095 2144
rect 10107 2110 10130 2144
rect 10130 2110 10159 2144
rect 10171 2110 10202 2144
rect 10202 2110 10223 2144
rect 9787 2102 9839 2110
rect 9851 2102 9903 2110
rect 9915 2102 9967 2110
rect 9979 2102 10031 2110
rect 10043 2102 10095 2110
rect 10107 2102 10159 2110
rect 10171 2102 10223 2110
rect 10235 2144 10287 2154
rect 10235 2110 10240 2144
rect 10240 2110 10274 2144
rect 10274 2110 10287 2144
rect 10235 2102 10287 2110
rect 10299 2144 10351 2154
rect 10299 2110 10312 2144
rect 10312 2110 10346 2144
rect 10346 2110 10351 2144
rect 10299 2102 10351 2110
rect 10363 2144 10415 2154
rect 10427 2144 10479 2154
rect 10491 2144 10543 2154
rect 10555 2144 10607 2154
rect 10619 2144 10671 2154
rect 10683 2144 10735 2154
rect 10747 2144 10799 2154
rect 10363 2110 10384 2144
rect 10384 2110 10415 2144
rect 10427 2110 10456 2144
rect 10456 2110 10479 2144
rect 10491 2110 10528 2144
rect 10528 2110 10543 2144
rect 10555 2110 10562 2144
rect 10562 2110 10600 2144
rect 10600 2110 10607 2144
rect 10619 2110 10634 2144
rect 10634 2110 10671 2144
rect 10683 2110 10706 2144
rect 10706 2110 10735 2144
rect 10747 2110 10778 2144
rect 10778 2110 10799 2144
rect 10363 2102 10415 2110
rect 10427 2102 10479 2110
rect 10491 2102 10543 2110
rect 10555 2102 10607 2110
rect 10619 2102 10671 2110
rect 10683 2102 10735 2110
rect 10747 2102 10799 2110
rect 10811 2144 10863 2154
rect 10811 2110 10816 2144
rect 10816 2110 10850 2144
rect 10850 2110 10863 2144
rect 10811 2102 10863 2110
rect 10875 2144 10927 2154
rect 10875 2110 10888 2144
rect 10888 2110 10922 2144
rect 10922 2110 10927 2144
rect 10875 2102 10927 2110
rect 6582 2069 6634 2075
rect 6646 2069 6698 2075
rect 6710 2069 6762 2075
rect 6774 2069 6826 2075
rect 6582 2035 6629 2069
rect 6629 2035 6634 2069
rect 6646 2035 6663 2069
rect 6663 2035 6698 2069
rect 6710 2035 6735 2069
rect 6735 2035 6762 2069
rect 6774 2035 6807 2069
rect 6807 2035 6826 2069
rect 6582 2023 6634 2035
rect 6646 2023 6698 2035
rect 6710 2023 6762 2035
rect 6774 2023 6826 2035
rect 6838 2069 6890 2075
rect 6838 2035 6845 2069
rect 6845 2035 6879 2069
rect 6879 2035 6890 2069
rect 6838 2023 6890 2035
rect 6902 2069 6954 2075
rect 6902 2035 6917 2069
rect 6917 2035 6951 2069
rect 6951 2035 6954 2069
rect 6902 2023 6954 2035
rect 6966 2069 7018 2075
rect 7030 2069 7082 2075
rect 7094 2069 7146 2075
rect 7158 2069 7210 2075
rect 7222 2069 7274 2075
rect 7286 2069 7338 2075
rect 7350 2069 7402 2075
rect 6966 2035 6989 2069
rect 6989 2035 7018 2069
rect 7030 2035 7061 2069
rect 7061 2035 7082 2069
rect 7094 2035 7095 2069
rect 7095 2035 7133 2069
rect 7133 2035 7146 2069
rect 7158 2035 7167 2069
rect 7167 2035 7205 2069
rect 7205 2035 7210 2069
rect 7222 2035 7239 2069
rect 7239 2035 7274 2069
rect 7286 2035 7311 2069
rect 7311 2035 7338 2069
rect 7350 2035 7383 2069
rect 7383 2035 7402 2069
rect 6966 2023 7018 2035
rect 7030 2023 7082 2035
rect 7094 2023 7146 2035
rect 7158 2023 7210 2035
rect 7222 2023 7274 2035
rect 7286 2023 7338 2035
rect 7350 2023 7402 2035
rect 7414 2069 7466 2075
rect 7414 2035 7421 2069
rect 7421 2035 7455 2069
rect 7455 2035 7466 2069
rect 7414 2023 7466 2035
rect 7478 2069 7530 2075
rect 7478 2035 7493 2069
rect 7493 2035 7527 2069
rect 7527 2035 7530 2069
rect 7478 2023 7530 2035
rect 7542 2069 7594 2075
rect 7606 2069 7658 2075
rect 7670 2069 7722 2075
rect 7734 2069 7786 2075
rect 7798 2069 7850 2075
rect 7862 2069 7914 2075
rect 7926 2069 7978 2075
rect 7542 2035 7565 2069
rect 7565 2035 7594 2069
rect 7606 2035 7637 2069
rect 7637 2035 7658 2069
rect 7670 2035 7671 2069
rect 7671 2035 7709 2069
rect 7709 2035 7722 2069
rect 7734 2035 7743 2069
rect 7743 2035 7781 2069
rect 7781 2035 7786 2069
rect 7798 2035 7815 2069
rect 7815 2035 7850 2069
rect 7862 2035 7887 2069
rect 7887 2035 7914 2069
rect 7926 2035 7959 2069
rect 7959 2035 7978 2069
rect 7542 2023 7594 2035
rect 7606 2023 7658 2035
rect 7670 2023 7722 2035
rect 7734 2023 7786 2035
rect 7798 2023 7850 2035
rect 7862 2023 7914 2035
rect 7926 2023 7978 2035
rect 7990 2069 8042 2075
rect 7990 2035 7997 2069
rect 7997 2035 8031 2069
rect 8031 2035 8042 2069
rect 7990 2023 8042 2035
rect 8054 2069 8106 2075
rect 8054 2035 8069 2069
rect 8069 2035 8103 2069
rect 8103 2035 8106 2069
rect 8054 2023 8106 2035
rect 8118 2069 8170 2075
rect 8182 2069 8234 2075
rect 8246 2069 8298 2075
rect 8310 2069 8362 2075
rect 8374 2069 8426 2075
rect 8438 2069 8490 2075
rect 8502 2069 8554 2075
rect 8118 2035 8141 2069
rect 8141 2035 8170 2069
rect 8182 2035 8213 2069
rect 8213 2035 8234 2069
rect 8246 2035 8247 2069
rect 8247 2035 8285 2069
rect 8285 2035 8298 2069
rect 8310 2035 8319 2069
rect 8319 2035 8357 2069
rect 8357 2035 8362 2069
rect 8374 2035 8391 2069
rect 8391 2035 8426 2069
rect 8438 2035 8463 2069
rect 8463 2035 8490 2069
rect 8502 2035 8535 2069
rect 8535 2035 8554 2069
rect 8118 2023 8170 2035
rect 8182 2023 8234 2035
rect 8246 2023 8298 2035
rect 8310 2023 8362 2035
rect 8374 2023 8426 2035
rect 8438 2023 8490 2035
rect 8502 2023 8554 2035
rect 8566 2069 8618 2075
rect 8566 2035 8573 2069
rect 8573 2035 8607 2069
rect 8607 2035 8618 2069
rect 8566 2023 8618 2035
rect 8630 2069 8682 2075
rect 8630 2035 8645 2069
rect 8645 2035 8679 2069
rect 8679 2035 8682 2069
rect 8630 2023 8682 2035
rect 8694 2069 8746 2075
rect 8758 2069 8810 2075
rect 8822 2069 8874 2075
rect 8886 2069 8938 2075
rect 8950 2069 9002 2075
rect 9014 2069 9066 2075
rect 9078 2069 9130 2075
rect 8694 2035 8717 2069
rect 8717 2035 8746 2069
rect 8758 2035 8789 2069
rect 8789 2035 8810 2069
rect 8822 2035 8823 2069
rect 8823 2035 8861 2069
rect 8861 2035 8874 2069
rect 8886 2035 8895 2069
rect 8895 2035 8933 2069
rect 8933 2035 8938 2069
rect 8950 2035 8967 2069
rect 8967 2035 9002 2069
rect 9014 2035 9039 2069
rect 9039 2035 9066 2069
rect 9078 2035 9111 2069
rect 9111 2035 9130 2069
rect 8694 2023 8746 2035
rect 8758 2023 8810 2035
rect 8822 2023 8874 2035
rect 8886 2023 8938 2035
rect 8950 2023 9002 2035
rect 9014 2023 9066 2035
rect 9078 2023 9130 2035
rect 9142 2069 9194 2075
rect 9142 2035 9149 2069
rect 9149 2035 9183 2069
rect 9183 2035 9194 2069
rect 9142 2023 9194 2035
rect 9206 2069 9258 2075
rect 9206 2035 9221 2069
rect 9221 2035 9255 2069
rect 9255 2035 9258 2069
rect 9206 2023 9258 2035
rect 9270 2069 9322 2075
rect 9334 2069 9386 2075
rect 9398 2069 9450 2075
rect 9462 2069 9514 2075
rect 9526 2069 9578 2075
rect 9590 2069 9642 2075
rect 9654 2069 9706 2075
rect 9270 2035 9293 2069
rect 9293 2035 9322 2069
rect 9334 2035 9365 2069
rect 9365 2035 9386 2069
rect 9398 2035 9399 2069
rect 9399 2035 9437 2069
rect 9437 2035 9450 2069
rect 9462 2035 9471 2069
rect 9471 2035 9509 2069
rect 9509 2035 9514 2069
rect 9526 2035 9543 2069
rect 9543 2035 9578 2069
rect 9590 2035 9615 2069
rect 9615 2035 9642 2069
rect 9654 2035 9687 2069
rect 9687 2035 9706 2069
rect 9270 2023 9322 2035
rect 9334 2023 9386 2035
rect 9398 2023 9450 2035
rect 9462 2023 9514 2035
rect 9526 2023 9578 2035
rect 9590 2023 9642 2035
rect 9654 2023 9706 2035
rect 9718 2069 9770 2075
rect 9718 2035 9725 2069
rect 9725 2035 9759 2069
rect 9759 2035 9770 2069
rect 9718 2023 9770 2035
rect 9782 2069 9834 2075
rect 9782 2035 9797 2069
rect 9797 2035 9831 2069
rect 9831 2035 9834 2069
rect 9782 2023 9834 2035
rect 9846 2069 9898 2075
rect 9910 2069 9962 2075
rect 9974 2069 10026 2075
rect 10038 2069 10090 2075
rect 10102 2069 10154 2075
rect 10166 2069 10218 2075
rect 10230 2069 10282 2075
rect 9846 2035 9869 2069
rect 9869 2035 9898 2069
rect 9910 2035 9941 2069
rect 9941 2035 9962 2069
rect 9974 2035 9975 2069
rect 9975 2035 10013 2069
rect 10013 2035 10026 2069
rect 10038 2035 10047 2069
rect 10047 2035 10085 2069
rect 10085 2035 10090 2069
rect 10102 2035 10119 2069
rect 10119 2035 10154 2069
rect 10166 2035 10191 2069
rect 10191 2035 10218 2069
rect 10230 2035 10263 2069
rect 10263 2035 10282 2069
rect 9846 2023 9898 2035
rect 9910 2023 9962 2035
rect 9974 2023 10026 2035
rect 10038 2023 10090 2035
rect 10102 2023 10154 2035
rect 10166 2023 10218 2035
rect 10230 2023 10282 2035
rect 10294 2069 10346 2075
rect 10294 2035 10301 2069
rect 10301 2035 10335 2069
rect 10335 2035 10346 2069
rect 10294 2023 10346 2035
rect 10358 2069 10410 2075
rect 10358 2035 10373 2069
rect 10373 2035 10407 2069
rect 10407 2035 10410 2069
rect 10358 2023 10410 2035
rect 10422 2069 10474 2075
rect 10486 2069 10538 2075
rect 10550 2069 10602 2075
rect 10614 2069 10666 2075
rect 10678 2069 10730 2075
rect 10742 2069 10794 2075
rect 10806 2069 10858 2075
rect 10422 2035 10445 2069
rect 10445 2035 10474 2069
rect 10486 2035 10517 2069
rect 10517 2035 10538 2069
rect 10550 2035 10551 2069
rect 10551 2035 10589 2069
rect 10589 2035 10602 2069
rect 10614 2035 10623 2069
rect 10623 2035 10661 2069
rect 10661 2035 10666 2069
rect 10678 2035 10695 2069
rect 10695 2035 10730 2069
rect 10742 2035 10767 2069
rect 10767 2035 10794 2069
rect 10806 2035 10839 2069
rect 10839 2035 10858 2069
rect 10422 2023 10474 2035
rect 10486 2023 10538 2035
rect 10550 2023 10602 2035
rect 10614 2023 10666 2035
rect 10678 2023 10730 2035
rect 10742 2023 10794 2035
rect 10806 2023 10858 2035
rect 10870 2069 10922 2075
rect 10870 2035 10877 2069
rect 10877 2035 10911 2069
rect 10911 2035 10922 2069
rect 10870 2023 10922 2035
rect 11619 5872 11671 5882
rect 11619 5838 11624 5872
rect 11624 5838 11658 5872
rect 11658 5838 11671 5872
rect 11619 5830 11671 5838
rect 11683 5872 11735 5882
rect 11683 5838 11696 5872
rect 11696 5838 11730 5872
rect 11730 5838 11735 5872
rect 11683 5830 11735 5838
rect 14355 5845 14407 5897
rect 14419 5845 14471 5897
rect 11619 5734 11671 5743
rect 11619 5700 11624 5734
rect 11624 5700 11658 5734
rect 11658 5700 11671 5734
rect 11619 5691 11671 5700
rect 11683 5734 11735 5743
rect 11683 5700 11696 5734
rect 11696 5700 11730 5734
rect 11730 5700 11735 5734
rect 11683 5691 11735 5700
rect 14359 5691 14411 5743
rect 14423 5691 14475 5743
rect 11619 5580 11671 5589
rect 11619 5546 11624 5580
rect 11624 5546 11658 5580
rect 11658 5546 11671 5580
rect 11619 5537 11671 5546
rect 11683 5580 11735 5589
rect 11683 5546 11696 5580
rect 11696 5546 11730 5580
rect 11730 5546 11735 5580
rect 11683 5537 11735 5546
rect 14355 5537 14407 5589
rect 14419 5537 14471 5589
rect 11619 5426 11671 5435
rect 11619 5392 11624 5426
rect 11624 5392 11658 5426
rect 11658 5392 11671 5426
rect 11619 5383 11671 5392
rect 11683 5426 11735 5435
rect 11683 5392 11696 5426
rect 11696 5392 11730 5426
rect 11730 5392 11735 5426
rect 11683 5383 11735 5392
rect 14359 5383 14411 5435
rect 14423 5383 14475 5435
rect 11619 5272 11671 5281
rect 11619 5238 11624 5272
rect 11624 5238 11658 5272
rect 11658 5238 11671 5272
rect 11619 5229 11671 5238
rect 11683 5272 11735 5281
rect 11683 5238 11696 5272
rect 11696 5238 11730 5272
rect 11730 5238 11735 5272
rect 11683 5229 11735 5238
rect 14355 5229 14407 5281
rect 14419 5229 14471 5281
rect 11619 5118 11671 5127
rect 11619 5084 11624 5118
rect 11624 5084 11658 5118
rect 11658 5084 11671 5118
rect 11619 5075 11671 5084
rect 11683 5118 11735 5127
rect 11683 5084 11696 5118
rect 11696 5084 11730 5118
rect 11730 5084 11735 5118
rect 11683 5075 11735 5084
rect 14359 5075 14411 5127
rect 14423 5075 14475 5127
rect 11619 4964 11671 4973
rect 11619 4930 11624 4964
rect 11624 4930 11658 4964
rect 11658 4930 11671 4964
rect 11619 4921 11671 4930
rect 11683 4964 11735 4973
rect 11683 4930 11696 4964
rect 11696 4930 11730 4964
rect 11730 4930 11735 4964
rect 11683 4921 11735 4930
rect 14355 4921 14407 4973
rect 14419 4921 14471 4973
rect 11619 4810 11671 4819
rect 11619 4776 11624 4810
rect 11624 4776 11658 4810
rect 11658 4776 11671 4810
rect 11619 4767 11671 4776
rect 11683 4810 11735 4819
rect 11683 4776 11696 4810
rect 11696 4776 11730 4810
rect 11730 4776 11735 4810
rect 11683 4767 11735 4776
rect 14359 4767 14411 4819
rect 14423 4767 14475 4819
rect 11619 4656 11671 4665
rect 11619 4622 11624 4656
rect 11624 4622 11658 4656
rect 11658 4622 11671 4656
rect 11619 4613 11671 4622
rect 11683 4656 11735 4665
rect 11683 4622 11696 4656
rect 11696 4622 11730 4656
rect 11730 4622 11735 4656
rect 11683 4613 11735 4622
rect 14355 4613 14407 4665
rect 14419 4613 14471 4665
rect 11619 4502 11671 4511
rect 11619 4468 11624 4502
rect 11624 4468 11658 4502
rect 11658 4468 11671 4502
rect 11619 4459 11671 4468
rect 11683 4502 11735 4511
rect 11683 4468 11696 4502
rect 11696 4468 11730 4502
rect 11730 4468 11735 4502
rect 11683 4459 11735 4468
rect 14359 4459 14411 4511
rect 14423 4459 14475 4511
rect 11619 4348 11671 4357
rect 11619 4314 11624 4348
rect 11624 4314 11658 4348
rect 11658 4314 11671 4348
rect 11619 4305 11671 4314
rect 11683 4348 11735 4357
rect 11683 4314 11696 4348
rect 11696 4314 11730 4348
rect 11730 4314 11735 4348
rect 11683 4305 11735 4314
rect 14355 4305 14407 4357
rect 14419 4305 14471 4357
rect 11619 4194 11671 4203
rect 11619 4160 11624 4194
rect 11624 4160 11658 4194
rect 11658 4160 11671 4194
rect 11619 4151 11671 4160
rect 11683 4194 11735 4203
rect 11683 4160 11696 4194
rect 11696 4160 11730 4194
rect 11730 4160 11735 4194
rect 11683 4151 11735 4160
rect 14359 4151 14411 4203
rect 14423 4151 14475 4203
rect 11619 3908 11671 3917
rect 11619 3874 11624 3908
rect 11624 3874 11658 3908
rect 11658 3874 11671 3908
rect 11619 3865 11671 3874
rect 11683 3908 11735 3917
rect 11683 3874 11696 3908
rect 11696 3874 11730 3908
rect 11730 3874 11735 3908
rect 11683 3865 11735 3874
rect 14359 3865 14411 3917
rect 14423 3865 14475 3917
rect 15173 3865 15225 3917
rect 15237 3865 15289 3917
rect 11619 3754 11671 3763
rect 11619 3720 11624 3754
rect 11624 3720 11658 3754
rect 11658 3720 11671 3754
rect 11619 3711 11671 3720
rect 11683 3754 11735 3763
rect 11683 3720 11696 3754
rect 11696 3720 11730 3754
rect 11730 3720 11735 3754
rect 11683 3711 11735 3720
rect 14355 3711 14407 3763
rect 14419 3711 14471 3763
rect 15005 3711 15057 3763
rect 15069 3711 15121 3763
rect 11619 3600 11671 3609
rect 11619 3566 11624 3600
rect 11624 3566 11658 3600
rect 11658 3566 11671 3600
rect 11619 3557 11671 3566
rect 11683 3600 11735 3609
rect 11683 3566 11696 3600
rect 11696 3566 11730 3600
rect 11730 3566 11735 3600
rect 11683 3557 11735 3566
rect 14359 3557 14411 3609
rect 14423 3557 14475 3609
rect 11619 3446 11671 3455
rect 11619 3412 11624 3446
rect 11624 3412 11658 3446
rect 11658 3412 11671 3446
rect 11619 3403 11671 3412
rect 11683 3446 11735 3455
rect 11683 3412 11696 3446
rect 11696 3412 11730 3446
rect 11730 3412 11735 3446
rect 11683 3403 11735 3412
rect 14355 3403 14407 3455
rect 14419 3403 14471 3455
rect 11619 3292 11671 3301
rect 11619 3258 11624 3292
rect 11624 3258 11658 3292
rect 11658 3258 11671 3292
rect 11619 3249 11671 3258
rect 11683 3292 11735 3301
rect 11683 3258 11696 3292
rect 11696 3258 11730 3292
rect 11730 3258 11735 3292
rect 11683 3249 11735 3258
rect 14359 3249 14411 3301
rect 14423 3249 14475 3301
rect 11619 3138 11671 3147
rect 11619 3104 11624 3138
rect 11624 3104 11658 3138
rect 11658 3104 11671 3138
rect 11619 3095 11671 3104
rect 11683 3138 11735 3147
rect 11683 3104 11696 3138
rect 11696 3104 11730 3138
rect 11730 3104 11735 3138
rect 11683 3095 11735 3104
rect 14355 3095 14407 3147
rect 14419 3095 14471 3147
rect 11619 2984 11671 2993
rect 11619 2950 11624 2984
rect 11624 2950 11658 2984
rect 11658 2950 11671 2984
rect 11619 2941 11671 2950
rect 11683 2984 11735 2993
rect 11683 2950 11696 2984
rect 11696 2950 11730 2984
rect 11730 2950 11735 2984
rect 11683 2941 11735 2950
rect 14359 2941 14411 2993
rect 14423 2941 14475 2993
rect 11619 2830 11671 2839
rect 11619 2796 11624 2830
rect 11624 2796 11658 2830
rect 11658 2796 11671 2830
rect 11619 2787 11671 2796
rect 11683 2830 11735 2839
rect 11683 2796 11696 2830
rect 11696 2796 11730 2830
rect 11730 2796 11735 2830
rect 11683 2787 11735 2796
rect 14355 2787 14407 2839
rect 14419 2787 14471 2839
rect 11619 2676 11671 2685
rect 11619 2642 11624 2676
rect 11624 2642 11658 2676
rect 11658 2642 11671 2676
rect 11619 2633 11671 2642
rect 11683 2676 11735 2685
rect 11683 2642 11696 2676
rect 11696 2642 11730 2676
rect 11730 2642 11735 2676
rect 11683 2633 11735 2642
rect 14359 2633 14411 2685
rect 14423 2633 14475 2685
rect 11619 2522 11671 2531
rect 11619 2488 11624 2522
rect 11624 2488 11658 2522
rect 11658 2488 11671 2522
rect 11619 2479 11671 2488
rect 11683 2522 11735 2531
rect 11683 2488 11696 2522
rect 11696 2488 11730 2522
rect 11730 2488 11735 2522
rect 11683 2479 11735 2488
rect 14355 2479 14407 2531
rect 14419 2479 14471 2531
rect 11619 2368 11671 2377
rect 11619 2334 11624 2368
rect 11624 2334 11658 2368
rect 11658 2334 11671 2368
rect 11619 2325 11671 2334
rect 11683 2368 11735 2377
rect 11683 2334 11696 2368
rect 11696 2334 11730 2368
rect 11730 2334 11735 2368
rect 11683 2325 11735 2334
rect 14359 2325 14411 2377
rect 14423 2325 14475 2377
rect 11619 2214 11671 2223
rect 11619 2180 11624 2214
rect 11624 2180 11658 2214
rect 11658 2180 11671 2214
rect 11619 2171 11671 2180
rect 11683 2214 11735 2223
rect 11683 2180 11696 2214
rect 11696 2180 11730 2214
rect 11730 2180 11735 2214
rect 11683 2171 11735 2180
rect 14355 2171 14407 2223
rect 14419 2171 14471 2223
rect 11585 2069 11637 2078
rect 11649 2069 11701 2078
rect 11713 2069 11765 2078
rect 11777 2069 11829 2078
rect 11841 2069 11893 2078
rect 11905 2069 11957 2078
rect 11969 2069 12021 2078
rect 11585 2035 11608 2069
rect 11608 2035 11637 2069
rect 11649 2035 11680 2069
rect 11680 2035 11701 2069
rect 11713 2035 11714 2069
rect 11714 2035 11752 2069
rect 11752 2035 11765 2069
rect 11777 2035 11786 2069
rect 11786 2035 11824 2069
rect 11824 2035 11829 2069
rect 11841 2035 11858 2069
rect 11858 2035 11893 2069
rect 11905 2035 11930 2069
rect 11930 2035 11957 2069
rect 11969 2035 12002 2069
rect 12002 2035 12021 2069
rect 11585 2026 11637 2035
rect 11649 2026 11701 2035
rect 11713 2026 11765 2035
rect 11777 2026 11829 2035
rect 11841 2026 11893 2035
rect 11905 2026 11957 2035
rect 11969 2026 12021 2035
rect 12033 2069 12085 2078
rect 12033 2035 12040 2069
rect 12040 2035 12074 2069
rect 12074 2035 12085 2069
rect 12033 2026 12085 2035
rect 12097 2069 12149 2078
rect 12097 2035 12112 2069
rect 12112 2035 12146 2069
rect 12146 2035 12149 2069
rect 12097 2026 12149 2035
rect 12161 2069 12213 2078
rect 12225 2069 12277 2078
rect 12289 2069 12341 2078
rect 12353 2069 12405 2078
rect 12417 2069 12469 2078
rect 12481 2069 12533 2078
rect 12545 2069 12597 2078
rect 12161 2035 12184 2069
rect 12184 2035 12213 2069
rect 12225 2035 12256 2069
rect 12256 2035 12277 2069
rect 12289 2035 12290 2069
rect 12290 2035 12328 2069
rect 12328 2035 12341 2069
rect 12353 2035 12362 2069
rect 12362 2035 12400 2069
rect 12400 2035 12405 2069
rect 12417 2035 12434 2069
rect 12434 2035 12469 2069
rect 12481 2035 12506 2069
rect 12506 2035 12533 2069
rect 12545 2035 12578 2069
rect 12578 2035 12597 2069
rect 12161 2026 12213 2035
rect 12225 2026 12277 2035
rect 12289 2026 12341 2035
rect 12353 2026 12405 2035
rect 12417 2026 12469 2035
rect 12481 2026 12533 2035
rect 12545 2026 12597 2035
rect 12609 2069 12661 2078
rect 12609 2035 12616 2069
rect 12616 2035 12650 2069
rect 12650 2035 12661 2069
rect 12609 2026 12661 2035
rect 12673 2069 12725 2078
rect 12673 2035 12688 2069
rect 12688 2035 12722 2069
rect 12722 2035 12725 2069
rect 12673 2026 12725 2035
rect 12737 2069 12789 2078
rect 12801 2069 12853 2078
rect 12865 2069 12917 2078
rect 12929 2069 12981 2078
rect 12993 2069 13045 2078
rect 13057 2069 13109 2078
rect 13121 2069 13173 2078
rect 12737 2035 12760 2069
rect 12760 2035 12789 2069
rect 12801 2035 12832 2069
rect 12832 2035 12853 2069
rect 12865 2035 12866 2069
rect 12866 2035 12904 2069
rect 12904 2035 12917 2069
rect 12929 2035 12938 2069
rect 12938 2035 12976 2069
rect 12976 2035 12981 2069
rect 12993 2035 13010 2069
rect 13010 2035 13045 2069
rect 13057 2035 13082 2069
rect 13082 2035 13109 2069
rect 13121 2035 13154 2069
rect 13154 2035 13173 2069
rect 12737 2026 12789 2035
rect 12801 2026 12853 2035
rect 12865 2026 12917 2035
rect 12929 2026 12981 2035
rect 12993 2026 13045 2035
rect 13057 2026 13109 2035
rect 13121 2026 13173 2035
rect 13185 2069 13237 2078
rect 13185 2035 13192 2069
rect 13192 2035 13226 2069
rect 13226 2035 13237 2069
rect 13185 2026 13237 2035
rect 13249 2069 13301 2078
rect 13249 2035 13264 2069
rect 13264 2035 13298 2069
rect 13298 2035 13301 2069
rect 13249 2026 13301 2035
rect 13313 2069 13365 2078
rect 13377 2069 13429 2078
rect 13441 2069 13493 2078
rect 13505 2069 13557 2078
rect 13569 2069 13621 2078
rect 13633 2069 13685 2078
rect 13697 2069 13749 2078
rect 13313 2035 13336 2069
rect 13336 2035 13365 2069
rect 13377 2035 13408 2069
rect 13408 2035 13429 2069
rect 13441 2035 13442 2069
rect 13442 2035 13480 2069
rect 13480 2035 13493 2069
rect 13505 2035 13514 2069
rect 13514 2035 13552 2069
rect 13552 2035 13557 2069
rect 13569 2035 13586 2069
rect 13586 2035 13621 2069
rect 13633 2035 13658 2069
rect 13658 2035 13685 2069
rect 13697 2035 13730 2069
rect 13730 2035 13749 2069
rect 13313 2026 13365 2035
rect 13377 2026 13429 2035
rect 13441 2026 13493 2035
rect 13505 2026 13557 2035
rect 13569 2026 13621 2035
rect 13633 2026 13685 2035
rect 13697 2026 13749 2035
rect 13761 2069 13813 2078
rect 13761 2035 13768 2069
rect 13768 2035 13802 2069
rect 13802 2035 13813 2069
rect 13761 2026 13813 2035
rect 13825 2069 13877 2078
rect 13825 2035 13840 2069
rect 13840 2035 13874 2069
rect 13874 2035 13877 2069
rect 13825 2026 13877 2035
rect 13889 2069 13941 2078
rect 13953 2069 14005 2078
rect 14017 2069 14069 2078
rect 14081 2069 14133 2078
rect 14145 2069 14197 2078
rect 14209 2069 14261 2078
rect 14273 2069 14325 2078
rect 13889 2035 13912 2069
rect 13912 2035 13941 2069
rect 13953 2035 13984 2069
rect 13984 2035 14005 2069
rect 14017 2035 14018 2069
rect 14018 2035 14056 2069
rect 14056 2035 14069 2069
rect 14081 2035 14090 2069
rect 14090 2035 14128 2069
rect 14128 2035 14133 2069
rect 14145 2035 14162 2069
rect 14162 2035 14197 2069
rect 14209 2035 14234 2069
rect 14234 2035 14261 2069
rect 14273 2035 14306 2069
rect 14306 2035 14325 2069
rect 13889 2026 13941 2035
rect 13953 2026 14005 2035
rect 14017 2026 14069 2035
rect 14081 2026 14133 2035
rect 14145 2026 14197 2035
rect 14209 2026 14261 2035
rect 14273 2026 14325 2035
rect 14337 2069 14389 2078
rect 14337 2035 14344 2069
rect 14344 2035 14378 2069
rect 14378 2035 14389 2069
rect 14337 2026 14389 2035
rect 14401 2069 14453 2078
rect 14401 2035 14416 2069
rect 14416 2035 14450 2069
rect 14450 2035 14453 2069
rect 14401 2026 14453 2035
rect 14465 2069 14517 2078
rect 14529 2069 14581 2078
rect 14593 2069 14645 2078
rect 14657 2069 14709 2078
rect 14721 2069 14773 2078
rect 14465 2035 14488 2069
rect 14488 2035 14517 2069
rect 14529 2035 14560 2069
rect 14560 2035 14581 2069
rect 14593 2035 14594 2069
rect 14594 2035 14632 2069
rect 14632 2035 14645 2069
rect 14657 2035 14666 2069
rect 14666 2035 14704 2069
rect 14704 2035 14709 2069
rect 14721 2035 14738 2069
rect 14738 2035 14773 2069
rect 14465 2026 14517 2035
rect 14529 2026 14581 2035
rect 14593 2026 14645 2035
rect 14657 2026 14709 2035
rect 14721 2026 14773 2035
rect 13254 1847 13306 1856
rect 13322 1847 13374 1856
rect 13254 1813 13278 1847
rect 13278 1813 13306 1847
rect 13322 1813 13354 1847
rect 13354 1813 13374 1847
rect 13254 1804 13306 1813
rect 13322 1804 13374 1813
rect 13390 1847 13442 1856
rect 13390 1813 13396 1847
rect 13396 1813 13430 1847
rect 13430 1813 13442 1847
rect 13390 1804 13442 1813
rect 13458 1847 13510 1856
rect 13458 1813 13472 1847
rect 13472 1813 13506 1847
rect 13506 1813 13510 1847
rect 13458 1804 13510 1813
rect 13526 1847 13578 1856
rect 13594 1847 13646 1856
rect 13662 1847 13714 1856
rect 13730 1847 13782 1856
rect 13526 1813 13548 1847
rect 13548 1813 13578 1847
rect 13594 1813 13624 1847
rect 13624 1813 13646 1847
rect 13662 1813 13700 1847
rect 13700 1813 13714 1847
rect 13730 1813 13734 1847
rect 13734 1813 13776 1847
rect 13776 1813 13782 1847
rect 13526 1804 13578 1813
rect 13594 1804 13646 1813
rect 13662 1804 13714 1813
rect 13730 1804 13782 1813
rect 10789 1727 10841 1779
rect 10853 1727 10905 1779
rect 10789 1419 10841 1471
rect 10853 1419 10905 1471
rect 13254 1385 13306 1394
rect 13322 1385 13374 1394
rect 13254 1351 13278 1385
rect 13278 1351 13306 1385
rect 13322 1351 13354 1385
rect 13354 1351 13374 1385
rect 13254 1342 13306 1351
rect 13322 1342 13374 1351
rect 13390 1385 13442 1394
rect 13390 1351 13396 1385
rect 13396 1351 13430 1385
rect 13430 1351 13442 1385
rect 13390 1342 13442 1351
rect 13458 1385 13510 1394
rect 13458 1351 13472 1385
rect 13472 1351 13506 1385
rect 13506 1351 13510 1385
rect 13458 1342 13510 1351
rect 13526 1385 13578 1394
rect 13594 1385 13646 1394
rect 13662 1385 13714 1394
rect 13730 1385 13782 1394
rect 13526 1351 13548 1385
rect 13548 1351 13578 1385
rect 13594 1351 13624 1385
rect 13624 1351 13646 1385
rect 13662 1351 13700 1385
rect 13700 1351 13714 1385
rect 13730 1351 13734 1385
rect 13734 1351 13776 1385
rect 13776 1351 13782 1385
rect 13526 1342 13578 1351
rect 13594 1342 13646 1351
rect 13662 1342 13714 1351
rect 13730 1342 13782 1351
rect 10789 1111 10841 1163
rect 10853 1111 10905 1163
rect 13254 1077 13306 1086
rect 13322 1077 13374 1086
rect 13254 1043 13278 1077
rect 13278 1043 13306 1077
rect 13322 1043 13354 1077
rect 13354 1043 13374 1077
rect 13254 1034 13306 1043
rect 13322 1034 13374 1043
rect 13390 1077 13442 1086
rect 13390 1043 13396 1077
rect 13396 1043 13430 1077
rect 13430 1043 13442 1077
rect 13390 1034 13442 1043
rect 13458 1077 13510 1086
rect 13458 1043 13472 1077
rect 13472 1043 13506 1077
rect 13506 1043 13510 1077
rect 13458 1034 13510 1043
rect 13526 1077 13578 1086
rect 13594 1077 13646 1086
rect 13662 1077 13714 1086
rect 13730 1077 13782 1086
rect 13526 1043 13548 1077
rect 13548 1043 13578 1077
rect 13594 1043 13624 1077
rect 13624 1043 13646 1077
rect 13662 1043 13700 1077
rect 13700 1043 13714 1077
rect 13730 1043 13734 1077
rect 13734 1043 13776 1077
rect 13776 1043 13782 1077
rect 13526 1034 13578 1043
rect 13594 1034 13646 1043
rect 13662 1034 13714 1043
rect 13730 1034 13782 1043
rect 10789 803 10841 855
rect 10853 803 10905 855
rect 13254 769 13306 778
rect 13322 769 13374 778
rect 13254 735 13278 769
rect 13278 735 13306 769
rect 13322 735 13354 769
rect 13354 735 13374 769
rect 13254 726 13306 735
rect 13322 726 13374 735
rect 13390 769 13442 778
rect 13390 735 13396 769
rect 13396 735 13430 769
rect 13430 735 13442 769
rect 13390 726 13442 735
rect 13458 769 13510 778
rect 13458 735 13472 769
rect 13472 735 13506 769
rect 13506 735 13510 769
rect 13458 726 13510 735
rect 13526 769 13578 778
rect 13594 769 13646 778
rect 13662 769 13714 778
rect 13730 769 13782 778
rect 13526 735 13548 769
rect 13548 735 13578 769
rect 13594 735 13624 769
rect 13624 735 13646 769
rect 13662 735 13700 769
rect 13700 735 13714 769
rect 13730 735 13734 769
rect 13734 735 13776 769
rect 13776 735 13782 769
rect 13526 726 13578 735
rect 13594 726 13646 735
rect 13662 726 13714 735
rect 13730 726 13782 735
rect 10789 495 10841 547
rect 10853 495 10905 547
rect 6451 341 6503 393
rect 6515 341 6567 393
rect 13162 461 13214 470
rect 13162 427 13168 461
rect 13168 427 13202 461
rect 13202 427 13214 461
rect 13162 418 13214 427
rect 13232 461 13284 470
rect 13232 427 13241 461
rect 13241 427 13275 461
rect 13275 427 13284 461
rect 13232 418 13284 427
rect 13302 461 13354 470
rect 13302 427 13314 461
rect 13314 427 13348 461
rect 13348 427 13354 461
rect 13302 418 13354 427
rect 13372 461 13424 470
rect 13372 427 13387 461
rect 13387 427 13421 461
rect 13421 427 13424 461
rect 13372 418 13424 427
rect 13442 461 13494 470
rect 13442 427 13460 461
rect 13460 427 13494 461
rect 13442 418 13494 427
rect 13511 461 13563 470
rect 13580 461 13632 470
rect 13649 461 13701 470
rect 13718 461 13770 470
rect 13787 461 13839 470
rect 13856 461 13908 470
rect 13925 461 13977 470
rect 13511 427 13533 461
rect 13533 427 13563 461
rect 13580 427 13606 461
rect 13606 427 13632 461
rect 13649 427 13679 461
rect 13679 427 13701 461
rect 13718 427 13752 461
rect 13752 427 13770 461
rect 13787 427 13825 461
rect 13825 427 13839 461
rect 13856 427 13859 461
rect 13859 427 13898 461
rect 13898 427 13908 461
rect 13925 427 13932 461
rect 13932 427 13971 461
rect 13971 427 13977 461
rect 13511 418 13563 427
rect 13580 418 13632 427
rect 13649 418 13701 427
rect 13718 418 13770 427
rect 13787 418 13839 427
rect 13856 418 13908 427
rect 13925 418 13977 427
rect 15005 341 15057 393
rect 15069 341 15121 393
rect 473 230 525 239
rect 473 196 478 230
rect 478 196 512 230
rect 512 196 525 230
rect 473 187 525 196
rect 537 230 589 239
rect 537 196 550 230
rect 550 196 584 230
rect 584 196 589 230
rect 537 187 589 196
rect 3209 187 3261 239
rect 3273 187 3325 239
rect 5149 187 5201 239
rect 5213 187 5265 239
rect 10789 187 10841 239
rect 10853 187 10905 239
rect 15173 187 15225 239
rect 15237 187 15289 239
rect 363 84 415 93
rect 427 84 479 93
rect 491 84 543 93
rect 555 84 607 93
rect 619 84 671 93
rect 683 84 735 93
rect 363 50 389 84
rect 389 50 415 84
rect 427 50 461 84
rect 461 50 479 84
rect 491 50 495 84
rect 495 50 533 84
rect 533 50 543 84
rect 555 50 567 84
rect 567 50 605 84
rect 605 50 607 84
rect 619 50 639 84
rect 639 50 671 84
rect 683 50 711 84
rect 711 50 735 84
rect 363 41 415 50
rect 427 41 479 50
rect 491 41 543 50
rect 555 41 607 50
rect 619 41 671 50
rect 683 41 735 50
rect 886 84 938 93
rect 950 84 1002 93
rect 1014 84 1066 93
rect 1078 84 1130 93
rect 1142 84 1194 93
rect 1206 84 1258 93
rect 886 50 915 84
rect 915 50 938 84
rect 950 50 987 84
rect 987 50 1002 84
rect 1014 50 1021 84
rect 1021 50 1059 84
rect 1059 50 1066 84
rect 1078 50 1093 84
rect 1093 50 1130 84
rect 1142 50 1165 84
rect 1165 50 1194 84
rect 1206 50 1237 84
rect 1237 50 1258 84
rect 886 41 938 50
rect 950 41 1002 50
rect 1014 41 1066 50
rect 1078 41 1130 50
rect 1142 41 1194 50
rect 1206 41 1258 50
rect 1270 84 1322 93
rect 1270 50 1275 84
rect 1275 50 1309 84
rect 1309 50 1322 84
rect 1270 41 1322 50
rect 1334 84 1386 93
rect 1334 50 1347 84
rect 1347 50 1381 84
rect 1381 50 1386 84
rect 1334 41 1386 50
rect 1398 84 1450 93
rect 1462 84 1514 93
rect 1526 84 1578 93
rect 1590 84 1642 93
rect 1654 84 1706 93
rect 1718 84 1770 93
rect 1782 84 1834 93
rect 1398 50 1419 84
rect 1419 50 1450 84
rect 1462 50 1491 84
rect 1491 50 1514 84
rect 1526 50 1563 84
rect 1563 50 1578 84
rect 1590 50 1597 84
rect 1597 50 1635 84
rect 1635 50 1642 84
rect 1654 50 1669 84
rect 1669 50 1706 84
rect 1718 50 1741 84
rect 1741 50 1770 84
rect 1782 50 1813 84
rect 1813 50 1834 84
rect 1398 41 1450 50
rect 1462 41 1514 50
rect 1526 41 1578 50
rect 1590 41 1642 50
rect 1654 41 1706 50
rect 1718 41 1770 50
rect 1782 41 1834 50
rect 1846 84 1898 93
rect 1846 50 1851 84
rect 1851 50 1885 84
rect 1885 50 1898 84
rect 1846 41 1898 50
rect 1910 84 1962 93
rect 1910 50 1923 84
rect 1923 50 1957 84
rect 1957 50 1962 84
rect 1910 41 1962 50
rect 1974 84 2026 93
rect 2038 84 2090 93
rect 2102 84 2154 93
rect 2166 84 2218 93
rect 2230 84 2282 93
rect 2294 84 2346 93
rect 2358 84 2410 93
rect 1974 50 1995 84
rect 1995 50 2026 84
rect 2038 50 2067 84
rect 2067 50 2090 84
rect 2102 50 2139 84
rect 2139 50 2154 84
rect 2166 50 2173 84
rect 2173 50 2211 84
rect 2211 50 2218 84
rect 2230 50 2245 84
rect 2245 50 2282 84
rect 2294 50 2317 84
rect 2317 50 2346 84
rect 2358 50 2389 84
rect 2389 50 2410 84
rect 1974 41 2026 50
rect 2038 41 2090 50
rect 2102 41 2154 50
rect 2166 41 2218 50
rect 2230 41 2282 50
rect 2294 41 2346 50
rect 2358 41 2410 50
rect 2422 84 2474 93
rect 2422 50 2427 84
rect 2427 50 2461 84
rect 2461 50 2474 84
rect 2422 41 2474 50
rect 2486 84 2538 93
rect 2486 50 2499 84
rect 2499 50 2533 84
rect 2533 50 2538 84
rect 2486 41 2538 50
rect 2550 84 2602 93
rect 2614 84 2666 93
rect 2678 84 2730 93
rect 2742 84 2794 93
rect 2806 84 2858 93
rect 2870 84 2922 93
rect 2934 84 2986 93
rect 2550 50 2571 84
rect 2571 50 2602 84
rect 2614 50 2643 84
rect 2643 50 2666 84
rect 2678 50 2715 84
rect 2715 50 2730 84
rect 2742 50 2749 84
rect 2749 50 2787 84
rect 2787 50 2794 84
rect 2806 50 2821 84
rect 2821 50 2858 84
rect 2870 50 2893 84
rect 2893 50 2922 84
rect 2934 50 2965 84
rect 2965 50 2986 84
rect 2550 41 2602 50
rect 2614 41 2666 50
rect 2678 41 2730 50
rect 2742 41 2794 50
rect 2806 41 2858 50
rect 2870 41 2922 50
rect 2934 41 2986 50
rect 2998 84 3050 93
rect 2998 50 3003 84
rect 3003 50 3037 84
rect 3037 50 3050 84
rect 2998 41 3050 50
rect 3062 84 3114 93
rect 3062 50 3075 84
rect 3075 50 3109 84
rect 3109 50 3114 84
rect 3062 41 3114 50
rect 3126 84 3178 93
rect 3190 84 3242 93
rect 3254 84 3306 93
rect 3318 84 3370 93
rect 3382 84 3434 93
rect 3446 84 3498 93
rect 3510 84 3562 93
rect 3126 50 3147 84
rect 3147 50 3178 84
rect 3190 50 3219 84
rect 3219 50 3242 84
rect 3254 50 3291 84
rect 3291 50 3306 84
rect 3318 50 3325 84
rect 3325 50 3363 84
rect 3363 50 3370 84
rect 3382 50 3397 84
rect 3397 50 3434 84
rect 3446 50 3469 84
rect 3469 50 3498 84
rect 3510 50 3541 84
rect 3541 50 3562 84
rect 3126 41 3178 50
rect 3190 41 3242 50
rect 3254 41 3306 50
rect 3318 41 3370 50
rect 3382 41 3434 50
rect 3446 41 3498 50
rect 3510 41 3562 50
rect 3574 84 3626 93
rect 3574 50 3579 84
rect 3579 50 3613 84
rect 3613 50 3626 84
rect 3574 41 3626 50
rect 3638 84 3690 93
rect 3638 50 3651 84
rect 3651 50 3685 84
rect 3685 50 3690 84
rect 3638 41 3690 50
rect 3702 84 3754 93
rect 3766 84 3818 93
rect 3830 84 3882 93
rect 3894 84 3946 93
rect 3958 84 4010 93
rect 4022 84 4074 93
rect 4086 84 4138 93
rect 3702 50 3723 84
rect 3723 50 3754 84
rect 3766 50 3795 84
rect 3795 50 3818 84
rect 3830 50 3867 84
rect 3867 50 3882 84
rect 3894 50 3901 84
rect 3901 50 3939 84
rect 3939 50 3946 84
rect 3958 50 3973 84
rect 3973 50 4010 84
rect 4022 50 4045 84
rect 4045 50 4074 84
rect 4086 50 4117 84
rect 4117 50 4138 84
rect 3702 41 3754 50
rect 3766 41 3818 50
rect 3830 41 3882 50
rect 3894 41 3946 50
rect 3958 41 4010 50
rect 4022 41 4074 50
rect 4086 41 4138 50
rect 4150 84 4202 93
rect 4150 50 4155 84
rect 4155 50 4189 84
rect 4189 50 4202 84
rect 4150 41 4202 50
rect 4214 84 4266 93
rect 4214 50 4227 84
rect 4227 50 4261 84
rect 4261 50 4266 84
rect 4214 41 4266 50
rect 4278 84 4330 93
rect 4342 84 4394 93
rect 4406 84 4458 93
rect 4470 84 4522 93
rect 4534 84 4586 93
rect 4598 84 4650 93
rect 4662 84 4714 93
rect 4278 50 4299 84
rect 4299 50 4330 84
rect 4342 50 4371 84
rect 4371 50 4394 84
rect 4406 50 4443 84
rect 4443 50 4458 84
rect 4470 50 4477 84
rect 4477 50 4515 84
rect 4515 50 4522 84
rect 4534 50 4549 84
rect 4549 50 4586 84
rect 4598 50 4621 84
rect 4621 50 4650 84
rect 4662 50 4693 84
rect 4693 50 4714 84
rect 4278 41 4330 50
rect 4342 41 4394 50
rect 4406 41 4458 50
rect 4470 41 4522 50
rect 4534 41 4586 50
rect 4598 41 4650 50
rect 4662 41 4714 50
rect 4726 84 4778 93
rect 4726 50 4731 84
rect 4731 50 4765 84
rect 4765 50 4778 84
rect 4726 41 4778 50
rect 4790 84 4842 93
rect 4790 50 4803 84
rect 4803 50 4837 84
rect 4837 50 4842 84
rect 4790 41 4842 50
rect 4854 84 4906 93
rect 4918 84 4970 93
rect 4982 84 5034 93
rect 5046 84 5098 93
rect 5110 84 5162 93
rect 5174 84 5226 93
rect 5238 84 5290 93
rect 4854 50 4875 84
rect 4875 50 4906 84
rect 4918 50 4947 84
rect 4947 50 4970 84
rect 4982 50 5019 84
rect 5019 50 5034 84
rect 5046 50 5053 84
rect 5053 50 5091 84
rect 5091 50 5098 84
rect 5110 50 5125 84
rect 5125 50 5162 84
rect 5174 50 5197 84
rect 5197 50 5226 84
rect 5238 50 5269 84
rect 5269 50 5290 84
rect 4854 41 4906 50
rect 4918 41 4970 50
rect 4982 41 5034 50
rect 5046 41 5098 50
rect 5110 41 5162 50
rect 5174 41 5226 50
rect 5238 41 5290 50
rect 5302 84 5354 93
rect 5302 50 5307 84
rect 5307 50 5341 84
rect 5341 50 5354 84
rect 5302 41 5354 50
rect 5366 84 5418 93
rect 5366 50 5379 84
rect 5379 50 5413 84
rect 5413 50 5418 84
rect 5366 41 5418 50
rect 5430 84 5482 93
rect 5494 84 5546 93
rect 5558 84 5610 93
rect 5622 84 5674 93
rect 5686 84 5738 93
rect 5750 84 5802 93
rect 5814 84 5866 93
rect 5430 50 5451 84
rect 5451 50 5482 84
rect 5494 50 5523 84
rect 5523 50 5546 84
rect 5558 50 5595 84
rect 5595 50 5610 84
rect 5622 50 5629 84
rect 5629 50 5667 84
rect 5667 50 5674 84
rect 5686 50 5701 84
rect 5701 50 5738 84
rect 5750 50 5773 84
rect 5773 50 5802 84
rect 5814 50 5845 84
rect 5845 50 5866 84
rect 5430 41 5482 50
rect 5494 41 5546 50
rect 5558 41 5610 50
rect 5622 41 5674 50
rect 5686 41 5738 50
rect 5750 41 5802 50
rect 5814 41 5866 50
rect 5878 84 5930 93
rect 5878 50 5883 84
rect 5883 50 5917 84
rect 5917 50 5930 84
rect 5878 41 5930 50
rect 5942 84 5994 93
rect 5942 50 5955 84
rect 5955 50 5989 84
rect 5989 50 5994 84
rect 5942 41 5994 50
rect 6006 84 6058 93
rect 6070 84 6122 93
rect 6134 84 6186 93
rect 6198 84 6250 93
rect 6262 84 6314 93
rect 6326 84 6378 93
rect 6390 84 6442 93
rect 6006 50 6027 84
rect 6027 50 6058 84
rect 6070 50 6099 84
rect 6099 50 6122 84
rect 6134 50 6171 84
rect 6171 50 6186 84
rect 6198 50 6205 84
rect 6205 50 6243 84
rect 6243 50 6250 84
rect 6262 50 6277 84
rect 6277 50 6314 84
rect 6326 50 6349 84
rect 6349 50 6378 84
rect 6390 50 6421 84
rect 6421 50 6442 84
rect 6006 41 6058 50
rect 6070 41 6122 50
rect 6134 41 6186 50
rect 6198 41 6250 50
rect 6262 41 6314 50
rect 6326 41 6378 50
rect 6390 41 6442 50
rect 6454 84 6506 93
rect 6454 50 6459 84
rect 6459 50 6493 84
rect 6493 50 6506 84
rect 6454 41 6506 50
rect 6518 84 6570 93
rect 6518 50 6531 84
rect 6531 50 6565 84
rect 6565 50 6570 84
rect 6518 41 6570 50
rect 6582 84 6634 93
rect 6646 84 6698 93
rect 6710 84 6762 93
rect 6774 84 6826 93
rect 6838 84 6890 93
rect 6902 84 6954 93
rect 6966 84 7018 93
rect 6582 50 6603 84
rect 6603 50 6634 84
rect 6646 50 6675 84
rect 6675 50 6698 84
rect 6710 50 6747 84
rect 6747 50 6762 84
rect 6774 50 6781 84
rect 6781 50 6819 84
rect 6819 50 6826 84
rect 6838 50 6853 84
rect 6853 50 6890 84
rect 6902 50 6925 84
rect 6925 50 6954 84
rect 6966 50 6997 84
rect 6997 50 7018 84
rect 6582 41 6634 50
rect 6646 41 6698 50
rect 6710 41 6762 50
rect 6774 41 6826 50
rect 6838 41 6890 50
rect 6902 41 6954 50
rect 6966 41 7018 50
rect 7030 84 7082 93
rect 7030 50 7035 84
rect 7035 50 7069 84
rect 7069 50 7082 84
rect 7030 41 7082 50
rect 7094 84 7146 93
rect 7094 50 7107 84
rect 7107 50 7141 84
rect 7141 50 7146 84
rect 7094 41 7146 50
rect 7158 84 7210 93
rect 7222 84 7274 93
rect 7286 84 7338 93
rect 7350 84 7402 93
rect 7414 84 7466 93
rect 7478 84 7530 93
rect 7542 84 7594 93
rect 7158 50 7179 84
rect 7179 50 7210 84
rect 7222 50 7251 84
rect 7251 50 7274 84
rect 7286 50 7323 84
rect 7323 50 7338 84
rect 7350 50 7357 84
rect 7357 50 7395 84
rect 7395 50 7402 84
rect 7414 50 7429 84
rect 7429 50 7466 84
rect 7478 50 7501 84
rect 7501 50 7530 84
rect 7542 50 7573 84
rect 7573 50 7594 84
rect 7158 41 7210 50
rect 7222 41 7274 50
rect 7286 41 7338 50
rect 7350 41 7402 50
rect 7414 41 7466 50
rect 7478 41 7530 50
rect 7542 41 7594 50
rect 7606 84 7658 93
rect 7606 50 7611 84
rect 7611 50 7645 84
rect 7645 50 7658 84
rect 7606 41 7658 50
rect 7670 84 7722 93
rect 7670 50 7683 84
rect 7683 50 7717 84
rect 7717 50 7722 84
rect 7670 41 7722 50
rect 7734 84 7786 93
rect 7798 84 7850 93
rect 7862 84 7914 93
rect 7926 84 7978 93
rect 7990 84 8042 93
rect 8054 84 8106 93
rect 8118 84 8170 93
rect 7734 50 7755 84
rect 7755 50 7786 84
rect 7798 50 7827 84
rect 7827 50 7850 84
rect 7862 50 7899 84
rect 7899 50 7914 84
rect 7926 50 7933 84
rect 7933 50 7971 84
rect 7971 50 7978 84
rect 7990 50 8005 84
rect 8005 50 8042 84
rect 8054 50 8077 84
rect 8077 50 8106 84
rect 8118 50 8149 84
rect 8149 50 8170 84
rect 7734 41 7786 50
rect 7798 41 7850 50
rect 7862 41 7914 50
rect 7926 41 7978 50
rect 7990 41 8042 50
rect 8054 41 8106 50
rect 8118 41 8170 50
rect 8182 84 8234 93
rect 8182 50 8187 84
rect 8187 50 8221 84
rect 8221 50 8234 84
rect 8182 41 8234 50
rect 8246 84 8298 93
rect 8246 50 8259 84
rect 8259 50 8293 84
rect 8293 50 8298 84
rect 8246 41 8298 50
rect 8310 84 8362 93
rect 8374 84 8426 93
rect 8438 84 8490 93
rect 8502 84 8554 93
rect 8566 84 8618 93
rect 8630 84 8682 93
rect 8694 84 8746 93
rect 8310 50 8331 84
rect 8331 50 8362 84
rect 8374 50 8403 84
rect 8403 50 8426 84
rect 8438 50 8475 84
rect 8475 50 8490 84
rect 8502 50 8509 84
rect 8509 50 8547 84
rect 8547 50 8554 84
rect 8566 50 8581 84
rect 8581 50 8618 84
rect 8630 50 8653 84
rect 8653 50 8682 84
rect 8694 50 8725 84
rect 8725 50 8746 84
rect 8310 41 8362 50
rect 8374 41 8426 50
rect 8438 41 8490 50
rect 8502 41 8554 50
rect 8566 41 8618 50
rect 8630 41 8682 50
rect 8694 41 8746 50
rect 8758 84 8810 93
rect 8758 50 8763 84
rect 8763 50 8797 84
rect 8797 50 8810 84
rect 8758 41 8810 50
rect 8822 84 8874 93
rect 8822 50 8835 84
rect 8835 50 8869 84
rect 8869 50 8874 84
rect 8822 41 8874 50
rect 8886 84 8938 93
rect 8950 84 9002 93
rect 9014 84 9066 93
rect 9078 84 9130 93
rect 9142 84 9194 93
rect 9206 84 9258 93
rect 9270 84 9322 93
rect 8886 50 8907 84
rect 8907 50 8938 84
rect 8950 50 8979 84
rect 8979 50 9002 84
rect 9014 50 9051 84
rect 9051 50 9066 84
rect 9078 50 9085 84
rect 9085 50 9123 84
rect 9123 50 9130 84
rect 9142 50 9157 84
rect 9157 50 9194 84
rect 9206 50 9229 84
rect 9229 50 9258 84
rect 9270 50 9301 84
rect 9301 50 9322 84
rect 8886 41 8938 50
rect 8950 41 9002 50
rect 9014 41 9066 50
rect 9078 41 9130 50
rect 9142 41 9194 50
rect 9206 41 9258 50
rect 9270 41 9322 50
rect 9334 84 9386 93
rect 9334 50 9339 84
rect 9339 50 9373 84
rect 9373 50 9386 84
rect 9334 41 9386 50
rect 9398 84 9450 93
rect 9398 50 9411 84
rect 9411 50 9445 84
rect 9445 50 9450 84
rect 9398 41 9450 50
rect 9462 84 9514 93
rect 9526 84 9578 93
rect 9590 84 9642 93
rect 9654 84 9706 93
rect 9718 84 9770 93
rect 9782 84 9834 93
rect 9846 84 9898 93
rect 9462 50 9483 84
rect 9483 50 9514 84
rect 9526 50 9555 84
rect 9555 50 9578 84
rect 9590 50 9627 84
rect 9627 50 9642 84
rect 9654 50 9661 84
rect 9661 50 9699 84
rect 9699 50 9706 84
rect 9718 50 9733 84
rect 9733 50 9770 84
rect 9782 50 9805 84
rect 9805 50 9834 84
rect 9846 50 9877 84
rect 9877 50 9898 84
rect 9462 41 9514 50
rect 9526 41 9578 50
rect 9590 41 9642 50
rect 9654 41 9706 50
rect 9718 41 9770 50
rect 9782 41 9834 50
rect 9846 41 9898 50
rect 9910 84 9962 93
rect 9910 50 9915 84
rect 9915 50 9949 84
rect 9949 50 9962 84
rect 9910 41 9962 50
rect 9974 84 10026 93
rect 9974 50 9987 84
rect 9987 50 10021 84
rect 10021 50 10026 84
rect 9974 41 10026 50
rect 10038 84 10090 93
rect 10102 84 10154 93
rect 10166 84 10218 93
rect 10230 84 10282 93
rect 10294 84 10346 93
rect 10358 84 10410 93
rect 10422 84 10474 93
rect 10038 50 10059 84
rect 10059 50 10090 84
rect 10102 50 10131 84
rect 10131 50 10154 84
rect 10166 50 10203 84
rect 10203 50 10218 84
rect 10230 50 10237 84
rect 10237 50 10275 84
rect 10275 50 10282 84
rect 10294 50 10309 84
rect 10309 50 10346 84
rect 10358 50 10381 84
rect 10381 50 10410 84
rect 10422 50 10453 84
rect 10453 50 10474 84
rect 10038 41 10090 50
rect 10102 41 10154 50
rect 10166 41 10218 50
rect 10230 41 10282 50
rect 10294 41 10346 50
rect 10358 41 10410 50
rect 10422 41 10474 50
rect 10486 84 10538 93
rect 10486 50 10491 84
rect 10491 50 10525 84
rect 10525 50 10538 84
rect 10486 41 10538 50
rect 10550 84 10602 93
rect 10550 50 10563 84
rect 10563 50 10597 84
rect 10597 50 10602 84
rect 10550 41 10602 50
rect 10614 84 10666 93
rect 10678 84 10730 93
rect 10742 84 10794 93
rect 10806 84 10858 93
rect 10870 84 10922 93
rect 10934 84 10986 93
rect 10998 84 11050 93
rect 10614 50 10635 84
rect 10635 50 10666 84
rect 10678 50 10707 84
rect 10707 50 10730 84
rect 10742 50 10779 84
rect 10779 50 10794 84
rect 10806 50 10813 84
rect 10813 50 10851 84
rect 10851 50 10858 84
rect 10870 50 10885 84
rect 10885 50 10922 84
rect 10934 50 10957 84
rect 10957 50 10986 84
rect 10998 50 11029 84
rect 11029 50 11050 84
rect 10614 41 10666 50
rect 10678 41 10730 50
rect 10742 41 10794 50
rect 10806 41 10858 50
rect 10870 41 10922 50
rect 10934 41 10986 50
rect 10998 41 11050 50
rect 11062 84 11114 93
rect 11062 50 11067 84
rect 11067 50 11101 84
rect 11101 50 11114 84
rect 11062 41 11114 50
rect 11126 84 11178 93
rect 11126 50 11139 84
rect 11139 50 11173 84
rect 11173 50 11178 84
rect 11126 41 11178 50
rect 11190 84 11242 93
rect 11254 84 11306 93
rect 11318 84 11370 93
rect 11382 84 11434 93
rect 11446 84 11498 93
rect 11510 84 11562 93
rect 11574 84 11626 93
rect 11190 50 11211 84
rect 11211 50 11242 84
rect 11254 50 11283 84
rect 11283 50 11306 84
rect 11318 50 11355 84
rect 11355 50 11370 84
rect 11382 50 11389 84
rect 11389 50 11427 84
rect 11427 50 11434 84
rect 11446 50 11461 84
rect 11461 50 11498 84
rect 11510 50 11533 84
rect 11533 50 11562 84
rect 11574 50 11605 84
rect 11605 50 11626 84
rect 11190 41 11242 50
rect 11254 41 11306 50
rect 11318 41 11370 50
rect 11382 41 11434 50
rect 11446 41 11498 50
rect 11510 41 11562 50
rect 11574 41 11626 50
rect 11638 84 11690 93
rect 11638 50 11643 84
rect 11643 50 11677 84
rect 11677 50 11690 84
rect 11638 41 11690 50
rect 11702 84 11754 93
rect 11702 50 11715 84
rect 11715 50 11749 84
rect 11749 50 11754 84
rect 11702 41 11754 50
rect 11766 84 11818 93
rect 11830 84 11882 93
rect 11894 84 11946 93
rect 11958 84 12010 93
rect 12022 84 12074 93
rect 12086 84 12138 93
rect 12150 84 12202 93
rect 11766 50 11787 84
rect 11787 50 11818 84
rect 11830 50 11859 84
rect 11859 50 11882 84
rect 11894 50 11931 84
rect 11931 50 11946 84
rect 11958 50 11965 84
rect 11965 50 12003 84
rect 12003 50 12010 84
rect 12022 50 12037 84
rect 12037 50 12074 84
rect 12086 50 12109 84
rect 12109 50 12138 84
rect 12150 50 12181 84
rect 12181 50 12202 84
rect 11766 41 11818 50
rect 11830 41 11882 50
rect 11894 41 11946 50
rect 11958 41 12010 50
rect 12022 41 12074 50
rect 12086 41 12138 50
rect 12150 41 12202 50
rect 12214 84 12266 93
rect 12214 50 12219 84
rect 12219 50 12253 84
rect 12253 50 12266 84
rect 12214 41 12266 50
rect 12278 84 12330 93
rect 12278 50 12291 84
rect 12291 50 12325 84
rect 12325 50 12330 84
rect 12278 41 12330 50
rect 12342 84 12394 93
rect 12406 84 12458 93
rect 12470 84 12522 93
rect 12534 84 12586 93
rect 12598 84 12650 93
rect 12662 84 12714 93
rect 12726 84 12778 93
rect 12342 50 12363 84
rect 12363 50 12394 84
rect 12406 50 12435 84
rect 12435 50 12458 84
rect 12470 50 12507 84
rect 12507 50 12522 84
rect 12534 50 12541 84
rect 12541 50 12579 84
rect 12579 50 12586 84
rect 12598 50 12613 84
rect 12613 50 12650 84
rect 12662 50 12685 84
rect 12685 50 12714 84
rect 12726 50 12757 84
rect 12757 50 12778 84
rect 12342 41 12394 50
rect 12406 41 12458 50
rect 12470 41 12522 50
rect 12534 41 12586 50
rect 12598 41 12650 50
rect 12662 41 12714 50
rect 12726 41 12778 50
rect 12790 84 12842 93
rect 12790 50 12795 84
rect 12795 50 12829 84
rect 12829 50 12842 84
rect 12790 41 12842 50
rect 12854 84 12906 93
rect 12854 50 12867 84
rect 12867 50 12901 84
rect 12901 50 12906 84
rect 12854 41 12906 50
rect 12918 84 12970 93
rect 12982 84 13034 93
rect 13046 84 13098 93
rect 13110 84 13162 93
rect 13174 84 13226 93
rect 13238 84 13290 93
rect 13302 84 13354 93
rect 12918 50 12939 84
rect 12939 50 12970 84
rect 12982 50 13011 84
rect 13011 50 13034 84
rect 13046 50 13083 84
rect 13083 50 13098 84
rect 13110 50 13117 84
rect 13117 50 13155 84
rect 13155 50 13162 84
rect 13174 50 13189 84
rect 13189 50 13226 84
rect 13238 50 13261 84
rect 13261 50 13290 84
rect 13302 50 13333 84
rect 13333 50 13354 84
rect 12918 41 12970 50
rect 12982 41 13034 50
rect 13046 41 13098 50
rect 13110 41 13162 50
rect 13174 41 13226 50
rect 13238 41 13290 50
rect 13302 41 13354 50
rect 13366 84 13418 93
rect 13366 50 13371 84
rect 13371 50 13405 84
rect 13405 50 13418 84
rect 13366 41 13418 50
rect 13430 84 13482 93
rect 13430 50 13443 84
rect 13443 50 13477 84
rect 13477 50 13482 84
rect 13430 41 13482 50
rect 13494 84 13546 93
rect 13558 84 13610 93
rect 13622 84 13674 93
rect 13686 84 13738 93
rect 13750 84 13802 93
rect 13814 84 13866 93
rect 13878 84 13930 93
rect 13494 50 13515 84
rect 13515 50 13546 84
rect 13558 50 13587 84
rect 13587 50 13610 84
rect 13622 50 13659 84
rect 13659 50 13674 84
rect 13686 50 13693 84
rect 13693 50 13731 84
rect 13731 50 13738 84
rect 13750 50 13765 84
rect 13765 50 13802 84
rect 13814 50 13837 84
rect 13837 50 13866 84
rect 13878 50 13909 84
rect 13909 50 13930 84
rect 13494 41 13546 50
rect 13558 41 13610 50
rect 13622 41 13674 50
rect 13686 41 13738 50
rect 13750 41 13802 50
rect 13814 41 13866 50
rect 13878 41 13930 50
rect 13942 84 13994 93
rect 13942 50 13947 84
rect 13947 50 13981 84
rect 13981 50 13994 84
rect 13942 41 13994 50
rect 14006 84 14058 93
rect 14006 50 14019 84
rect 14019 50 14053 84
rect 14053 50 14058 84
rect 14006 41 14058 50
rect 14070 84 14122 93
rect 14134 84 14186 93
rect 14198 84 14250 93
rect 14262 84 14314 93
rect 14326 84 14378 93
rect 14070 50 14091 84
rect 14091 50 14122 84
rect 14134 50 14163 84
rect 14163 50 14186 84
rect 14198 50 14235 84
rect 14235 50 14250 84
rect 14262 50 14269 84
rect 14269 50 14307 84
rect 14307 50 14314 84
rect 14326 50 14341 84
rect 14341 50 14378 84
rect 14070 41 14122 50
rect 14134 41 14186 50
rect 14198 41 14250 50
rect 14262 41 14314 50
rect 14326 41 14378 50
<< metal2 >>
rect 348 7975 354 8027
rect 406 7975 418 8027
rect 470 7975 482 8027
rect 534 7975 546 8027
rect 598 7975 610 8027
rect 662 7975 674 8027
rect 726 7975 857 8027
rect 909 7975 921 8027
rect 973 7975 985 8027
rect 1037 7975 1049 8027
rect 1101 7975 1113 8027
rect 1165 7975 1177 8027
rect 1229 7975 1241 8027
rect 1293 7975 1305 8027
rect 1357 7975 1369 8027
rect 1421 7975 1433 8027
rect 1485 7975 1497 8027
rect 1549 7975 1561 8027
rect 1613 7975 1625 8027
rect 1677 7975 1689 8027
rect 1741 7975 1753 8027
rect 1805 7975 1817 8027
rect 1869 7975 1881 8027
rect 1933 7975 1945 8027
rect 1997 7975 2009 8027
rect 2061 7975 2073 8027
rect 2125 7975 2137 8027
rect 2189 7975 2201 8027
rect 2253 7975 2265 8027
rect 2317 7975 2329 8027
rect 2381 7975 2393 8027
rect 2445 7975 2457 8027
rect 2509 7975 2521 8027
rect 2573 7975 2585 8027
rect 2637 7975 2649 8027
rect 2701 7975 2713 8027
rect 2765 7975 2777 8027
rect 2829 7975 2841 8027
rect 2893 7975 2905 8027
rect 2957 7975 2969 8027
rect 3021 7975 3033 8027
rect 3085 7975 3097 8027
rect 3149 7975 3161 8027
rect 3213 7975 3225 8027
rect 3277 7975 3289 8027
rect 3341 7975 3353 8027
rect 3405 7975 3417 8027
rect 3469 7975 3481 8027
rect 3533 7975 3545 8027
rect 3597 7975 3609 8027
rect 3661 7975 3673 8027
rect 3725 7975 3737 8027
rect 3789 7975 3801 8027
rect 3853 7975 3865 8027
rect 3917 7975 3929 8027
rect 3981 7975 3993 8027
rect 4045 7975 4057 8027
rect 4109 7975 4121 8027
rect 4173 7975 4185 8027
rect 4237 7975 4249 8027
rect 4301 7975 4313 8027
rect 4365 7975 4377 8027
rect 4429 7975 4441 8027
rect 4493 7975 4505 8027
rect 4557 7975 4722 8027
rect 4774 7975 4786 8027
rect 4838 7975 4850 8027
rect 4902 7975 4914 8027
rect 4966 7975 4978 8027
rect 5030 7975 5042 8027
rect 5094 7975 5106 8027
rect 5158 7975 5170 8027
rect 5222 7975 5234 8027
rect 5286 7975 5298 8027
rect 5350 7975 5362 8027
rect 5414 7975 5426 8027
rect 5478 7975 5490 8027
rect 5542 7975 5554 8027
rect 5606 7975 5618 8027
rect 5670 7975 5682 8027
rect 5734 7975 5746 8027
rect 5798 7975 5810 8027
rect 5862 7975 5874 8027
rect 5926 7975 5938 8027
rect 5990 7975 6002 8027
rect 6054 7975 6066 8027
rect 6118 7975 6130 8027
rect 6182 7975 6194 8027
rect 6246 7975 6258 8027
rect 6310 7975 6322 8027
rect 6374 7975 6386 8027
rect 6438 7975 6450 8027
rect 6502 7975 6514 8027
rect 6566 7975 6578 8027
rect 6630 7975 6810 8027
rect 6862 7975 6874 8027
rect 6926 7975 6938 8027
rect 6990 7975 7002 8027
rect 7054 7975 7066 8027
rect 7118 7975 7130 8027
rect 7182 7975 7194 8027
rect 7246 7975 7258 8027
rect 7310 7975 7322 8027
rect 7374 7975 7386 8027
rect 7438 7975 7450 8027
rect 7502 7975 7514 8027
rect 7566 7975 7578 8027
rect 7630 7975 7642 8027
rect 7694 7975 7706 8027
rect 7758 7975 7770 8027
rect 7822 7975 7834 8027
rect 7886 7975 7898 8027
rect 7950 7975 7962 8027
rect 8014 7975 8026 8027
rect 8078 7975 8090 8027
rect 8142 7975 8154 8027
rect 8206 7975 8218 8027
rect 8270 7975 8282 8027
rect 8334 7975 8346 8027
rect 8398 7975 8410 8027
rect 8462 7975 8474 8027
rect 8526 7975 8538 8027
rect 8590 7975 8602 8027
rect 8654 7975 8666 8027
rect 8718 7975 8730 8027
rect 8782 7975 8794 8027
rect 8846 7975 8858 8027
rect 8910 7975 8922 8027
rect 8974 7975 8986 8027
rect 9038 7975 9050 8027
rect 9102 7975 9114 8027
rect 9166 7975 9178 8027
rect 9230 7975 9242 8027
rect 9294 7975 9306 8027
rect 9358 7975 9370 8027
rect 9422 7975 9434 8027
rect 9486 7975 9498 8027
rect 9550 7975 9562 8027
rect 9614 7975 9626 8027
rect 9678 7975 9690 8027
rect 9742 7975 9754 8027
rect 9806 7975 9818 8027
rect 9870 7975 9882 8027
rect 9934 7975 9946 8027
rect 9998 7975 10010 8027
rect 10062 7975 10074 8027
rect 10126 7975 10138 8027
rect 10190 7975 10202 8027
rect 10254 7975 10266 8027
rect 10318 7975 10330 8027
rect 10382 7975 10394 8027
rect 10446 7975 10458 8027
rect 10510 7975 10522 8027
rect 10574 7975 10586 8027
rect 10638 7975 10650 8027
rect 10702 7975 10714 8027
rect 10766 7975 10778 8027
rect 10830 7975 10842 8027
rect 10894 7975 10906 8027
rect 10958 7975 10970 8027
rect 11022 7975 11034 8027
rect 11086 7975 11098 8027
rect 11150 7975 11162 8027
rect 11214 7975 11226 8027
rect 11278 7975 11290 8027
rect 11342 7975 11354 8027
rect 11406 7975 11418 8027
rect 11470 7975 11482 8027
rect 11534 7975 11546 8027
rect 11598 7975 11610 8027
rect 11662 7975 11674 8027
rect 11726 7975 11738 8027
rect 11790 7975 11802 8027
rect 11854 7975 11866 8027
rect 11918 7975 11930 8027
rect 11982 7975 11994 8027
rect 12046 7975 12058 8027
rect 12110 7975 12122 8027
rect 12174 7975 12186 8027
rect 12238 7975 12250 8027
rect 12302 7975 12314 8027
rect 12366 7975 12378 8027
rect 12430 7975 12442 8027
rect 12494 7975 12506 8027
rect 12558 7975 12570 8027
rect 12622 7975 12634 8027
rect 12686 7975 12698 8027
rect 12750 7975 12762 8027
rect 12814 7975 12826 8027
rect 12878 7975 12890 8027
rect 12942 7975 12954 8027
rect 13006 7975 13018 8027
rect 13070 7975 13082 8027
rect 13134 7975 13146 8027
rect 13198 7975 13210 8027
rect 13262 7975 13274 8027
rect 13326 7975 13338 8027
rect 13390 7975 13402 8027
rect 13454 7975 13466 8027
rect 13518 7975 13530 8027
rect 13582 7975 13594 8027
rect 13646 7975 16020 8027
rect 467 7830 473 7882
rect 525 7830 537 7882
rect 589 7830 3209 7882
rect 3261 7830 3273 7882
rect 3325 7830 3331 7882
rect 467 7676 473 7728
rect 525 7676 537 7728
rect 589 7676 3213 7728
rect 3265 7676 3277 7728
rect 3329 7676 3335 7728
rect 10279 7676 10285 7728
rect 10337 7676 10349 7728
rect 10401 7708 14963 7728
tri 14963 7708 14983 7728 sw
rect 10401 7676 14983 7708
tri 14941 7634 14983 7676 ne
tri 14983 7634 15057 7708 sw
tri 14983 7574 15043 7634 ne
rect 15043 7574 15057 7634
tri 15057 7574 15117 7634 sw
rect 467 7522 473 7574
rect 525 7522 537 7574
rect 589 7522 3209 7574
rect 3261 7522 3273 7574
rect 3325 7522 3331 7574
tri 15043 7560 15057 7574 ne
rect 15057 7560 15117 7574
tri 15117 7560 15131 7574 sw
tri 15057 7522 15095 7560 ne
rect 15095 7522 15131 7560
tri 15131 7522 15169 7560 sw
tri 15095 7486 15131 7522 ne
rect 15131 7486 15169 7522
tri 15169 7486 15205 7522 sw
tri 15131 7420 15197 7486 ne
rect 15197 7420 15205 7486
tri 15205 7420 15271 7486 sw
rect 467 7368 473 7420
rect 525 7368 537 7420
rect 589 7368 3213 7420
rect 3265 7368 3277 7420
rect 3329 7368 3335 7420
rect 9423 7368 9429 7420
rect 9481 7368 9493 7420
rect 9545 7368 15005 7420
tri 15005 7368 15057 7420 sw
tri 15197 7412 15205 7420 ne
rect 15205 7412 15271 7420
tri 15271 7412 15279 7420 sw
tri 15205 7368 15249 7412 ne
rect 15249 7368 15279 7412
tri 15279 7368 15323 7412 sw
tri 14983 7356 14995 7368 ne
rect 14995 7356 15057 7368
tri 15057 7356 15069 7368 sw
tri 15249 7356 15261 7368 ne
rect 15261 7356 15323 7368
tri 15323 7356 15335 7368 sw
tri 14995 7346 15005 7356 ne
rect 15005 7346 15069 7356
tri 15005 7282 15069 7346 ne
tri 15069 7282 15143 7356 sw
tri 15261 7338 15279 7356 ne
rect 15279 7338 15335 7356
tri 15335 7338 15353 7356 sw
tri 15279 7282 15335 7338 ne
rect 15335 7282 15353 7338
tri 15353 7282 15409 7338 sw
tri 15069 7266 15085 7282 ne
rect 15085 7266 15143 7282
rect 467 7214 473 7266
rect 525 7214 537 7266
rect 589 7214 3209 7266
rect 3261 7214 3273 7266
rect 3325 7214 3331 7266
tri 15085 7214 15137 7266 ne
rect 15137 7214 15143 7266
tri 15137 7208 15143 7214 ne
tri 15143 7208 15217 7282 sw
tri 15335 7264 15353 7282 ne
rect 15353 7264 15409 7282
tri 15409 7264 15427 7282 sw
tri 15353 7208 15409 7264 ne
rect 15409 7208 15427 7264
tri 15427 7208 15483 7264 sw
tri 15143 7134 15217 7208 ne
tri 15217 7134 15291 7208 sw
tri 15409 7190 15427 7208 ne
rect 15427 7190 15483 7208
tri 15483 7190 15501 7208 sw
tri 15427 7134 15483 7190 ne
rect 15483 7134 15501 7190
tri 15501 7134 15557 7190 sw
tri 15217 7112 15239 7134 ne
rect 15239 7112 15291 7134
tri 15291 7112 15313 7134 sw
tri 15483 7116 15501 7134 ne
rect 15501 7116 15557 7134
tri 15557 7116 15575 7134 sw
tri 15501 7112 15505 7116 ne
rect 15505 7112 15575 7116
rect 467 7060 473 7112
rect 525 7060 537 7112
rect 589 7060 3213 7112
rect 3265 7060 3277 7112
rect 3329 7060 3335 7112
rect 8567 7060 8573 7112
rect 8625 7060 8637 7112
rect 8689 7065 15121 7112
tri 15121 7065 15168 7112 sw
tri 15239 7065 15286 7112 ne
rect 15286 7065 15313 7112
tri 15313 7065 15360 7112 sw
tri 15505 7094 15523 7112 ne
rect 8689 7060 15168 7065
tri 15168 7060 15173 7065 sw
tri 15286 7060 15291 7065 ne
rect 15291 7060 15360 7065
tri 15360 7060 15365 7065 sw
tri 15099 6991 15168 7060 ne
rect 15168 6991 15173 7060
tri 15173 6991 15242 7060 sw
tri 15291 6991 15360 7060 ne
rect 15360 6991 15365 7060
tri 15365 6991 15434 7060 sw
tri 15168 6958 15201 6991 ne
rect 15201 6986 15242 6991
tri 15242 6986 15247 6991 sw
tri 15360 6986 15365 6991 ne
rect 15365 6986 15434 6991
tri 15434 6986 15439 6991 sw
rect 15201 6958 15247 6986
rect 467 6906 473 6958
rect 525 6906 537 6958
rect 589 6906 3209 6958
rect 3261 6906 3273 6958
rect 3325 6906 3331 6958
tri 15201 6917 15242 6958 ne
rect 15242 6917 15247 6958
tri 15247 6917 15316 6986 sw
tri 15365 6964 15387 6986 ne
tri 15242 6906 15253 6917 ne
rect 15253 6906 15316 6917
tri 15253 6895 15264 6906 ne
rect 467 6752 473 6804
rect 525 6752 537 6804
rect 589 6752 3213 6804
rect 3265 6752 3277 6804
rect 3329 6752 3335 6804
rect 7711 6752 7717 6804
rect 7769 6752 7781 6804
rect 7833 6800 15105 6804
tri 15105 6800 15109 6804 sw
rect 7833 6752 15109 6800
tri 15083 6726 15109 6752 ne
tri 15109 6726 15183 6800 sw
tri 15109 6704 15131 6726 ne
rect 467 6598 473 6650
rect 525 6598 537 6650
rect 589 6598 3209 6650
rect 3261 6598 3273 6650
rect 3325 6598 3331 6650
rect 467 6444 473 6496
rect 525 6444 537 6496
rect 589 6444 3213 6496
rect 3265 6444 3277 6496
rect 3329 6444 3335 6496
rect 6855 6444 6861 6496
rect 6913 6444 6925 6496
rect 6977 6444 14799 6496
tri 14777 6442 14779 6444 ne
rect 14779 6442 14799 6444
tri 14799 6442 14853 6496 sw
tri 14779 6422 14799 6442 ne
rect 14799 6422 14853 6442
tri 14799 6368 14853 6422 ne
tri 14853 6368 14927 6442 sw
tri 14853 6342 14879 6368 ne
rect 14879 6342 14927 6368
rect 467 6290 473 6342
rect 525 6290 537 6342
rect 589 6290 3209 6342
rect 3261 6290 3273 6342
rect 3325 6290 3331 6342
tri 14879 6294 14927 6342 ne
tri 14927 6294 15001 6368 sw
tri 14927 6290 14931 6294 ne
rect 14931 6290 15001 6294
tri 14931 6220 15001 6290 ne
tri 15001 6220 15075 6294 sw
tri 15001 6198 15023 6220 ne
rect 467 6136 473 6188
rect 525 6136 537 6188
rect 589 6136 3213 6188
rect 3265 6136 3277 6188
rect 3329 6136 3335 6188
rect 5999 6136 6005 6188
rect 6057 6136 6069 6188
rect 6121 6164 14669 6188
tri 14669 6164 14693 6188 sw
rect 6121 6136 14693 6164
tri 14693 6136 14721 6164 sw
tri 14647 6090 14693 6136 ne
rect 14693 6090 14721 6136
tri 14721 6090 14767 6136 sw
tri 14693 6068 14715 6090 ne
rect 348 5990 354 6042
rect 406 5990 418 6042
rect 470 5990 482 6042
rect 534 5990 546 6042
rect 598 5990 610 6042
rect 662 5990 674 6042
rect 726 5990 869 6042
rect 921 5990 933 6042
rect 985 5990 997 6042
rect 1049 5990 1061 6042
rect 1113 5990 1125 6042
rect 1177 5990 1189 6042
rect 1241 5990 1253 6042
rect 1305 5990 1317 6042
rect 1369 5990 1381 6042
rect 1433 5990 1445 6042
rect 1497 5990 1509 6042
rect 1561 5990 1573 6042
rect 1625 5990 1637 6042
rect 1689 5990 1701 6042
rect 1753 5990 1765 6042
rect 1817 5990 1829 6042
rect 1881 5990 1893 6042
rect 1945 5990 1957 6042
rect 2009 5990 2021 6042
rect 2073 5990 2085 6042
rect 2137 5990 2149 6042
rect 2201 5990 2213 6042
rect 2265 5990 2277 6042
rect 2329 5990 2341 6042
rect 2393 5990 2405 6042
rect 2457 5990 2469 6042
rect 2521 5990 2533 6042
rect 2585 5990 2597 6042
rect 2649 5990 2661 6042
rect 2713 5990 2725 6042
rect 2777 5990 2789 6042
rect 2841 5990 2853 6042
rect 2905 5990 2917 6042
rect 2969 5990 2981 6042
rect 3033 5990 3045 6042
rect 3097 5990 3109 6042
rect 3161 5990 3173 6042
rect 3225 5990 3237 6042
rect 3289 5990 3301 6042
rect 3353 5990 3365 6042
rect 3417 5990 3429 6042
rect 3481 5990 3493 6042
rect 3545 5990 3557 6042
rect 3609 5990 3621 6042
rect 3673 5990 3685 6042
rect 3737 5990 3749 6042
rect 3801 5990 3813 6042
rect 3865 5990 3877 6042
rect 3929 5990 3941 6042
rect 3993 5990 4005 6042
rect 4057 5990 4069 6042
rect 4121 5990 4133 6042
rect 4185 5990 4197 6042
rect 4249 5990 4261 6042
rect 4313 5990 4325 6042
rect 4377 5990 4389 6042
rect 4441 5990 4453 6042
rect 4505 5990 4517 6042
rect 4569 5990 4757 6042
rect 4809 5990 4821 6042
rect 4873 5990 4885 6042
rect 4937 5990 4949 6042
rect 5001 5990 5013 6042
rect 5065 5990 5077 6042
rect 5129 5990 5141 6042
rect 5193 5990 5205 6042
rect 5257 5990 5269 6042
rect 5321 5990 5333 6042
rect 5385 5990 5397 6042
rect 5449 5990 5461 6042
rect 5513 5990 5525 6042
rect 5577 5990 5589 6042
rect 5641 5990 5653 6042
rect 5705 5990 5717 6042
rect 5769 5990 5781 6042
rect 5833 5990 5845 6042
rect 5897 5990 6189 6042
rect 6241 5990 6254 6042
rect 6306 5990 6319 6042
rect 6371 5990 6384 6042
rect 6436 5990 6448 6042
rect 6500 5990 6512 6042
rect 6564 5990 6576 6042
rect 6628 5990 6640 6042
rect 6692 5990 6704 6042
rect 6756 5990 6768 6042
rect 6820 5990 7060 6042
rect 7112 5990 7124 6042
rect 7176 5990 7188 6042
rect 7240 5990 7252 6042
rect 7304 5990 7316 6042
rect 7368 5990 7380 6042
rect 7432 5990 7444 6042
rect 7496 5990 7508 6042
rect 7560 5990 7572 6042
rect 7624 5990 7923 6042
rect 7975 5990 7987 6042
rect 8039 5990 8051 6042
rect 8103 5990 8115 6042
rect 8167 5990 8179 6042
rect 8231 5990 8243 6042
rect 8295 5990 8307 6042
rect 8359 5990 8371 6042
rect 8423 5990 8435 6042
rect 8487 5990 8781 6042
rect 8833 5990 8845 6042
rect 8897 5990 8909 6042
rect 8961 5990 8973 6042
rect 9025 5990 9037 6042
rect 9089 5990 9101 6042
rect 9153 5990 9165 6042
rect 9217 5990 9229 6042
rect 9281 5990 9293 6042
rect 9345 5990 9619 6042
rect 9671 5990 9683 6042
rect 9735 5990 9747 6042
rect 9799 5990 9811 6042
rect 9863 5990 9875 6042
rect 9927 5990 9939 6042
rect 9991 5990 10003 6042
rect 10055 5990 10067 6042
rect 10119 5990 10131 6042
rect 10183 5990 10465 6042
rect 10517 5990 10529 6042
rect 10581 5990 10593 6042
rect 10645 5990 10657 6042
rect 10709 5990 10721 6042
rect 10773 5990 10785 6042
rect 10837 5990 10849 6042
rect 10901 5990 10913 6042
rect 10965 5990 10977 6042
rect 11029 5990 11041 6042
rect 11093 5990 11105 6042
rect 11157 5990 11169 6042
rect 11221 5990 11233 6042
rect 11285 5990 11297 6042
rect 11349 5990 11361 6042
rect 11413 5990 11425 6042
rect 11477 5990 11489 6042
rect 11541 5990 11553 6042
rect 11605 5990 11617 6042
rect 11669 5990 11681 6042
rect 11733 5990 11745 6042
rect 11797 5990 11809 6042
rect 11861 5990 11873 6042
rect 11925 5990 11937 6042
rect 11989 5990 12001 6042
rect 12053 5990 12065 6042
rect 12117 5990 12129 6042
rect 12181 5990 12193 6042
rect 12245 5990 12257 6042
rect 12309 5990 12321 6042
rect 12373 5990 12385 6042
rect 12437 5990 12449 6042
rect 12501 5990 12513 6042
rect 12565 5990 12577 6042
rect 12629 5990 12641 6042
rect 12693 5990 12705 6042
rect 12757 5990 12769 6042
rect 12821 5990 12833 6042
rect 12885 5990 12897 6042
rect 12949 5990 12961 6042
rect 13013 5990 13025 6042
rect 13077 5990 13089 6042
rect 13141 5990 13153 6042
rect 13205 5990 13217 6042
rect 13269 5990 13281 6042
rect 13333 5990 13345 6042
rect 13397 5990 13409 6042
rect 13461 5990 13473 6042
rect 13525 5990 13537 6042
rect 13589 5990 13601 6042
rect 13653 5990 13665 6042
rect 13717 5990 13729 6042
rect 13781 5990 13793 6042
rect 13845 5990 13857 6042
rect 13909 5990 13921 6042
rect 13973 5990 13985 6042
rect 14037 5990 14049 6042
rect 14101 5990 14114 6042
rect 14166 5990 14179 6042
rect 14231 5990 14244 6042
rect 14296 5990 14309 6042
rect 14361 5990 14374 6042
rect 14426 5990 14439 6042
rect 14491 5990 14504 6042
rect 14556 5990 14562 6042
tri 14709 5962 14715 5968 se
rect 14715 5962 14767 6090
rect 10986 5910 10992 5962
rect 11044 5910 11056 5962
rect 11108 5910 11390 5962
rect 11442 5910 11454 5962
rect 11506 5910 11512 5962
tri 14657 5910 14709 5962 se
rect 14709 5946 14767 5962
rect 14709 5910 14718 5946
tri 14644 5897 14657 5910 se
rect 14657 5897 14718 5910
tri 14718 5897 14767 5946 nw
tri 11878 5882 11893 5897 se
rect 11893 5882 14355 5897
rect 11613 5830 11619 5882
rect 11671 5830 11683 5882
rect 11735 5845 14355 5882
rect 14407 5845 14419 5897
rect 14471 5882 14703 5897
tri 14703 5882 14718 5897 nw
rect 14471 5845 14666 5882
tri 14666 5845 14703 5882 nw
rect 11735 5830 11900 5845
tri 11900 5830 11915 5845 nw
tri 15015 5830 15023 5838 se
rect 15023 5830 15075 6220
tri 14993 5808 15015 5830 se
rect 15015 5816 15075 5830
rect 15015 5808 15023 5816
rect 348 5756 354 5808
rect 406 5756 418 5808
rect 470 5756 482 5808
rect 534 5756 546 5808
rect 598 5756 610 5808
rect 662 5756 674 5808
rect 726 5756 738 5808
rect 790 5756 802 5808
rect 854 5756 866 5808
rect 918 5756 930 5808
rect 982 5756 994 5808
rect 1046 5756 1058 5808
rect 1110 5756 1122 5808
rect 1174 5756 1186 5808
rect 1238 5756 1250 5808
rect 1302 5756 1314 5808
rect 1366 5756 1378 5808
rect 1430 5756 1442 5808
rect 1494 5756 1506 5808
rect 1558 5756 1570 5808
rect 1622 5756 1634 5808
rect 1686 5756 1698 5808
rect 1750 5756 1762 5808
rect 1814 5756 1826 5808
rect 1878 5756 1890 5808
rect 1942 5756 1954 5808
rect 2006 5756 2018 5808
rect 2070 5756 2082 5808
rect 2134 5756 2146 5808
rect 2198 5756 2210 5808
rect 2262 5756 2274 5808
rect 2326 5756 2338 5808
rect 2390 5756 2402 5808
rect 2454 5756 2466 5808
rect 2518 5756 2530 5808
rect 2582 5756 2594 5808
rect 2646 5756 2658 5808
rect 2710 5756 2722 5808
rect 2774 5756 2786 5808
rect 2838 5756 2850 5808
rect 2902 5756 2914 5808
rect 2966 5756 2978 5808
rect 3030 5756 3042 5808
rect 3094 5756 3106 5808
rect 3158 5756 3170 5808
rect 3222 5756 3234 5808
rect 3286 5756 3298 5808
rect 3350 5756 3362 5808
rect 3414 5756 3427 5808
rect 3479 5756 3492 5808
rect 3544 5756 3557 5808
rect 3609 5756 3622 5808
rect 3674 5756 3687 5808
rect 3739 5756 3752 5808
rect 3804 5756 3817 5808
rect 3869 5756 3882 5808
rect 3934 5756 3947 5808
rect 3999 5756 4012 5808
rect 4064 5756 4077 5808
rect 4129 5756 4142 5808
rect 4194 5756 4207 5808
rect 4259 5756 4272 5808
rect 4324 5756 4337 5808
rect 4389 5756 4402 5808
rect 4454 5756 4467 5808
rect 4519 5756 4532 5808
rect 4584 5756 4597 5808
rect 4649 5756 4662 5808
rect 4714 5756 4727 5808
rect 4779 5756 4792 5808
rect 4844 5756 4857 5808
rect 4909 5756 4922 5808
rect 4974 5756 4987 5808
rect 5039 5756 5052 5808
rect 5104 5756 5117 5808
rect 5169 5756 5182 5808
rect 5234 5756 5247 5808
rect 5299 5756 5312 5808
rect 5364 5756 5377 5808
rect 5429 5756 5442 5808
rect 5494 5756 5507 5808
rect 5559 5756 5572 5808
rect 5624 5756 5637 5808
rect 5689 5756 5702 5808
rect 5754 5756 5767 5808
rect 5819 5756 5832 5808
rect 5884 5756 5897 5808
rect 5949 5756 6189 5808
rect 6241 5756 6254 5808
rect 6306 5756 6319 5808
rect 6371 5756 6384 5808
rect 6436 5756 6448 5808
rect 6500 5756 6512 5808
rect 6564 5756 6576 5808
rect 6628 5756 6640 5808
rect 6692 5756 6704 5808
rect 6756 5756 6768 5808
rect 6820 5756 7060 5808
rect 7112 5756 7124 5808
rect 7176 5756 7188 5808
rect 7240 5756 7252 5808
rect 7304 5756 7316 5808
rect 7368 5756 7380 5808
rect 7432 5756 7444 5808
rect 7496 5756 7508 5808
rect 7560 5756 7572 5808
rect 7624 5756 7923 5808
rect 7975 5756 7987 5808
rect 8039 5756 8051 5808
rect 8103 5756 8115 5808
rect 8167 5756 8179 5808
rect 8231 5756 8243 5808
rect 8295 5756 8307 5808
rect 8359 5756 8371 5808
rect 8423 5756 8435 5808
rect 8487 5756 8781 5808
rect 8833 5756 8845 5808
rect 8897 5756 8909 5808
rect 8961 5756 8973 5808
rect 9025 5756 9037 5808
rect 9089 5756 9101 5808
rect 9153 5756 9165 5808
rect 9217 5756 9229 5808
rect 9281 5756 9293 5808
rect 9345 5756 9619 5808
rect 9671 5756 9683 5808
rect 9735 5756 9747 5808
rect 9799 5756 9811 5808
rect 9863 5756 9875 5808
rect 9927 5756 9939 5808
rect 9991 5756 10003 5808
rect 10055 5756 10067 5808
rect 10119 5756 10131 5808
rect 10183 5756 10476 5808
rect 10528 5756 10540 5808
rect 10592 5756 10604 5808
rect 10656 5756 10668 5808
rect 10720 5756 10732 5808
rect 10784 5756 10796 5808
rect 10848 5756 10860 5808
rect 10912 5756 10918 5808
tri 14949 5764 14993 5808 se
rect 14993 5764 15023 5808
tri 15023 5764 15075 5816 nw
tri 14941 5756 14949 5764 se
tri 14928 5743 14941 5756 se
rect 14941 5743 14949 5756
rect 11613 5691 11619 5743
rect 11671 5691 11683 5743
rect 11735 5691 14359 5743
rect 14411 5691 14423 5743
rect 14475 5691 14481 5743
tri 14876 5691 14928 5743 se
rect 14928 5691 14949 5743
tri 14875 5690 14876 5691 se
rect 14876 5690 14949 5691
tri 14949 5690 15023 5764 nw
tri 14801 5616 14875 5690 se
tri 14875 5616 14949 5690 nw
tri 14774 5589 14801 5616 se
rect 14801 5589 14848 5616
tri 14848 5589 14875 5616 nw
rect 11613 5537 11619 5589
rect 11671 5537 11683 5589
rect 11735 5537 14355 5589
rect 14407 5537 14419 5589
rect 14471 5537 14796 5589
tri 14796 5537 14848 5589 nw
rect 292 5402 11553 5408
rect 292 5350 351 5402
rect 403 5350 471 5402
rect 523 5350 1327 5402
rect 1379 5350 2183 5402
rect 2235 5350 3039 5402
rect 3091 5350 3895 5402
rect 3947 5350 4751 5402
rect 4803 5350 5607 5402
rect 5659 5350 6463 5402
rect 6515 5350 7319 5402
rect 7371 5350 8175 5402
rect 8227 5350 9031 5402
rect 9083 5350 9887 5402
rect 9939 5350 10743 5402
rect 10795 5350 10863 5402
rect 10915 5350 11553 5402
rect 11613 5383 11619 5435
rect 11671 5383 11683 5435
rect 11735 5383 14359 5435
rect 14411 5383 14423 5435
rect 14475 5383 14481 5435
tri 15121 5383 15131 5393 se
rect 15131 5383 15183 6726
rect 292 5338 11553 5350
rect 292 5286 351 5338
rect 403 5286 471 5338
rect 523 5286 1327 5338
rect 1379 5286 2183 5338
rect 2235 5286 3039 5338
rect 3091 5286 3895 5338
rect 3947 5286 4751 5338
rect 4803 5286 5607 5338
rect 5659 5286 6463 5338
rect 6515 5286 7319 5338
rect 7371 5286 8175 5338
rect 8227 5286 9031 5338
rect 9083 5286 9887 5338
rect 9939 5286 10743 5338
rect 10795 5286 10863 5338
rect 10915 5286 11553 5338
tri 15057 5319 15121 5383 se
rect 15121 5371 15183 5383
rect 15121 5319 15131 5371
tri 15131 5319 15183 5371 nw
tri 15236 5319 15264 5347 se
rect 15264 5325 15316 6906
rect 292 5274 11553 5286
tri 15019 5281 15057 5319 se
rect 15057 5281 15093 5319
tri 15093 5281 15131 5319 nw
tri 15198 5281 15236 5319 se
rect 15236 5281 15264 5319
rect 292 5222 351 5274
rect 403 5222 471 5274
rect 523 5222 1327 5274
rect 1379 5222 2183 5274
rect 2235 5222 3039 5274
rect 3091 5222 3895 5274
rect 3947 5222 4751 5274
rect 4803 5222 5607 5274
rect 5659 5222 6463 5274
rect 6515 5222 7319 5274
rect 7371 5222 8175 5274
rect 8227 5222 9031 5274
rect 9083 5222 9887 5274
rect 9939 5222 10743 5274
rect 10795 5222 10863 5274
rect 10915 5222 11553 5274
rect 11613 5229 11619 5281
rect 11671 5229 11683 5281
rect 11735 5229 14355 5281
rect 14407 5229 14419 5281
rect 14471 5229 15041 5281
tri 15041 5229 15093 5281 nw
tri 15190 5273 15198 5281 se
rect 15198 5273 15264 5281
tri 15264 5273 15316 5325 nw
tri 15146 5229 15190 5273 se
rect 292 5210 11553 5222
rect 292 5158 351 5210
rect 403 5158 471 5210
rect 523 5158 1327 5210
rect 1379 5158 2183 5210
rect 2235 5158 3039 5210
rect 3091 5158 3895 5210
rect 3947 5158 4751 5210
rect 4803 5158 5607 5210
rect 5659 5158 6463 5210
rect 6515 5158 7319 5210
rect 7371 5158 8175 5210
rect 8227 5158 9031 5210
rect 9083 5158 9887 5210
rect 9939 5158 10743 5210
rect 10795 5158 10863 5210
rect 10915 5158 11553 5210
tri 15116 5199 15146 5229 se
rect 15146 5199 15190 5229
tri 15190 5199 15264 5273 nw
rect 292 5146 11553 5158
rect 292 5094 351 5146
rect 403 5094 471 5146
rect 523 5094 1327 5146
rect 1379 5094 2183 5146
rect 2235 5094 3039 5146
rect 3091 5094 3895 5146
rect 3947 5094 4751 5146
rect 4803 5094 5607 5146
rect 5659 5094 6463 5146
rect 6515 5094 7319 5146
rect 7371 5094 8175 5146
rect 8227 5094 9031 5146
rect 9083 5094 9887 5146
rect 9939 5094 10743 5146
rect 10795 5094 10863 5146
rect 10915 5094 11553 5146
tri 15044 5127 15116 5199 se
rect 292 5082 11553 5094
rect 292 5030 351 5082
rect 403 5030 471 5082
rect 523 5030 1327 5082
rect 1379 5030 2183 5082
rect 2235 5030 3039 5082
rect 3091 5030 3895 5082
rect 3947 5030 4751 5082
rect 4803 5030 5607 5082
rect 5659 5030 6463 5082
rect 6515 5030 7319 5082
rect 7371 5030 8175 5082
rect 8227 5030 9031 5082
rect 9083 5030 9887 5082
rect 9939 5030 10743 5082
rect 10795 5030 10863 5082
rect 10915 5030 11553 5082
rect 11613 5075 11619 5127
rect 11671 5075 11683 5127
rect 11735 5075 14359 5127
rect 14411 5075 14423 5127
rect 14475 5075 14481 5127
tri 15042 5125 15044 5127 se
rect 15044 5125 15116 5127
tri 15116 5125 15190 5199 nw
tri 15364 5125 15387 5148 se
rect 15387 5126 15439 6986
tri 14992 5075 15042 5125 se
tri 14968 5051 14992 5075 se
rect 14992 5051 15042 5075
tri 15042 5051 15116 5125 nw
tri 15313 5074 15364 5125 se
rect 15364 5074 15387 5125
tri 15387 5074 15439 5126 nw
tri 15290 5051 15313 5074 se
rect 292 5018 11553 5030
rect 292 4966 351 5018
rect 403 4966 471 5018
rect 523 4966 1327 5018
rect 1379 4966 2183 5018
rect 2235 4966 3039 5018
rect 3091 4966 3895 5018
rect 3947 4966 4751 5018
rect 4803 4966 5607 5018
rect 5659 4966 6463 5018
rect 6515 4966 7319 5018
rect 7371 4966 8175 5018
rect 8227 4966 9031 5018
rect 9083 4966 9887 5018
rect 9939 4966 10743 5018
rect 10795 4966 10863 5018
rect 10915 4966 11553 5018
tri 14894 4977 14968 5051 se
tri 14968 4977 15042 5051 nw
tri 15239 5000 15290 5051 se
rect 15290 5000 15313 5051
tri 15313 5000 15387 5074 nw
tri 15520 5000 15523 5003 se
rect 15523 5000 15575 7112
tri 15216 4977 15239 5000 se
tri 14890 4973 14894 4977 se
rect 14894 4973 14964 4977
tri 14964 4973 14968 4977 nw
tri 15212 4973 15216 4977 se
rect 15216 4973 15239 4977
rect 292 4954 11553 4966
rect 292 4902 351 4954
rect 403 4902 471 4954
rect 523 4902 1327 4954
rect 1379 4902 2183 4954
rect 2235 4902 3039 4954
rect 3091 4902 3895 4954
rect 3947 4902 4751 4954
rect 4803 4902 5607 4954
rect 5659 4902 6463 4954
rect 6515 4902 7319 4954
rect 7371 4902 8175 4954
rect 8227 4902 9031 4954
rect 9083 4902 9887 4954
rect 9939 4902 10743 4954
rect 10795 4902 10863 4954
rect 10915 4902 11553 4954
rect 11613 4921 11619 4973
rect 11671 4921 11683 4973
rect 11735 4921 14355 4973
rect 14407 4921 14419 4973
rect 14471 4921 14912 4973
tri 14912 4921 14964 4973 nw
tri 15165 4926 15212 4973 se
rect 15212 4926 15239 4973
tri 15239 4926 15313 5000 nw
tri 15449 4929 15520 5000 se
rect 15520 4981 15575 5000
rect 15520 4929 15523 4981
tri 15523 4929 15575 4981 nw
tri 15446 4926 15449 4929 se
tri 15160 4921 15165 4926 se
rect 292 4890 11553 4902
rect 292 4838 351 4890
rect 403 4838 471 4890
rect 523 4838 1327 4890
rect 1379 4838 2183 4890
rect 2235 4838 3039 4890
rect 3091 4838 3895 4890
rect 3947 4838 4751 4890
rect 4803 4838 5607 4890
rect 5659 4838 6463 4890
rect 6515 4838 7319 4890
rect 7371 4838 8175 4890
rect 8227 4838 9031 4890
rect 9083 4838 9887 4890
rect 9939 4838 10743 4890
rect 10795 4838 10863 4890
rect 10915 4838 11553 4890
tri 15091 4852 15160 4921 se
rect 15160 4852 15165 4921
tri 15165 4852 15239 4926 nw
tri 15375 4855 15446 4926 se
rect 15446 4855 15449 4926
tri 15449 4855 15523 4929 nw
tri 15372 4852 15375 4855 se
rect 292 4826 11553 4838
rect 292 4774 351 4826
rect 403 4774 471 4826
rect 523 4774 1327 4826
rect 1379 4774 2183 4826
rect 2235 4774 3039 4826
rect 3091 4774 3895 4826
rect 3947 4774 4751 4826
rect 4803 4774 5607 4826
rect 5659 4774 6463 4826
rect 6515 4774 7319 4826
rect 7371 4774 8175 4826
rect 8227 4774 9031 4826
rect 9083 4774 9887 4826
rect 9939 4774 10743 4826
rect 10795 4774 10863 4826
rect 10915 4774 11553 4826
tri 15058 4819 15091 4852 se
rect 292 4762 11553 4774
rect 11613 4767 11619 4819
rect 11671 4767 11683 4819
rect 11735 4767 14359 4819
rect 14411 4767 14423 4819
rect 14475 4767 14481 4819
tri 15017 4778 15058 4819 se
rect 15058 4778 15091 4819
tri 15091 4778 15165 4852 nw
tri 15301 4781 15372 4852 se
rect 15372 4781 15375 4852
tri 15375 4781 15449 4855 nw
tri 15298 4778 15301 4781 se
tri 15006 4767 15017 4778 se
rect 292 4710 351 4762
rect 403 4710 471 4762
rect 523 4710 1327 4762
rect 1379 4710 2183 4762
rect 2235 4710 3039 4762
rect 3091 4710 3895 4762
rect 3947 4710 4751 4762
rect 4803 4710 5607 4762
rect 5659 4710 6463 4762
rect 6515 4710 7319 4762
rect 7371 4710 8175 4762
rect 8227 4710 9031 4762
rect 9083 4710 9887 4762
rect 9939 4710 10743 4762
rect 10795 4710 10863 4762
rect 10915 4710 11553 4762
rect 292 4698 11553 4710
tri 14943 4704 15006 4767 se
rect 15006 4704 15017 4767
tri 15017 4704 15091 4778 nw
tri 15227 4707 15298 4778 se
rect 15298 4707 15301 4778
tri 15301 4707 15375 4781 nw
tri 15224 4704 15227 4707 se
rect 292 4646 351 4698
rect 403 4646 471 4698
rect 523 4646 1327 4698
rect 1379 4646 2183 4698
rect 2235 4646 3039 4698
rect 3091 4646 3895 4698
rect 3947 4646 4751 4698
rect 4803 4646 5607 4698
rect 5659 4646 6463 4698
rect 6515 4646 7319 4698
rect 7371 4646 8175 4698
rect 8227 4646 9031 4698
rect 9083 4646 9887 4698
rect 9939 4646 10743 4698
rect 10795 4646 10863 4698
rect 10915 4646 11553 4698
tri 14904 4665 14943 4704 se
rect 14943 4665 14978 4704
tri 14978 4665 15017 4704 nw
tri 15185 4665 15224 4704 se
rect 15224 4665 15227 4704
rect 292 4634 11553 4646
rect 292 4582 351 4634
rect 403 4582 471 4634
rect 523 4582 1327 4634
rect 1379 4582 2183 4634
rect 2235 4582 3039 4634
rect 3091 4582 3895 4634
rect 3947 4582 4751 4634
rect 4803 4582 5607 4634
rect 5659 4582 6463 4634
rect 6515 4582 7319 4634
rect 7371 4582 8175 4634
rect 8227 4582 9031 4634
rect 9083 4582 9887 4634
rect 9939 4582 10743 4634
rect 10795 4582 10863 4634
rect 10915 4582 11553 4634
rect 11613 4613 11619 4665
rect 11671 4613 11683 4665
rect 11735 4613 14355 4665
rect 14407 4613 14419 4665
rect 14471 4613 14926 4665
tri 14926 4613 14978 4665 nw
tri 15153 4633 15185 4665 se
rect 15185 4633 15227 4665
tri 15227 4633 15301 4707 nw
tri 15133 4613 15153 4633 se
rect 292 4570 11553 4582
rect 292 4518 351 4570
rect 403 4518 471 4570
rect 523 4518 1327 4570
rect 1379 4518 2183 4570
rect 2235 4518 3039 4570
rect 3091 4518 3895 4570
rect 3947 4518 4751 4570
rect 4803 4518 5607 4570
rect 5659 4518 6463 4570
rect 6515 4518 7319 4570
rect 7371 4518 8175 4570
rect 8227 4518 9031 4570
rect 9083 4518 9887 4570
rect 9939 4518 10743 4570
rect 10795 4518 10863 4570
rect 10915 4518 11553 4570
tri 15079 4559 15133 4613 se
rect 15133 4559 15153 4613
tri 15153 4559 15227 4633 nw
rect 292 4512 11553 4518
tri 15032 4512 15079 4559 se
tri 15031 4511 15032 4512 se
rect 15032 4511 15079 4512
rect 11613 4459 11619 4511
rect 11671 4459 11683 4511
rect 11735 4459 14359 4511
rect 14411 4459 14423 4511
rect 14475 4459 14481 4511
tri 15005 4485 15031 4511 se
rect 15031 4485 15079 4511
tri 15079 4485 15153 4559 nw
tri 14979 4459 15005 4485 se
tri 14931 4411 14979 4459 se
rect 14979 4411 15005 4459
tri 15005 4411 15079 4485 nw
tri 14877 4357 14931 4411 se
rect 14931 4357 14951 4411
tri 14951 4357 15005 4411 nw
rect 11613 4305 11619 4357
rect 11671 4305 11683 4357
rect 11735 4305 14355 4357
rect 14407 4305 14419 4357
rect 14471 4305 14899 4357
tri 14899 4305 14951 4357 nw
rect 11613 4151 11619 4203
rect 11671 4151 11683 4203
rect 11735 4151 14359 4203
rect 14411 4151 14423 4203
rect 14475 4151 14481 4203
rect 11613 3865 11619 3917
rect 11671 3865 11683 3917
rect 11735 3865 14359 3917
rect 14411 3865 14423 3917
rect 14475 3865 14481 3917
rect 15167 3865 15173 3917
rect 15225 3865 15237 3917
rect 15289 3865 15295 3917
rect 11613 3711 11619 3763
rect 11671 3711 11683 3763
rect 11735 3711 14355 3763
rect 14407 3711 14419 3763
rect 14471 3711 14477 3763
rect 14999 3711 15005 3763
rect 15057 3711 15069 3763
rect 15121 3711 15127 3763
rect 292 3637 11146 3643
rect 292 3585 491 3637
rect 543 3585 1347 3637
rect 1399 3585 2203 3637
rect 2255 3585 3059 3637
rect 3111 3585 3915 3637
rect 3967 3585 4771 3637
rect 4823 3585 5627 3637
rect 5679 3585 6483 3637
rect 6535 3585 7339 3637
rect 7391 3585 8195 3637
rect 8247 3585 9051 3637
rect 9103 3585 9907 3637
rect 9959 3585 10763 3637
rect 10815 3585 11146 3637
rect 292 3573 11146 3585
rect 292 3521 491 3573
rect 543 3521 1347 3573
rect 1399 3521 2203 3573
rect 2255 3521 3059 3573
rect 3111 3521 3915 3573
rect 3967 3521 4771 3573
rect 4823 3521 5627 3573
rect 5679 3521 6483 3573
rect 6535 3521 7339 3573
rect 7391 3521 8195 3573
rect 8247 3521 9051 3573
rect 9103 3521 9907 3573
rect 9959 3521 10763 3573
rect 10815 3521 11146 3573
rect 11613 3557 11619 3609
rect 11671 3557 11683 3609
rect 11735 3557 14359 3609
rect 14411 3557 14423 3609
rect 14475 3557 14481 3609
rect 292 3509 11146 3521
rect 292 3457 491 3509
rect 543 3457 1347 3509
rect 1399 3457 2203 3509
rect 2255 3457 3059 3509
rect 3111 3457 3915 3509
rect 3967 3457 4771 3509
rect 4823 3457 5627 3509
rect 5679 3457 6483 3509
rect 6535 3457 7339 3509
rect 7391 3457 8195 3509
rect 8247 3457 9051 3509
rect 9103 3457 9907 3509
rect 9959 3457 10763 3509
rect 10815 3457 11146 3509
rect 292 3445 11146 3457
rect 292 3393 491 3445
rect 543 3393 1347 3445
rect 1399 3393 2203 3445
rect 2255 3393 3059 3445
rect 3111 3393 3915 3445
rect 3967 3393 4771 3445
rect 4823 3393 5627 3445
rect 5679 3393 6483 3445
rect 6535 3393 7339 3445
rect 7391 3393 8195 3445
rect 8247 3393 9051 3445
rect 9103 3393 9907 3445
rect 9959 3393 10763 3445
rect 10815 3393 11146 3445
rect 11613 3403 11619 3455
rect 11671 3403 11683 3455
rect 11735 3403 14355 3455
rect 14407 3403 14419 3455
rect 14471 3403 14477 3455
rect 292 3381 11146 3393
rect 292 3329 491 3381
rect 543 3329 1347 3381
rect 1399 3329 2203 3381
rect 2255 3329 3059 3381
rect 3111 3329 3915 3381
rect 3967 3329 4771 3381
rect 4823 3329 5627 3381
rect 5679 3329 6483 3381
rect 6535 3329 7339 3381
rect 7391 3329 8195 3381
rect 8247 3329 9051 3381
rect 9103 3329 9907 3381
rect 9959 3329 10763 3381
rect 10815 3329 11146 3381
rect 292 3317 11146 3329
rect 292 3265 491 3317
rect 543 3265 1347 3317
rect 1399 3265 2203 3317
rect 2255 3265 3059 3317
rect 3111 3265 3915 3317
rect 3967 3265 4771 3317
rect 4823 3265 5627 3317
rect 5679 3265 6483 3317
rect 6535 3265 7339 3317
rect 7391 3265 8195 3317
rect 8247 3265 9051 3317
rect 9103 3265 9907 3317
rect 9959 3265 10763 3317
rect 10815 3265 11146 3317
rect 292 3253 11146 3265
rect 292 3201 491 3253
rect 543 3201 1347 3253
rect 1399 3201 2203 3253
rect 2255 3201 3059 3253
rect 3111 3201 3915 3253
rect 3967 3201 4771 3253
rect 4823 3201 5627 3253
rect 5679 3201 6483 3253
rect 6535 3201 7339 3253
rect 7391 3201 8195 3253
rect 8247 3201 9051 3253
rect 9103 3201 9907 3253
rect 9959 3201 10763 3253
rect 10815 3201 11146 3253
rect 11613 3249 11619 3301
rect 11671 3249 11683 3301
rect 11735 3249 14359 3301
rect 14411 3249 14423 3301
rect 14475 3249 14481 3301
rect 292 3189 11146 3201
rect 292 3137 491 3189
rect 543 3137 1347 3189
rect 1399 3137 2203 3189
rect 2255 3137 3059 3189
rect 3111 3137 3915 3189
rect 3967 3137 4771 3189
rect 4823 3137 5627 3189
rect 5679 3137 6483 3189
rect 6535 3137 7339 3189
rect 7391 3137 8195 3189
rect 8247 3137 9051 3189
rect 9103 3137 9907 3189
rect 9959 3137 10763 3189
rect 10815 3137 11146 3189
rect 292 3125 11146 3137
rect 292 3073 491 3125
rect 543 3073 1347 3125
rect 1399 3073 2203 3125
rect 2255 3073 3059 3125
rect 3111 3073 3915 3125
rect 3967 3073 4771 3125
rect 4823 3073 5627 3125
rect 5679 3073 6483 3125
rect 6535 3073 7339 3125
rect 7391 3073 8195 3125
rect 8247 3073 9051 3125
rect 9103 3073 9907 3125
rect 9959 3073 10763 3125
rect 10815 3073 11146 3125
rect 11613 3095 11619 3147
rect 11671 3095 11683 3147
rect 11735 3095 14355 3147
rect 14407 3095 14419 3147
rect 14471 3095 14477 3147
rect 292 3061 11146 3073
rect 292 3009 491 3061
rect 543 3009 1347 3061
rect 1399 3009 2203 3061
rect 2255 3009 3059 3061
rect 3111 3009 3915 3061
rect 3967 3009 4771 3061
rect 4823 3009 5627 3061
rect 5679 3009 6483 3061
rect 6535 3009 7339 3061
rect 7391 3009 8195 3061
rect 8247 3009 9051 3061
rect 9103 3009 9907 3061
rect 9959 3009 10763 3061
rect 10815 3009 11146 3061
rect 292 2997 11146 3009
rect 292 2945 491 2997
rect 543 2945 1347 2997
rect 1399 2945 2203 2997
rect 2255 2945 3059 2997
rect 3111 2945 3915 2997
rect 3967 2945 4771 2997
rect 4823 2945 5627 2997
rect 5679 2945 6483 2997
rect 6535 2945 7339 2997
rect 7391 2945 8195 2997
rect 8247 2945 9051 2997
rect 9103 2945 9907 2997
rect 9959 2945 10763 2997
rect 10815 2945 11146 2997
rect 292 2933 11146 2945
rect 11613 2941 11619 2993
rect 11671 2941 11683 2993
rect 11735 2941 14359 2993
rect 14411 2941 14423 2993
rect 14475 2941 14481 2993
rect 292 2881 491 2933
rect 543 2881 1347 2933
rect 1399 2881 2203 2933
rect 2255 2881 3059 2933
rect 3111 2881 3915 2933
rect 3967 2881 4771 2933
rect 4823 2881 5627 2933
rect 5679 2881 6483 2933
rect 6535 2881 7339 2933
rect 7391 2881 8195 2933
rect 8247 2881 9051 2933
rect 9103 2881 9907 2933
rect 9959 2881 10763 2933
rect 10815 2881 11146 2933
rect 292 2869 11146 2881
rect 292 2817 491 2869
rect 543 2817 1347 2869
rect 1399 2817 2203 2869
rect 2255 2817 3059 2869
rect 3111 2817 3915 2869
rect 3967 2817 4771 2869
rect 4823 2817 5627 2869
rect 5679 2817 6483 2869
rect 6535 2817 7339 2869
rect 7391 2817 8195 2869
rect 8247 2817 9051 2869
rect 9103 2817 9907 2869
rect 9959 2817 10763 2869
rect 10815 2817 11146 2869
rect 292 2805 11146 2817
rect 292 2753 491 2805
rect 543 2753 1347 2805
rect 1399 2753 2203 2805
rect 2255 2753 3059 2805
rect 3111 2753 3915 2805
rect 3967 2753 4771 2805
rect 4823 2753 5627 2805
rect 5679 2753 6483 2805
rect 6535 2753 7339 2805
rect 7391 2753 8195 2805
rect 8247 2753 9051 2805
rect 9103 2753 9907 2805
rect 9959 2753 10763 2805
rect 10815 2753 11146 2805
rect 11613 2787 11619 2839
rect 11671 2787 11683 2839
rect 11735 2787 14355 2839
rect 14407 2787 14419 2839
rect 14471 2787 14477 2839
rect 292 2747 11146 2753
rect 292 2685 11346 2691
rect 292 2633 351 2685
rect 403 2679 11346 2685
rect 403 2633 10904 2679
rect 292 2627 10904 2633
rect 10956 2627 11346 2679
rect 11613 2633 11619 2685
rect 11671 2633 11683 2685
rect 11735 2633 14359 2685
rect 14411 2633 14423 2685
rect 14475 2633 14481 2685
rect 292 2621 11346 2627
rect 292 2569 351 2621
rect 403 2615 11346 2621
rect 403 2569 10904 2615
rect 292 2563 10904 2569
rect 10956 2563 11346 2615
rect 292 2557 11346 2563
rect 292 2505 351 2557
rect 403 2550 11346 2557
rect 403 2505 10904 2550
rect 292 2498 10904 2505
rect 10956 2498 11346 2550
rect 292 2493 11346 2498
rect 292 2441 351 2493
rect 403 2485 11346 2493
rect 403 2441 10904 2485
rect 292 2433 10904 2441
rect 10956 2433 11346 2485
rect 11613 2479 11619 2531
rect 11671 2479 11683 2531
rect 11735 2479 14355 2531
rect 14407 2479 14419 2531
rect 14471 2479 14477 2531
rect 292 2429 11346 2433
rect 292 2377 351 2429
rect 403 2420 11346 2429
rect 403 2377 10904 2420
rect 292 2368 10904 2377
rect 10956 2368 11346 2420
rect 292 2365 11346 2368
rect 292 2313 351 2365
rect 403 2355 11346 2365
rect 403 2313 10904 2355
rect 292 2303 10904 2313
rect 10956 2303 11346 2355
rect 11613 2325 11619 2377
rect 11671 2325 11683 2377
rect 11735 2325 14359 2377
rect 14411 2325 14423 2377
rect 14475 2325 14481 2377
rect 292 2301 11346 2303
rect 292 2249 351 2301
rect 403 2249 11346 2301
rect 292 2232 11346 2249
rect 292 2180 381 2232
rect 433 2180 445 2232
rect 497 2180 509 2232
rect 561 2180 573 2232
rect 625 2180 637 2232
rect 689 2229 3209 2232
rect 689 2180 1047 2229
rect 292 2177 1047 2180
rect 1099 2177 1111 2229
rect 1163 2177 1175 2229
rect 1227 2177 1239 2229
rect 1291 2177 1436 2229
rect 1488 2177 1500 2229
rect 1552 2177 1564 2229
rect 1616 2177 1628 2229
rect 1680 2177 1890 2229
rect 1942 2177 1954 2229
rect 2006 2177 2018 2229
rect 2070 2177 2082 2229
rect 2134 2177 2295 2229
rect 2347 2177 2359 2229
rect 2411 2177 2423 2229
rect 2475 2177 2487 2229
rect 2539 2177 2759 2229
rect 2811 2177 2823 2229
rect 2875 2177 2887 2229
rect 2939 2177 2951 2229
rect 3003 2180 3209 2229
rect 3261 2180 3273 2232
rect 3325 2180 3337 2232
rect 3389 2180 3401 2232
rect 3453 2180 3465 2232
rect 3517 2180 3529 2232
rect 3581 2180 3593 2232
rect 3645 2229 11346 2232
rect 3645 2180 3971 2229
rect 3003 2177 3971 2180
rect 4023 2177 4035 2229
rect 4087 2177 4099 2229
rect 4151 2177 4163 2229
rect 4215 2177 4466 2229
rect 4518 2177 4530 2229
rect 4582 2177 4594 2229
rect 4646 2177 4658 2229
rect 4710 2177 4860 2229
rect 4912 2177 4924 2229
rect 4976 2177 4988 2229
rect 5040 2177 5052 2229
rect 5104 2177 5325 2229
rect 5377 2177 5389 2229
rect 5441 2177 5453 2229
rect 5505 2177 5517 2229
rect 5569 2177 5719 2229
rect 5771 2177 5783 2229
rect 5835 2177 5847 2229
rect 5899 2177 5911 2229
rect 5963 2177 6189 2229
rect 6241 2177 6253 2229
rect 6305 2177 6317 2229
rect 6369 2177 6381 2229
rect 6433 2177 6576 2229
rect 6628 2177 6640 2229
rect 6692 2177 6704 2229
rect 6756 2177 6768 2229
rect 6820 2177 6832 2229
rect 6884 2177 6896 2229
rect 6948 2177 6960 2229
rect 7012 2177 7024 2229
rect 7076 2177 7088 2229
rect 7140 2177 7152 2229
rect 7204 2177 7216 2229
rect 7268 2177 7280 2229
rect 7332 2177 7344 2229
rect 7396 2177 7408 2229
rect 7460 2177 7472 2229
rect 7524 2177 7536 2229
rect 7588 2177 7600 2229
rect 7652 2177 7664 2229
rect 7716 2177 7728 2229
rect 7780 2177 7792 2229
rect 7844 2177 7856 2229
rect 7908 2177 7920 2229
rect 7972 2177 7984 2229
rect 8036 2177 8048 2229
rect 8100 2177 8112 2229
rect 8164 2177 8176 2229
rect 8228 2177 8240 2229
rect 8292 2177 8304 2229
rect 8356 2177 8368 2229
rect 8420 2177 8432 2229
rect 8484 2177 8496 2229
rect 8548 2177 8560 2229
rect 8612 2177 8624 2229
rect 8676 2177 8688 2229
rect 8740 2177 8752 2229
rect 8804 2177 8816 2229
rect 8868 2177 8880 2229
rect 8932 2177 8944 2229
rect 8996 2177 9008 2229
rect 9060 2177 9072 2229
rect 9124 2177 9136 2229
rect 9188 2177 9200 2229
rect 9252 2177 9264 2229
rect 9316 2177 9328 2229
rect 9380 2177 9392 2229
rect 9444 2177 9456 2229
rect 9508 2177 9520 2229
rect 9572 2177 9584 2229
rect 9636 2177 9648 2229
rect 9700 2177 9712 2229
rect 9764 2177 9776 2229
rect 9828 2177 9840 2229
rect 9892 2177 9904 2229
rect 9956 2177 9968 2229
rect 10020 2177 10032 2229
rect 10084 2177 10096 2229
rect 10148 2177 10160 2229
rect 10212 2177 10224 2229
rect 10276 2177 10288 2229
rect 10340 2177 10352 2229
rect 10404 2177 10416 2229
rect 10468 2177 10480 2229
rect 10532 2177 10544 2229
rect 10596 2177 10608 2229
rect 10660 2177 10672 2229
rect 10724 2177 10736 2229
rect 10788 2177 10800 2229
rect 10852 2177 10864 2229
rect 10916 2177 11346 2229
rect 292 2154 11346 2177
rect 11613 2171 11619 2223
rect 11671 2171 11683 2223
rect 11735 2171 14355 2223
rect 14407 2171 14419 2223
rect 14471 2171 14477 2223
rect 292 2102 354 2154
rect 406 2102 418 2154
rect 470 2102 482 2154
rect 534 2102 546 2154
rect 598 2102 610 2154
rect 662 2102 674 2154
rect 726 2102 1047 2154
rect 1099 2102 1111 2154
rect 1163 2102 1175 2154
rect 1227 2102 1239 2154
rect 1291 2102 1436 2154
rect 1488 2102 1500 2154
rect 1552 2102 1564 2154
rect 1616 2102 1628 2154
rect 1680 2102 1890 2154
rect 1942 2102 1954 2154
rect 2006 2102 2018 2154
rect 2070 2102 2082 2154
rect 2134 2102 2295 2154
rect 2347 2102 2359 2154
rect 2411 2102 2423 2154
rect 2475 2102 2487 2154
rect 2539 2102 2759 2154
rect 2811 2102 2823 2154
rect 2875 2102 2887 2154
rect 2939 2102 2951 2154
rect 3003 2102 3209 2154
rect 3261 2102 3273 2154
rect 3325 2102 3337 2154
rect 3389 2102 3401 2154
rect 3453 2102 3465 2154
rect 3517 2102 3529 2154
rect 3581 2102 3593 2154
rect 3645 2102 3971 2154
rect 4023 2102 4035 2154
rect 4087 2102 4099 2154
rect 4151 2102 4163 2154
rect 4215 2102 4466 2154
rect 4518 2102 4530 2154
rect 4582 2102 4594 2154
rect 4646 2102 4658 2154
rect 4710 2102 4860 2154
rect 4912 2102 4924 2154
rect 4976 2102 4988 2154
rect 5040 2102 5052 2154
rect 5104 2102 5325 2154
rect 5377 2102 5389 2154
rect 5441 2102 5453 2154
rect 5505 2102 5517 2154
rect 5569 2102 5719 2154
rect 5771 2102 5783 2154
rect 5835 2102 5847 2154
rect 5899 2102 5911 2154
rect 5963 2102 6189 2154
rect 6241 2102 6253 2154
rect 6305 2102 6317 2154
rect 6369 2102 6381 2154
rect 6433 2102 6576 2154
rect 6628 2102 6641 2154
rect 6693 2102 6706 2154
rect 6758 2102 6771 2154
rect 6823 2102 6836 2154
rect 6888 2102 6901 2154
rect 6953 2102 6966 2154
rect 7018 2102 7031 2154
rect 7083 2102 7096 2154
rect 7148 2102 7161 2154
rect 7213 2102 7226 2154
rect 7278 2102 7291 2154
rect 7343 2102 7355 2154
rect 7407 2102 7419 2154
rect 7471 2102 7483 2154
rect 7535 2102 7547 2154
rect 7599 2102 7611 2154
rect 7663 2102 7675 2154
rect 7727 2102 7739 2154
rect 7791 2102 7803 2154
rect 7855 2102 7867 2154
rect 7919 2102 7931 2154
rect 7983 2102 7995 2154
rect 8047 2102 8059 2154
rect 8111 2102 8123 2154
rect 8175 2102 8187 2154
rect 8239 2102 8251 2154
rect 8303 2102 8315 2154
rect 8367 2102 8379 2154
rect 8431 2102 8443 2154
rect 8495 2102 8507 2154
rect 8559 2102 8571 2154
rect 8623 2102 8635 2154
rect 8687 2102 8699 2154
rect 8751 2102 8763 2154
rect 8815 2102 8827 2154
rect 8879 2102 8891 2154
rect 8943 2102 8955 2154
rect 9007 2102 9019 2154
rect 9071 2102 9083 2154
rect 9135 2102 9147 2154
rect 9199 2102 9211 2154
rect 9263 2102 9275 2154
rect 9327 2102 9339 2154
rect 9391 2102 9403 2154
rect 9455 2102 9467 2154
rect 9519 2102 9531 2154
rect 9583 2102 9595 2154
rect 9647 2102 9659 2154
rect 9711 2102 9723 2154
rect 9775 2102 9787 2154
rect 9839 2102 9851 2154
rect 9903 2102 9915 2154
rect 9967 2102 9979 2154
rect 10031 2102 10043 2154
rect 10095 2102 10107 2154
rect 10159 2102 10171 2154
rect 10223 2102 10235 2154
rect 10287 2102 10299 2154
rect 10351 2102 10363 2154
rect 10415 2102 10427 2154
rect 10479 2102 10491 2154
rect 10543 2102 10555 2154
rect 10607 2102 10619 2154
rect 10671 2102 10683 2154
rect 10735 2102 10747 2154
rect 10799 2102 10811 2154
rect 10863 2102 10875 2154
rect 10927 2102 11346 2154
rect 292 2078 11346 2102
rect 292 2075 3209 2078
rect 292 2023 354 2075
rect 406 2023 418 2075
rect 470 2023 482 2075
rect 534 2023 546 2075
rect 598 2023 610 2075
rect 662 2023 674 2075
rect 726 2023 1047 2075
rect 1099 2023 1111 2075
rect 1163 2023 1175 2075
rect 1227 2023 1239 2075
rect 1291 2023 1436 2075
rect 1488 2023 1500 2075
rect 1552 2023 1564 2075
rect 1616 2023 1628 2075
rect 1680 2023 1890 2075
rect 1942 2023 1954 2075
rect 2006 2023 2018 2075
rect 2070 2023 2082 2075
rect 2134 2023 2295 2075
rect 2347 2023 2359 2075
rect 2411 2023 2423 2075
rect 2475 2023 2487 2075
rect 2539 2023 2759 2075
rect 2811 2023 2823 2075
rect 2875 2023 2887 2075
rect 2939 2023 2951 2075
rect 3003 2026 3209 2075
rect 3261 2026 3273 2078
rect 3325 2026 3337 2078
rect 3389 2026 3401 2078
rect 3453 2026 3465 2078
rect 3517 2026 3529 2078
rect 3581 2026 3593 2078
rect 3645 2075 11346 2078
rect 3645 2026 3971 2075
rect 3003 2023 3971 2026
rect 4023 2023 4035 2075
rect 4087 2023 4099 2075
rect 4151 2023 4163 2075
rect 4215 2023 4466 2075
rect 4518 2023 4530 2075
rect 4582 2023 4594 2075
rect 4646 2023 4658 2075
rect 4710 2023 4860 2075
rect 4912 2023 4924 2075
rect 4976 2023 4988 2075
rect 5040 2023 5052 2075
rect 5104 2023 5325 2075
rect 5377 2023 5389 2075
rect 5441 2023 5453 2075
rect 5505 2023 5517 2075
rect 5569 2023 5719 2075
rect 5771 2023 5783 2075
rect 5835 2023 5847 2075
rect 5899 2023 5911 2075
rect 5963 2023 6189 2075
rect 6241 2023 6253 2075
rect 6305 2023 6317 2075
rect 6369 2023 6381 2075
rect 6433 2023 6582 2075
rect 6634 2023 6646 2075
rect 6698 2023 6710 2075
rect 6762 2023 6774 2075
rect 6826 2023 6838 2075
rect 6890 2023 6902 2075
rect 6954 2023 6966 2075
rect 7018 2023 7030 2075
rect 7082 2023 7094 2075
rect 7146 2023 7158 2075
rect 7210 2023 7222 2075
rect 7274 2023 7286 2075
rect 7338 2023 7350 2075
rect 7402 2023 7414 2075
rect 7466 2023 7478 2075
rect 7530 2023 7542 2075
rect 7594 2023 7606 2075
rect 7658 2023 7670 2075
rect 7722 2023 7734 2075
rect 7786 2023 7798 2075
rect 7850 2023 7862 2075
rect 7914 2023 7926 2075
rect 7978 2023 7990 2075
rect 8042 2023 8054 2075
rect 8106 2023 8118 2075
rect 8170 2023 8182 2075
rect 8234 2023 8246 2075
rect 8298 2023 8310 2075
rect 8362 2023 8374 2075
rect 8426 2023 8438 2075
rect 8490 2023 8502 2075
rect 8554 2023 8566 2075
rect 8618 2023 8630 2075
rect 8682 2023 8694 2075
rect 8746 2023 8758 2075
rect 8810 2023 8822 2075
rect 8874 2023 8886 2075
rect 8938 2023 8950 2075
rect 9002 2023 9014 2075
rect 9066 2023 9078 2075
rect 9130 2023 9142 2075
rect 9194 2023 9206 2075
rect 9258 2023 9270 2075
rect 9322 2023 9334 2075
rect 9386 2023 9398 2075
rect 9450 2023 9462 2075
rect 9514 2023 9526 2075
rect 9578 2023 9590 2075
rect 9642 2023 9654 2075
rect 9706 2023 9718 2075
rect 9770 2023 9782 2075
rect 9834 2023 9846 2075
rect 9898 2023 9910 2075
rect 9962 2023 9974 2075
rect 10026 2023 10038 2075
rect 10090 2023 10102 2075
rect 10154 2023 10166 2075
rect 10218 2023 10230 2075
rect 10282 2023 10294 2075
rect 10346 2023 10358 2075
rect 10410 2023 10422 2075
rect 10474 2023 10486 2075
rect 10538 2023 10550 2075
rect 10602 2023 10614 2075
rect 10666 2023 10678 2075
rect 10730 2023 10742 2075
rect 10794 2023 10806 2075
rect 10858 2023 10870 2075
rect 10922 2023 11346 2075
rect 11579 2026 11585 2078
rect 11637 2026 11649 2078
rect 11701 2026 11713 2078
rect 11765 2026 11777 2078
rect 11829 2026 11841 2078
rect 11893 2026 11905 2078
rect 11957 2026 11969 2078
rect 12021 2026 12033 2078
rect 12085 2026 12097 2078
rect 12149 2026 12161 2078
rect 12213 2026 12225 2078
rect 12277 2026 12289 2078
rect 12341 2026 12353 2078
rect 12405 2026 12417 2078
rect 12469 2026 12481 2078
rect 12533 2026 12545 2078
rect 12597 2026 12609 2078
rect 12661 2026 12673 2078
rect 12725 2026 12737 2078
rect 12789 2026 12801 2078
rect 12853 2026 12865 2078
rect 12917 2026 12929 2078
rect 12981 2026 12993 2078
rect 13045 2026 13057 2078
rect 13109 2026 13121 2078
rect 13173 2026 13185 2078
rect 13237 2026 13249 2078
rect 13301 2026 13313 2078
rect 13365 2026 13377 2078
rect 13429 2026 13441 2078
rect 13493 2026 13505 2078
rect 13557 2026 13569 2078
rect 13621 2026 13633 2078
rect 13685 2026 13697 2078
rect 13749 2026 13761 2078
rect 13813 2026 13825 2078
rect 13877 2026 13889 2078
rect 13941 2026 13953 2078
rect 14005 2026 14017 2078
rect 14069 2026 14081 2078
rect 14133 2026 14145 2078
rect 14197 2026 14209 2078
rect 14261 2026 14273 2078
rect 14325 2026 14337 2078
rect 14389 2026 14401 2078
rect 14453 2026 14465 2078
rect 14517 2026 14529 2078
rect 14581 2026 14593 2078
rect 14645 2026 14657 2078
rect 14709 2026 14721 2078
rect 14773 2026 14779 2078
rect 292 2021 11346 2023
rect 467 1881 473 1933
rect 525 1881 537 1933
rect 589 1881 1315 1933
rect 1367 1881 1379 1933
rect 1431 1881 3213 1933
rect 3265 1881 3277 1933
rect 3329 1881 5807 1933
rect 5859 1881 5871 1933
rect 5923 1881 5929 1933
rect 13248 1804 13254 1856
rect 13306 1804 13322 1856
rect 13374 1804 13390 1856
rect 13442 1804 13458 1856
rect 13510 1804 13526 1856
rect 13578 1804 13594 1856
rect 13646 1804 13662 1856
rect 13714 1804 13730 1856
rect 13782 1804 13788 1856
rect 467 1727 473 1779
rect 525 1727 537 1779
rect 589 1727 869 1779
rect 921 1727 933 1779
rect 985 1727 3209 1779
rect 3261 1727 3273 1779
rect 3325 1727 10789 1779
rect 10841 1727 10853 1779
rect 10905 1727 10911 1779
rect 467 1573 473 1625
rect 525 1573 537 1625
rect 589 1573 2171 1625
rect 2223 1573 2235 1625
rect 2287 1573 3213 1625
rect 3265 1573 3277 1625
rect 3329 1573 3335 1625
rect 467 1419 473 1471
rect 525 1419 537 1471
rect 589 1419 1725 1471
rect 1777 1419 1789 1471
rect 1841 1419 3209 1471
rect 3261 1419 3273 1471
rect 3325 1419 10789 1471
rect 10841 1419 10853 1471
rect 10905 1419 10911 1471
rect 13248 1394 13788 1804
rect 13248 1342 13254 1394
rect 13306 1342 13322 1394
rect 13374 1342 13390 1394
rect 13442 1342 13458 1394
rect 13510 1342 13526 1394
rect 13578 1342 13594 1394
rect 13646 1342 13662 1394
rect 13714 1342 13730 1394
rect 13782 1342 13788 1394
rect 467 1265 473 1317
rect 525 1265 537 1317
rect 589 1265 3213 1317
rect 3265 1265 3277 1317
rect 3329 1265 3335 1317
rect 467 1111 473 1163
rect 525 1111 537 1163
rect 589 1111 2581 1163
rect 2633 1111 2645 1163
rect 2697 1111 3209 1163
rect 3261 1111 3273 1163
rect 3325 1111 10789 1163
rect 10841 1111 10853 1163
rect 10905 1111 10911 1163
rect 13248 1086 13788 1342
rect 13248 1034 13254 1086
rect 13306 1034 13322 1086
rect 13374 1034 13390 1086
rect 13442 1034 13458 1086
rect 13510 1034 13526 1086
rect 13578 1034 13594 1086
rect 13646 1034 13662 1086
rect 13714 1034 13730 1086
rect 13782 1034 13788 1086
rect 467 957 473 1009
rect 525 957 537 1009
rect 589 957 3213 1009
rect 3265 957 3277 1009
rect 3329 957 4739 1009
rect 4791 957 4803 1009
rect 4855 957 4861 1009
rect 467 803 473 855
rect 525 803 537 855
rect 589 803 3209 855
rect 3261 803 3273 855
rect 3325 803 3762 855
rect 3814 803 3826 855
rect 3878 803 10789 855
rect 10841 803 10853 855
rect 10905 803 10911 855
rect 13248 778 13788 1034
rect 13248 726 13254 778
rect 13306 726 13322 778
rect 13374 726 13390 778
rect 13442 726 13458 778
rect 13510 726 13526 778
rect 13578 726 13594 778
rect 13646 726 13662 778
rect 13714 726 13730 778
rect 13782 726 13788 778
rect 467 649 473 701
rect 525 649 537 701
rect 589 649 3213 701
rect 3265 649 3277 701
rect 3329 649 5595 701
rect 5647 649 5659 701
rect 5711 649 5717 701
tri 13226 649 13248 671 se
rect 13248 649 13788 726
tri 13788 649 13810 671 sw
tri 13124 547 13226 649 se
rect 13226 547 13810 649
tri 13810 547 13912 649 sw
rect 467 495 473 547
rect 525 495 537 547
rect 589 495 3209 547
rect 3261 495 3273 547
rect 3325 495 4293 547
rect 4345 495 4357 547
rect 4409 495 10789 547
rect 10841 495 10853 547
rect 10905 495 10911 547
tri 13072 495 13124 547 se
rect 13124 495 13912 547
tri 13912 495 13964 547 sw
tri 13047 470 13072 495 se
rect 13072 470 13964 495
tri 13964 470 13989 495 sw
tri 12995 418 13047 470 se
rect 13047 418 13162 470
rect 13214 418 13232 470
rect 13284 418 13302 470
rect 13354 418 13372 470
rect 13424 418 13442 470
rect 13494 418 13511 470
rect 13563 418 13580 470
rect 13632 418 13649 470
rect 13701 418 13718 470
rect 13770 418 13787 470
rect 13839 418 13856 470
rect 13908 418 13925 470
rect 13977 418 13989 470
tri 12970 393 12995 418 se
rect 12995 393 13989 418
tri 13989 393 14066 470 sw
rect 14999 393 15127 3711
rect 467 341 473 393
rect 525 341 537 393
rect 589 341 3213 393
rect 3265 341 3277 393
rect 3329 341 6451 393
rect 6503 341 6515 393
rect 6567 341 6573 393
tri 12918 341 12970 393 se
rect 12970 341 14066 393
tri 14066 341 14118 393 sw
rect 14999 341 15005 393
rect 15057 341 15069 393
rect 15121 341 15127 393
tri 12816 239 12918 341 se
rect 12918 239 14118 341
tri 14118 239 14220 341 sw
rect 15167 239 15295 3865
rect 467 187 473 239
rect 525 187 537 239
rect 589 187 3209 239
rect 3261 187 3273 239
rect 3325 187 5149 239
rect 5201 187 5213 239
rect 5265 187 10789 239
rect 10841 187 10853 239
rect 10905 187 10911 239
tri 12764 187 12816 239 se
rect 12816 187 14220 239
tri 14220 187 14272 239 sw
rect 15167 187 15173 239
rect 15225 187 15237 239
rect 15289 187 15295 239
tri 12670 93 12764 187 se
rect 12764 93 14272 187
tri 14272 93 14366 187 sw
rect 357 41 363 93
rect 415 41 427 93
rect 479 41 491 93
rect 543 41 555 93
rect 607 41 619 93
rect 671 41 683 93
rect 735 41 886 93
rect 938 41 950 93
rect 1002 41 1014 93
rect 1066 41 1078 93
rect 1130 41 1142 93
rect 1194 41 1206 93
rect 1258 41 1270 93
rect 1322 41 1334 93
rect 1386 41 1398 93
rect 1450 41 1462 93
rect 1514 41 1526 93
rect 1578 41 1590 93
rect 1642 41 1654 93
rect 1706 41 1718 93
rect 1770 41 1782 93
rect 1834 41 1846 93
rect 1898 41 1910 93
rect 1962 41 1974 93
rect 2026 41 2038 93
rect 2090 41 2102 93
rect 2154 41 2166 93
rect 2218 41 2230 93
rect 2282 41 2294 93
rect 2346 41 2358 93
rect 2410 41 2422 93
rect 2474 41 2486 93
rect 2538 41 2550 93
rect 2602 41 2614 93
rect 2666 41 2678 93
rect 2730 41 2742 93
rect 2794 41 2806 93
rect 2858 41 2870 93
rect 2922 41 2934 93
rect 2986 41 2998 93
rect 3050 41 3062 93
rect 3114 41 3126 93
rect 3178 41 3190 93
rect 3242 41 3254 93
rect 3306 41 3318 93
rect 3370 41 3382 93
rect 3434 41 3446 93
rect 3498 41 3510 93
rect 3562 41 3574 93
rect 3626 41 3638 93
rect 3690 41 3702 93
rect 3754 41 3766 93
rect 3818 41 3830 93
rect 3882 41 3894 93
rect 3946 41 3958 93
rect 4010 41 4022 93
rect 4074 41 4086 93
rect 4138 41 4150 93
rect 4202 41 4214 93
rect 4266 41 4278 93
rect 4330 41 4342 93
rect 4394 41 4406 93
rect 4458 41 4470 93
rect 4522 41 4534 93
rect 4586 41 4598 93
rect 4650 41 4662 93
rect 4714 41 4726 93
rect 4778 41 4790 93
rect 4842 41 4854 93
rect 4906 41 4918 93
rect 4970 41 4982 93
rect 5034 41 5046 93
rect 5098 41 5110 93
rect 5162 41 5174 93
rect 5226 41 5238 93
rect 5290 41 5302 93
rect 5354 41 5366 93
rect 5418 41 5430 93
rect 5482 41 5494 93
rect 5546 41 5558 93
rect 5610 41 5622 93
rect 5674 41 5686 93
rect 5738 41 5750 93
rect 5802 41 5814 93
rect 5866 41 5878 93
rect 5930 41 5942 93
rect 5994 41 6006 93
rect 6058 41 6070 93
rect 6122 41 6134 93
rect 6186 41 6198 93
rect 6250 41 6262 93
rect 6314 41 6326 93
rect 6378 41 6390 93
rect 6442 41 6454 93
rect 6506 41 6518 93
rect 6570 41 6582 93
rect 6634 41 6646 93
rect 6698 41 6710 93
rect 6762 41 6774 93
rect 6826 41 6838 93
rect 6890 41 6902 93
rect 6954 41 6966 93
rect 7018 41 7030 93
rect 7082 41 7094 93
rect 7146 41 7158 93
rect 7210 41 7222 93
rect 7274 41 7286 93
rect 7338 41 7350 93
rect 7402 41 7414 93
rect 7466 41 7478 93
rect 7530 41 7542 93
rect 7594 41 7606 93
rect 7658 41 7670 93
rect 7722 41 7734 93
rect 7786 41 7798 93
rect 7850 41 7862 93
rect 7914 41 7926 93
rect 7978 41 7990 93
rect 8042 41 8054 93
rect 8106 41 8118 93
rect 8170 41 8182 93
rect 8234 41 8246 93
rect 8298 41 8310 93
rect 8362 41 8374 93
rect 8426 41 8438 93
rect 8490 41 8502 93
rect 8554 41 8566 93
rect 8618 41 8630 93
rect 8682 41 8694 93
rect 8746 41 8758 93
rect 8810 41 8822 93
rect 8874 41 8886 93
rect 8938 41 8950 93
rect 9002 41 9014 93
rect 9066 41 9078 93
rect 9130 41 9142 93
rect 9194 41 9206 93
rect 9258 41 9270 93
rect 9322 41 9334 93
rect 9386 41 9398 93
rect 9450 41 9462 93
rect 9514 41 9526 93
rect 9578 41 9590 93
rect 9642 41 9654 93
rect 9706 41 9718 93
rect 9770 41 9782 93
rect 9834 41 9846 93
rect 9898 41 9910 93
rect 9962 41 9974 93
rect 10026 41 10038 93
rect 10090 41 10102 93
rect 10154 41 10166 93
rect 10218 41 10230 93
rect 10282 41 10294 93
rect 10346 41 10358 93
rect 10410 41 10422 93
rect 10474 41 10486 93
rect 10538 41 10550 93
rect 10602 41 10614 93
rect 10666 41 10678 93
rect 10730 41 10742 93
rect 10794 41 10806 93
rect 10858 41 10870 93
rect 10922 41 10934 93
rect 10986 41 10998 93
rect 11050 41 11062 93
rect 11114 41 11126 93
rect 11178 41 11190 93
rect 11242 41 11254 93
rect 11306 41 11318 93
rect 11370 41 11382 93
rect 11434 41 11446 93
rect 11498 41 11510 93
rect 11562 41 11574 93
rect 11626 41 11638 93
rect 11690 41 11702 93
rect 11754 41 11766 93
rect 11818 41 11830 93
rect 11882 41 11894 93
rect 11946 41 11958 93
rect 12010 41 12022 93
rect 12074 41 12086 93
rect 12138 41 12150 93
rect 12202 41 12214 93
rect 12266 41 12278 93
rect 12330 41 12342 93
rect 12394 41 12406 93
rect 12458 41 12470 93
rect 12522 41 12534 93
rect 12586 41 12598 93
rect 12650 41 12662 93
rect 12714 41 12726 93
rect 12778 41 12790 93
rect 12842 41 12854 93
rect 12906 41 12918 93
rect 12970 41 12982 93
rect 13034 41 13046 93
rect 13098 41 13110 93
rect 13162 41 13174 93
rect 13226 41 13238 93
rect 13290 41 13302 93
rect 13354 41 13366 93
rect 13418 41 13430 93
rect 13482 41 13494 93
rect 13546 41 13558 93
rect 13610 41 13622 93
rect 13674 41 13686 93
rect 13738 41 13750 93
rect 13802 41 13814 93
rect 13866 41 13878 93
rect 13930 41 13942 93
rect 13994 41 14006 93
rect 14058 41 14070 93
rect 14122 41 14134 93
rect 14186 41 14198 93
rect 14250 41 14262 93
rect 14314 41 14326 93
rect 14378 41 16032 93
use sky130_fd_pr__via_l1m1__example_55959141808752  sky130_fd_pr__via_l1m1__example_55959141808752_0
timestamp 1619729480
transform 1 0 9896 0 -1 5411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808752  sky130_fd_pr__via_l1m1__example_55959141808752_1
timestamp 1619729480
transform 1 0 7328 0 -1 5411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808752  sky130_fd_pr__via_l1m1__example_55959141808752_2
timestamp 1619729480
transform 1 0 5616 0 -1 5411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808752  sky130_fd_pr__via_l1m1__example_55959141808752_3
timestamp 1619729480
transform 1 0 3048 0 -1 5411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808752  sky130_fd_pr__via_l1m1__example_55959141808752_4
timestamp 1619729480
transform 1 0 3904 0 -1 5411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808752  sky130_fd_pr__via_l1m1__example_55959141808752_5
timestamp 1619729480
transform 1 0 9040 0 -1 5411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808752  sky130_fd_pr__via_l1m1__example_55959141808752_6
timestamp 1619729480
transform 1 0 8184 0 -1 5411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808752  sky130_fd_pr__via_l1m1__example_55959141808752_7
timestamp 1619729480
transform 1 0 6472 0 -1 5411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808752  sky130_fd_pr__via_l1m1__example_55959141808752_8
timestamp 1619729480
transform 1 0 4760 0 -1 5411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808752  sky130_fd_pr__via_l1m1__example_55959141808752_9
timestamp 1619729480
transform 1 0 2192 0 -1 5411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808752  sky130_fd_pr__via_l1m1__example_55959141808752_10
timestamp 1619729480
transform 1 0 1336 0 -1 5411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808752  sky130_fd_pr__via_l1m1__example_55959141808752_11
timestamp 1619729480
transform 1 0 480 0 -1 5411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808752  sky130_fd_pr__via_l1m1__example_55959141808752_12
timestamp 1619729480
transform 1 0 500 0 -1 3646
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808752  sky130_fd_pr__via_l1m1__example_55959141808752_13
timestamp 1619729480
transform 1 0 10752 0 -1 5411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1619729480
transform 1 0 12882 0 -1 6179
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1619729480
transform 1 0 12882 0 -1 7873
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1619729480
transform 1 0 12882 0 -1 6949
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1619729480
transform 1 0 12882 0 -1 7257
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1619729480
transform 1 0 12882 0 -1 6487
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1619729480
transform 1 0 12882 0 -1 6641
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1619729480
transform 1 0 12882 0 -1 7411
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1619729480
transform 1 0 12882 0 -1 7565
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1619729480
transform 1 0 12882 0 -1 7719
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1619729480
transform 1 0 12882 0 -1 6333
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1619729480
transform -1 0 584 0 1 7839
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1619729480
transform 1 0 11624 0 -1 4194
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_12
timestamp 1619729480
transform 1 0 14526 0 -1 4194
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_13
timestamp 1619729480
transform 1 0 3380 0 1 7839
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_14
timestamp 1619729480
transform -1 0 11730 0 -1 4348
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_15
timestamp 1619729480
transform 1 0 478 0 1 7685
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_16
timestamp 1619729480
transform 1 0 3380 0 1 7685
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_17
timestamp 1619729480
transform 1 0 14526 0 -1 4348
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_18
timestamp 1619729480
transform -1 0 584 0 1 7223
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_19
timestamp 1619729480
transform 1 0 11624 0 -1 4810
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_20
timestamp 1619729480
transform 1 0 14526 0 -1 4810
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_21
timestamp 1619729480
transform 1 0 3380 0 1 7223
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_22
timestamp 1619729480
transform -1 0 584 0 1 6915
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_23
timestamp 1619729480
transform 1 0 11624 0 -1 5118
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_24
timestamp 1619729480
transform 1 0 14526 0 -1 5118
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_25
timestamp 1619729480
transform 1 0 3380 0 1 6915
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_26
timestamp 1619729480
transform -1 0 584 0 1 6299
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_27
timestamp 1619729480
transform 1 0 11624 0 -1 5734
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_28
timestamp 1619729480
transform 1 0 14526 0 -1 5734
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_29
timestamp 1619729480
transform 1 0 3380 0 1 6299
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_30
timestamp 1619729480
transform -1 0 11730 0 -1 2830
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_31
timestamp 1619729480
transform 1 0 478 0 1 1274
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_32
timestamp 1619729480
transform 1 0 3380 0 1 1274
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_33
timestamp 1619729480
transform 1 0 14526 0 -1 2830
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_34
timestamp 1619729480
transform -1 0 584 0 1 1428
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_35
timestamp 1619729480
transform 1 0 11624 0 -1 2676
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_36
timestamp 1619729480
transform 1 0 14526 0 -1 2676
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_37
timestamp 1619729480
transform 1 0 3380 0 1 1428
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_38
timestamp 1619729480
transform -1 0 584 0 1 1120
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_39
timestamp 1619729480
transform 1 0 11624 0 -1 2984
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_40
timestamp 1619729480
transform 1 0 14526 0 -1 2984
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_41
timestamp 1619729480
transform 1 0 3380 0 1 1120
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_42
timestamp 1619729480
transform -1 0 584 0 1 196
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_43
timestamp 1619729480
transform 1 0 11624 0 -1 3908
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_44
timestamp 1619729480
transform 1 0 14526 0 -1 3908
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_45
timestamp 1619729480
transform 1 0 3380 0 1 196
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_46
timestamp 1619729480
transform -1 0 584 0 1 504
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_47
timestamp 1619729480
transform 1 0 11624 0 -1 3600
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_48
timestamp 1619729480
transform 1 0 14526 0 -1 3600
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_49
timestamp 1619729480
transform 1 0 3380 0 1 504
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_50
timestamp 1619729480
transform -1 0 11730 0 -1 3446
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_51
timestamp 1619729480
transform 1 0 478 0 1 658
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_52
timestamp 1619729480
transform 1 0 3380 0 1 658
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_53
timestamp 1619729480
transform 1 0 14526 0 -1 3446
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_54
timestamp 1619729480
transform -1 0 11730 0 -1 2214
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_55
timestamp 1619729480
transform 1 0 478 0 1 1890
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_56
timestamp 1619729480
transform 1 0 3380 0 1 1890
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_57
timestamp 1619729480
transform 1 0 14526 0 -1 2214
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_58
timestamp 1619729480
transform -1 0 584 0 1 1736
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_59
timestamp 1619729480
transform 1 0 11624 0 -1 2368
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_60
timestamp 1619729480
transform 1 0 14526 0 -1 2368
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_61
timestamp 1619729480
transform 1 0 3380 0 1 1736
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_62
timestamp 1619729480
transform -1 0 11730 0 -1 5580
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_63
timestamp 1619729480
transform 1 0 478 0 1 6453
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_64
timestamp 1619729480
transform 1 0 3380 0 1 6453
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_65
timestamp 1619729480
transform 1 0 14526 0 -1 5580
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_66
timestamp 1619729480
transform -1 0 584 0 1 6607
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_67
timestamp 1619729480
transform 1 0 11624 0 -1 5426
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_68
timestamp 1619729480
transform 1 0 14526 0 -1 5426
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_69
timestamp 1619729480
transform 1 0 3380 0 1 6607
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_70
timestamp 1619729480
transform -1 0 11730 0 -1 4656
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_71
timestamp 1619729480
transform 1 0 478 0 1 7377
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_72
timestamp 1619729480
transform 1 0 3380 0 1 7377
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_73
timestamp 1619729480
transform 1 0 14526 0 -1 4656
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_74
timestamp 1619729480
transform -1 0 584 0 1 7531
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_75
timestamp 1619729480
transform 1 0 11624 0 -1 4502
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_76
timestamp 1619729480
transform 1 0 14526 0 -1 4502
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_77
timestamp 1619729480
transform 1 0 3380 0 1 7531
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_78
timestamp 1619729480
transform -1 0 11730 0 -1 5272
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_79
timestamp 1619729480
transform 1 0 478 0 1 6761
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_80
timestamp 1619729480
transform 1 0 3380 0 1 6761
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_81
timestamp 1619729480
transform 1 0 14526 0 -1 5272
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_82
timestamp 1619729480
transform -1 0 11730 0 -1 4964
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_83
timestamp 1619729480
transform 1 0 478 0 1 7069
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_84
timestamp 1619729480
transform 1 0 3380 0 1 7069
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_85
timestamp 1619729480
transform 1 0 14526 0 -1 4964
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_86
timestamp 1619729480
transform -1 0 11730 0 -1 2522
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_87
timestamp 1619729480
transform 1 0 478 0 1 1582
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_88
timestamp 1619729480
transform 1 0 3380 0 1 1582
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_89
timestamp 1619729480
transform 1 0 14526 0 -1 2522
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_90
timestamp 1619729480
transform -1 0 11730 0 -1 3138
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_91
timestamp 1619729480
transform 1 0 478 0 1 966
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_92
timestamp 1619729480
transform 1 0 3380 0 1 966
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_93
timestamp 1619729480
transform 1 0 14526 0 -1 3138
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_94
timestamp 1619729480
transform -1 0 584 0 1 812
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_95
timestamp 1619729480
transform 1 0 11624 0 -1 3292
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_96
timestamp 1619729480
transform 1 0 14526 0 -1 3292
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_97
timestamp 1619729480
transform 1 0 3380 0 1 812
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_98
timestamp 1619729480
transform -1 0 11730 0 -1 3754
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_99
timestamp 1619729480
transform 1 0 478 0 1 350
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_100
timestamp 1619729480
transform 1 0 3380 0 1 350
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_101
timestamp 1619729480
transform 1 0 14526 0 -1 3754
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_102
timestamp 1619729480
transform -1 0 11730 0 -1 5872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_103
timestamp 1619729480
transform 1 0 478 0 1 6145
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_104
timestamp 1619729480
transform 1 0 3380 0 1 6145
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_105
timestamp 1619729480
transform 1 0 14526 0 -1 5888
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_106
timestamp 1619729480
transform 1 0 12882 0 -1 692
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_107
timestamp 1619729480
transform 1 0 12882 0 -1 1000
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_108
timestamp 1619729480
transform 1 0 12882 0 -1 1924
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_109
timestamp 1619729480
transform 1 0 12882 0 -1 1616
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_110
timestamp 1619729480
transform 1 0 12882 0 -1 1462
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_111
timestamp 1619729480
transform 1 0 12882 0 -1 1308
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_112
timestamp 1619729480
transform 1 0 12882 0 -1 1154
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_113
timestamp 1619729480
transform 1 0 12882 0 -1 538
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_114
timestamp 1619729480
transform 1 0 12882 0 -1 384
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_115
timestamp 1619729480
transform 1 0 12882 0 -1 230
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_116
timestamp 1619729480
transform 1 0 12882 0 -1 1770
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_117
timestamp 1619729480
transform 1 0 12882 0 -1 6795
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_118
timestamp 1619729480
transform 1 0 12882 0 -1 7103
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_119
timestamp 1619729480
transform 1 0 12882 0 -1 846
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808751  sky130_fd_pr__via_l1m1__example_55959141808751_0
timestamp 1619729480
transform 1 0 360 0 -1 3790
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808751  sky130_fd_pr__via_l1m1__example_55959141808751_1
timestamp 1619729480
transform 1 0 360 0 1 4219
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808750  sky130_fd_pr__via_l1m1__example_55959141808750_0
timestamp 1619729480
transform 1 0 2212 0 -1 3664
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808750  sky130_fd_pr__via_l1m1__example_55959141808750_1
timestamp 1619729480
transform 1 0 9916 0 -1 3664
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808750  sky130_fd_pr__via_l1m1__example_55959141808750_2
timestamp 1619729480
transform 1 0 9060 0 -1 3664
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808750  sky130_fd_pr__via_l1m1__example_55959141808750_3
timestamp 1619729480
transform 1 0 6492 0 -1 3664
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808750  sky130_fd_pr__via_l1m1__example_55959141808750_4
timestamp 1619729480
transform 1 0 5636 0 -1 3664
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808750  sky130_fd_pr__via_l1m1__example_55959141808750_5
timestamp 1619729480
transform 1 0 3068 0 -1 3664
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808750  sky130_fd_pr__via_l1m1__example_55959141808750_6
timestamp 1619729480
transform 1 0 3924 0 -1 3664
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808750  sky130_fd_pr__via_l1m1__example_55959141808750_7
timestamp 1619729480
transform 1 0 4780 0 -1 3664
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808750  sky130_fd_pr__via_l1m1__example_55959141808750_8
timestamp 1619729480
transform 1 0 7348 0 -1 3664
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808750  sky130_fd_pr__via_l1m1__example_55959141808750_9
timestamp 1619729480
transform 1 0 8204 0 -1 3664
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808750  sky130_fd_pr__via_l1m1__example_55959141808750_10
timestamp 1619729480
transform 1 0 10772 0 -1 3664
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808750  sky130_fd_pr__via_l1m1__example_55959141808750_11
timestamp 1619729480
transform 1 0 1356 0 -1 3664
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808270  sky130_fd_pr__via_l1m1__example_55959141808270_0
timestamp 1619729480
transform -1 0 10881 0 1 5765
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808270  sky130_fd_pr__via_l1m1__example_55959141808270_1
timestamp 1619729480
transform 1 0 3219 0 1 2035
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808270  sky130_fd_pr__via_l1m1__example_55959141808270_2
timestamp 1619729480
transform 1 0 3219 0 1 2189
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1619729480
transform 1 0 456 0 1 2189
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1619729480
transform 1 0 1069 0 1 2189
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_2
timestamp 1619729480
transform 1 0 1069 0 1 2035
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_3
timestamp 1619729480
transform 1 0 1912 0 1 2035
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_4
timestamp 1619729480
transform 1 0 2781 0 1 2189
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_5
timestamp 1619729480
transform 1 0 2781 0 1 2035
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_6
timestamp 1619729480
transform 1 0 2317 0 1 2189
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_7
timestamp 1619729480
transform 1 0 2317 0 1 2035
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_8
timestamp 1619729480
transform 1 0 3993 0 1 2189
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_9
timestamp 1619729480
transform 1 0 4882 0 1 2189
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_10
timestamp 1619729480
transform 1 0 5741 0 1 2189
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_11
timestamp 1619729480
transform 1 0 3993 0 1 2035
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_12
timestamp 1619729480
transform 1 0 4882 0 1 2035
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_13
timestamp 1619729480
transform 1 0 5741 0 1 2035
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_14
timestamp 1619729480
transform 1 0 4488 0 1 2189
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_15
timestamp 1619729480
transform 1 0 5347 0 1 2035
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_16
timestamp 1619729480
transform 1 0 6211 0 1 2035
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_17
timestamp 1619729480
transform 1 0 4488 0 1 2035
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_18
timestamp 1619729480
transform 1 0 5347 0 1 2189
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_19
timestamp 1619729480
transform 1 0 6211 0 1 2189
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_20
timestamp 1619729480
transform 1 0 1912 0 1 2189
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_21
timestamp 1619729480
transform 1 0 1458 0 1 2189
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_22
timestamp 1619729480
transform 1 0 1458 0 1 2035
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808749  sky130_fd_pr__via_l1m1__example_55959141808749_0
timestamp 1619729480
transform 1 0 360 0 1 6094
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808749  sky130_fd_pr__via_l1m1__example_55959141808749_1
timestamp 1619729480
transform 1 0 360 0 1 154
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808749  sky130_fd_pr__via_l1m1__example_55959141808749_2
timestamp 1619729480
transform -1 0 11540 0 -1 3950
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808748  sky130_fd_pr__via_l1m1__example_55959141808748_0
timestamp 1619729480
transform 1 0 10912 0 -1 3790
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808748  sky130_fd_pr__via_l1m1__example_55959141808748_1
timestamp 1619729480
transform 1 0 10872 0 -1 5710
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808127  sky130_fd_pr__via_l1m1__example_55959141808127_0
timestamp 1619729480
transform 1 0 445 0 1 7984
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808127  sky130_fd_pr__via_l1m1__example_55959141808127_1
timestamp 1619729480
transform 1 0 449 0 1 2035
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808747  sky130_fd_pr__via_l1m1__example_55959141808747_0
timestamp 1619729480
transform -1 0 4548 0 1 5999
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808747  sky130_fd_pr__via_l1m1__example_55959141808747_1
timestamp 1619729480
transform 1 0 876 0 -1 8018
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808746  sky130_fd_pr__via_l1m1__example_55959141808746_0
timestamp 1619729480
transform 1 0 4766 0 1 7984
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808745  sky130_fd_pr__via_l1m1__example_55959141808745_0
timestamp 1619729480
transform -1 0 13580 0 1 7984
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_0
timestamp 1619729480
transform 1 0 9628 0 1 5765
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_1
timestamp 1619729480
transform 1 0 7932 0 1 5765
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_2
timestamp 1619729480
transform 1 0 7069 0 1 5765
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_3
timestamp 1619729480
transform 1 0 8790 0 1 5765
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_4
timestamp 1619729480
transform 1 0 9628 0 1 5999
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_5
timestamp 1619729480
transform 1 0 8790 0 1 5999
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_6
timestamp 1619729480
transform 1 0 7932 0 1 5999
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_7
timestamp 1619729480
transform 1 0 7069 0 1 5999
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808324  sky130_fd_pr__via_l1m1__example_55959141808324_0
timestamp 1619729480
transform -1 0 5887 0 1 5999
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808372  sky130_fd_pr__via_l1m1__example_55959141808372_0
timestamp 1619729480
transform 1 0 389 0 1 50
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808372  sky130_fd_pr__via_l1m1__example_55959141808372_1
timestamp 1619729480
transform 1 0 389 0 1 5999
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808744  sky130_fd_pr__via_l1m1__example_55959141808744_0
timestamp 1619729480
transform -1 0 10911 0 1 2189
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808744  sky130_fd_pr__via_l1m1__example_55959141808744_1
timestamp 1619729480
transform -1 0 10911 0 1 2035
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808743  sky130_fd_pr__via_l1m1__example_55959141808743_0
timestamp 1619729480
transform 1 0 915 0 1 50
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808742  sky130_fd_pr__via_l1m1__example_55959141808742_0
timestamp 1619729480
transform 1 0 11608 0 1 2035
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808741  sky130_fd_pr__via_l1m1__example_55959141808741_0
timestamp 1619729480
transform 1 0 10538 0 1 5999
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_0
timestamp 1619729480
transform 0 1 5688 1 0 4189
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_1
timestamp 1619729480
transform 0 1 5708 1 0 3753
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_2
timestamp 1619729480
transform 0 1 4832 1 0 4189
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_3
timestamp 1619729480
transform 0 1 3976 1 0 4189
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_4
timestamp 1619729480
transform 0 1 3996 1 0 3753
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_5
timestamp 1619729480
transform 0 1 552 1 0 4189
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_6
timestamp 1619729480
transform 0 1 1408 1 0 4189
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_7
timestamp 1619729480
transform 0 1 6564 1 0 3753
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_8
timestamp 1619729480
transform 0 1 2264 1 0 4189
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_9
timestamp 1619729480
transform 0 1 8276 1 0 3753
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_10
timestamp 1619729480
transform 0 1 7420 1 0 3753
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_11
timestamp 1619729480
transform 0 1 7400 1 0 4189
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_12
timestamp 1619729480
transform 0 1 8256 1 0 4189
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_13
timestamp 1619729480
transform 0 1 9132 1 0 3753
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_14
timestamp 1619729480
transform 0 1 9112 1 0 4189
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_15
timestamp 1619729480
transform 0 1 9968 1 0 4189
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_16
timestamp 1619729480
transform 0 1 9988 1 0 3753
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_17
timestamp 1619729480
transform 0 1 3140 1 0 3753
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_18
timestamp 1619729480
transform 0 1 3120 1 0 4189
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_19
timestamp 1619729480
transform 0 1 2284 1 0 3753
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_20
timestamp 1619729480
transform 0 1 572 1 0 3753
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_21
timestamp 1619729480
transform 0 1 1428 1 0 3753
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_22
timestamp 1619729480
transform 0 1 6544 1 0 4189
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_23
timestamp 1619729480
transform 0 1 4852 1 0 3753
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_0
timestamp 1619729480
transform 0 -1 2255 -1 0 3643
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_1
timestamp 1619729480
transform 0 -1 10795 -1 0 5408
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_2
timestamp 1619729480
transform 0 -1 9939 -1 0 5408
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_3
timestamp 1619729480
transform 0 -1 7371 -1 0 5408
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_4
timestamp 1619729480
transform 0 -1 5659 -1 0 5408
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_5
timestamp 1619729480
transform 0 -1 3967 -1 0 3643
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_6
timestamp 1619729480
transform 0 -1 4823 -1 0 3643
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_7
timestamp 1619729480
transform 0 -1 7391 -1 0 3643
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_8
timestamp 1619729480
transform 0 -1 8247 -1 0 3643
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_9
timestamp 1619729480
transform 0 -1 10815 -1 0 3643
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_10
timestamp 1619729480
transform 0 -1 3947 -1 0 5408
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_11
timestamp 1619729480
transform 0 -1 3091 -1 0 5408
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_12
timestamp 1619729480
transform 0 -1 9083 -1 0 5408
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_13
timestamp 1619729480
transform 0 -1 8227 -1 0 5408
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_14
timestamp 1619729480
transform 0 -1 6515 -1 0 5408
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_15
timestamp 1619729480
transform 0 -1 4803 -1 0 5408
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_16
timestamp 1619729480
transform 0 -1 2235 -1 0 5408
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_17
timestamp 1619729480
transform 0 -1 1379 -1 0 5408
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_18
timestamp 1619729480
transform 0 -1 523 -1 0 5408
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_19
timestamp 1619729480
transform 0 -1 9959 -1 0 3643
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_20
timestamp 1619729480
transform 0 -1 9103 -1 0 3643
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_21
timestamp 1619729480
transform 0 -1 6535 -1 0 3643
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_22
timestamp 1619729480
transform 0 -1 5679 -1 0 3643
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_23
timestamp 1619729480
transform 0 -1 3111 -1 0 3643
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_24
timestamp 1619729480
transform 0 -1 1399 -1 0 3643
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_25
timestamp 1619729480
transform 0 -1 543 -1 0 3643
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_26
timestamp 1619729480
transform 0 -1 10915 -1 0 5408
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808740  sky130_fd_pr__via_m1m2__example_55959141808740_27
timestamp 1619729480
transform 0 -1 403 -1 0 5408
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1619729480
transform 1 0 11613 0 -1 4203
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1619729480
transform -1 0 14481 0 -1 4203
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1619729480
transform -1 0 3331 0 1 7830
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1619729480
transform 1 0 467 0 1 7830
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_4
timestamp 1619729480
transform 1 0 467 0 1 7676
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_5
timestamp 1619729480
transform -1 0 3335 0 1 7676
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_6
timestamp 1619729480
transform -1 0 14477 0 -1 4357
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_7
timestamp 1619729480
transform 1 0 11613 0 -1 4357
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_8
timestamp 1619729480
transform 1 0 11613 0 -1 4819
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_9
timestamp 1619729480
transform -1 0 14481 0 -1 4819
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_10
timestamp 1619729480
transform -1 0 3331 0 1 7214
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_11
timestamp 1619729480
transform 1 0 467 0 1 7214
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_12
timestamp 1619729480
transform 1 0 11613 0 -1 5127
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_13
timestamp 1619729480
transform -1 0 14481 0 -1 5127
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_14
timestamp 1619729480
transform -1 0 3331 0 1 6906
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_15
timestamp 1619729480
transform 1 0 467 0 1 6906
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_16
timestamp 1619729480
transform 1 0 11613 0 -1 5743
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_17
timestamp 1619729480
transform -1 0 14481 0 -1 5743
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_18
timestamp 1619729480
transform -1 0 3331 0 1 6290
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_19
timestamp 1619729480
transform 1 0 467 0 1 6290
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_20
timestamp 1619729480
transform 1 0 467 0 1 1265
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_21
timestamp 1619729480
transform -1 0 3335 0 1 1265
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_22
timestamp 1619729480
transform -1 0 14477 0 -1 2839
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_23
timestamp 1619729480
transform 1 0 11613 0 -1 2839
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_24
timestamp 1619729480
transform 1 0 11613 0 -1 2685
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_25
timestamp 1619729480
transform -1 0 14481 0 -1 2685
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_26
timestamp 1619729480
transform -1 0 3331 0 1 1419
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_27
timestamp 1619729480
transform 1 0 467 0 1 1419
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_28
timestamp 1619729480
transform 1 0 11613 0 -1 2993
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_29
timestamp 1619729480
transform -1 0 14481 0 -1 2993
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_30
timestamp 1619729480
transform -1 0 3331 0 1 1111
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_31
timestamp 1619729480
transform 1 0 467 0 1 1111
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_32
timestamp 1619729480
transform 1 0 11613 0 -1 3917
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_33
timestamp 1619729480
transform -1 0 14481 0 -1 3917
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_34
timestamp 1619729480
transform -1 0 3331 0 1 187
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_35
timestamp 1619729480
transform 1 0 467 0 1 187
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_36
timestamp 1619729480
transform 1 0 11613 0 -1 3609
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_37
timestamp 1619729480
transform -1 0 14481 0 -1 3609
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_38
timestamp 1619729480
transform -1 0 3331 0 1 495
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_39
timestamp 1619729480
transform 1 0 467 0 1 495
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_40
timestamp 1619729480
transform 1 0 467 0 1 649
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_41
timestamp 1619729480
transform -1 0 3335 0 1 649
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_42
timestamp 1619729480
transform -1 0 14477 0 -1 3455
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_43
timestamp 1619729480
transform 1 0 11613 0 -1 3455
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_44
timestamp 1619729480
transform 1 0 467 0 1 1881
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_45
timestamp 1619729480
transform -1 0 3335 0 1 1881
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_46
timestamp 1619729480
transform -1 0 14477 0 -1 2223
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_47
timestamp 1619729480
transform 1 0 11613 0 -1 2223
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_48
timestamp 1619729480
transform 1 0 11613 0 -1 2377
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_49
timestamp 1619729480
transform -1 0 14481 0 -1 2377
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_50
timestamp 1619729480
transform -1 0 3331 0 1 1727
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_51
timestamp 1619729480
transform 1 0 467 0 1 1727
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_52
timestamp 1619729480
transform 1 0 467 0 1 6444
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_53
timestamp 1619729480
transform -1 0 3335 0 1 6444
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_54
timestamp 1619729480
transform -1 0 14477 0 -1 5589
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_55
timestamp 1619729480
transform 1 0 11613 0 -1 5589
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_56
timestamp 1619729480
transform 1 0 11613 0 -1 5435
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_57
timestamp 1619729480
transform -1 0 14481 0 -1 5435
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_58
timestamp 1619729480
transform -1 0 3331 0 1 6598
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_59
timestamp 1619729480
transform 1 0 467 0 1 6598
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_60
timestamp 1619729480
transform 1 0 467 0 1 7368
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_61
timestamp 1619729480
transform -1 0 3335 0 1 7368
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_62
timestamp 1619729480
transform -1 0 14477 0 -1 4665
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_63
timestamp 1619729480
transform 1 0 11613 0 -1 4665
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_64
timestamp 1619729480
transform 1 0 11613 0 -1 4511
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_65
timestamp 1619729480
transform -1 0 14481 0 -1 4511
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_66
timestamp 1619729480
transform -1 0 3331 0 1 7522
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_67
timestamp 1619729480
transform 1 0 467 0 1 7522
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_68
timestamp 1619729480
transform 1 0 467 0 1 6752
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_69
timestamp 1619729480
transform -1 0 3335 0 1 6752
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_70
timestamp 1619729480
transform -1 0 14477 0 -1 5281
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_71
timestamp 1619729480
transform 1 0 11613 0 -1 5281
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_72
timestamp 1619729480
transform 1 0 467 0 1 7060
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_73
timestamp 1619729480
transform -1 0 3335 0 1 7060
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_74
timestamp 1619729480
transform -1 0 14477 0 -1 4973
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_75
timestamp 1619729480
transform 1 0 11613 0 -1 4973
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_76
timestamp 1619729480
transform 1 0 467 0 1 1573
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_77
timestamp 1619729480
transform -1 0 3335 0 1 1573
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_78
timestamp 1619729480
transform -1 0 14477 0 -1 2531
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_79
timestamp 1619729480
transform 1 0 11613 0 -1 2531
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_80
timestamp 1619729480
transform 1 0 467 0 1 957
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_81
timestamp 1619729480
transform -1 0 3335 0 1 957
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_82
timestamp 1619729480
transform -1 0 14477 0 -1 3147
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_83
timestamp 1619729480
transform 1 0 11613 0 -1 3147
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_84
timestamp 1619729480
transform 1 0 11613 0 -1 3301
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_85
timestamp 1619729480
transform -1 0 14481 0 -1 3301
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_86
timestamp 1619729480
transform -1 0 3331 0 1 803
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_87
timestamp 1619729480
transform 1 0 467 0 1 803
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_88
timestamp 1619729480
transform 1 0 467 0 1 341
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_89
timestamp 1619729480
transform -1 0 3335 0 1 341
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_90
timestamp 1619729480
transform -1 0 14477 0 -1 3763
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_91
timestamp 1619729480
transform 1 0 11613 0 -1 3763
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_92
timestamp 1619729480
transform 1 0 467 0 1 6136
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_93
timestamp 1619729480
transform -1 0 3335 0 1 6136
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_94
timestamp 1619729480
transform -1 0 14477 0 -1 5897
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_95
timestamp 1619729480
transform 1 0 11613 0 -1 5882
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_96
timestamp 1619729480
transform 1 0 10279 0 1 7676
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_97
timestamp 1619729480
transform 1 0 9423 0 1 7368
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_98
timestamp 1619729480
transform 1 0 8567 0 1 7060
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_99
timestamp 1619729480
transform 1 0 7711 0 1 6752
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_100
timestamp 1619729480
transform 1 0 6855 0 1 6444
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_101
timestamp 1619729480
transform 1 0 5999 0 1 6136
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_102
timestamp 1619729480
transform -1 0 5929 0 1 1881
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_103
timestamp 1619729480
transform 1 0 863 0 1 1727
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_104
timestamp 1619729480
transform 1 0 1719 0 1 1419
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_105
timestamp 1619729480
transform 1 0 2575 0 1 1111
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_106
timestamp 1619729480
transform 1 0 3756 0 1 803
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_107
timestamp 1619729480
transform 1 0 4287 0 1 495
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_108
timestamp 1619729480
transform 1 0 5143 0 1 187
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_109
timestamp 1619729480
transform -1 0 1437 0 1 1881
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_110
timestamp 1619729480
transform 1 0 10986 0 1 5910
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_111
timestamp 1619729480
transform -1 0 10911 0 1 1419
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_112
timestamp 1619729480
transform -1 0 10911 0 1 1727
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_113
timestamp 1619729480
transform -1 0 10911 0 1 1111
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_114
timestamp 1619729480
transform -1 0 10911 0 1 803
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_115
timestamp 1619729480
transform -1 0 10911 0 1 495
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_116
timestamp 1619729480
transform -1 0 10911 0 1 187
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_117
timestamp 1619729480
transform -1 0 2293 0 1 1573
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_118
timestamp 1619729480
transform -1 0 4861 0 1 957
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_119
timestamp 1619729480
transform -1 0 5717 0 1 649
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_120
timestamp 1619729480
transform -1 0 6573 0 1 341
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808739  sky130_fd_pr__via_m1m2__example_55959141808739_0
timestamp 1619729480
transform 0 -1 403 1 0 2243
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808739  sky130_fd_pr__via_m1m2__example_55959141808739_1
timestamp 1619729480
transform 1 0 3203 0 1 2180
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808739  sky130_fd_pr__via_m1m2__example_55959141808739_2
timestamp 1619729480
transform -1 0 10918 0 1 5756
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808739  sky130_fd_pr__via_m1m2__example_55959141808739_3
timestamp 1619729480
transform 1 0 3203 0 1 2026
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808553  sky130_fd_pr__via_m1m2__example_55959141808553_0
timestamp 1619729480
transform 1 0 348 0 1 7975
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808553  sky130_fd_pr__via_m1m2__example_55959141808553_1
timestamp 1619729480
transform 1 0 348 0 1 5990
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808553  sky130_fd_pr__via_m1m2__example_55959141808553_2
timestamp 1619729480
transform 1 0 357 0 1 41
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808553  sky130_fd_pr__via_m1m2__example_55959141808553_3
timestamp 1619729480
transform 1 0 348 0 1 2023
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808738  sky130_fd_pr__via_m1m2__example_55959141808738_0
timestamp 1619729480
transform 1 0 863 0 1 5990
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808738  sky130_fd_pr__via_m1m2__example_55959141808738_1
timestamp 1619729480
transform 1 0 851 0 1 7975
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808737  sky130_fd_pr__via_m1m2__example_55959141808737_0
timestamp 1619729480
transform 1 0 4716 0 1 7975
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808736  sky130_fd_pr__via_m1m2__example_55959141808736_0
timestamp 1619729480
transform 1 0 6804 0 1 7975
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_0
timestamp 1619729480
transform 1 0 2289 0 1 2177
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_1
timestamp 1619729480
transform 1 0 2289 0 1 2023
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_2
timestamp 1619729480
transform 1 0 1884 0 1 2177
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_3
timestamp 1619729480
transform 1 0 1884 0 1 2023
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_4
timestamp 1619729480
transform 1 0 2753 0 1 2177
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_5
timestamp 1619729480
transform 1 0 2753 0 1 2023
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_6
timestamp 1619729480
transform 1 0 4460 0 1 2023
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_7
timestamp 1619729480
transform 1 0 5319 0 1 2177
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_8
timestamp 1619729480
transform 1 0 3965 0 1 2177
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_9
timestamp 1619729480
transform 1 0 4854 0 1 2177
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_10
timestamp 1619729480
transform 1 0 5713 0 1 2177
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_11
timestamp 1619729480
transform 1 0 3965 0 1 2023
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_12
timestamp 1619729480
transform 1 0 4854 0 1 2023
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_13
timestamp 1619729480
transform 1 0 5713 0 1 2023
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_14
timestamp 1619729480
transform 1 0 4460 0 1 2177
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_15
timestamp 1619729480
transform 1 0 5319 0 1 2023
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_16
timestamp 1619729480
transform 1 0 6183 0 1 2023
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_17
timestamp 1619729480
transform 1 0 6183 0 1 2177
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_18
timestamp 1619729480
transform 1 0 1041 0 1 2177
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_19
timestamp 1619729480
transform 1 0 1430 0 1 2177
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_20
timestamp 1619729480
transform 1 0 1041 0 1 2023
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808735  sky130_fd_pr__via_m1m2__example_55959141808735_21
timestamp 1619729480
transform 1 0 1430 0 1 2023
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808734  sky130_fd_pr__via_m1m2__example_55959141808734_0
timestamp 1619729480
transform 1 0 9613 0 1 5756
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808734  sky130_fd_pr__via_m1m2__example_55959141808734_1
timestamp 1619729480
transform 1 0 8775 0 1 5756
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808734  sky130_fd_pr__via_m1m2__example_55959141808734_2
timestamp 1619729480
transform 1 0 7054 0 1 5756
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808734  sky130_fd_pr__via_m1m2__example_55959141808734_3
timestamp 1619729480
transform 1 0 7917 0 1 5756
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808734  sky130_fd_pr__via_m1m2__example_55959141808734_4
timestamp 1619729480
transform 1 0 9613 0 1 5990
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808734  sky130_fd_pr__via_m1m2__example_55959141808734_5
timestamp 1619729480
transform 1 0 8775 0 1 5990
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808734  sky130_fd_pr__via_m1m2__example_55959141808734_6
timestamp 1619729480
transform 1 0 7917 0 1 5990
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808734  sky130_fd_pr__via_m1m2__example_55959141808734_7
timestamp 1619729480
transform 1 0 7054 0 1 5990
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808733  sky130_fd_pr__via_m1m2__example_55959141808733_0
timestamp 1619729480
transform 1 0 4751 0 1 5990
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808259  sky130_fd_pr__via_m1m2__example_55959141808259_0
timestamp 1619729480
transform 1 0 375 0 1 2180
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808732  sky130_fd_pr__via_m1m2__example_55959141808732_0
timestamp 1619729480
transform -1 0 10922 0 1 2177
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808732  sky130_fd_pr__via_m1m2__example_55959141808732_1
timestamp 1619729480
transform -1 0 10928 0 1 2023
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808731  sky130_fd_pr__via_m1m2__example_55959141808731_0
timestamp 1619729480
transform 1 0 880 0 1 41
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808730  sky130_fd_pr__via_m1m2__example_55959141808730_0
timestamp 1619729480
transform 1 0 11579 0 1 2026
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_0
timestamp 1619729480
transform -1 0 12994 0 -1 1474
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_1
timestamp 1619729480
transform -1 0 12994 0 -1 6345
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_2
timestamp 1619729480
transform -1 0 12994 0 -1 6961
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_3
timestamp 1619729480
transform -1 0 12994 0 -1 7885
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_4
timestamp 1619729480
transform 1 0 14520 0 -1 4206
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_5
timestamp 1619729480
transform 1 0 11618 0 -1 4206
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_6
timestamp 1619729480
transform -1 0 3492 0 1 7827
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_7
timestamp 1619729480
transform -1 0 590 0 1 7827
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_8
timestamp 1619729480
transform 1 0 3374 0 1 7673
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_9
timestamp 1619729480
transform 1 0 472 0 1 7673
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_10
timestamp 1619729480
transform -1 0 14638 0 -1 4360
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_11
timestamp 1619729480
transform -1 0 11736 0 -1 4360
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_12
timestamp 1619729480
transform 1 0 14520 0 -1 4822
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_13
timestamp 1619729480
transform 1 0 11618 0 -1 4822
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_14
timestamp 1619729480
transform -1 0 3492 0 1 7211
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_15
timestamp 1619729480
transform -1 0 590 0 1 7211
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_16
timestamp 1619729480
transform 1 0 12876 0 -1 7731
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_17
timestamp 1619729480
transform 1 0 14520 0 -1 5130
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_18
timestamp 1619729480
transform 1 0 11618 0 -1 5130
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_19
timestamp 1619729480
transform -1 0 3492 0 1 6903
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_20
timestamp 1619729480
transform -1 0 590 0 1 6903
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_21
timestamp 1619729480
transform 1 0 12876 0 -1 7115
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_22
timestamp 1619729480
transform 1 0 14520 0 -1 5746
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_23
timestamp 1619729480
transform 1 0 11618 0 -1 5746
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_24
timestamp 1619729480
transform -1 0 3492 0 1 6287
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_25
timestamp 1619729480
transform -1 0 590 0 1 6287
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_26
timestamp 1619729480
transform 1 0 3374 0 1 1262
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_27
timestamp 1619729480
transform 1 0 472 0 1 1262
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_28
timestamp 1619729480
transform -1 0 14638 0 -1 2842
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_29
timestamp 1619729480
transform -1 0 11736 0 -1 2842
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_30
timestamp 1619729480
transform 1 0 14520 0 -1 2688
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_31
timestamp 1619729480
transform 1 0 11618 0 -1 2688
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_32
timestamp 1619729480
transform -1 0 3492 0 1 1416
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_33
timestamp 1619729480
transform -1 0 590 0 1 1416
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_34
timestamp 1619729480
transform 1 0 14520 0 -1 2996
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_35
timestamp 1619729480
transform 1 0 11618 0 -1 2996
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_36
timestamp 1619729480
transform -1 0 3492 0 1 1108
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_37
timestamp 1619729480
transform -1 0 590 0 1 1108
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_38
timestamp 1619729480
transform 1 0 14520 0 -1 3920
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_39
timestamp 1619729480
transform 1 0 11618 0 -1 3920
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_40
timestamp 1619729480
transform -1 0 3492 0 1 184
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_41
timestamp 1619729480
transform -1 0 590 0 1 184
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_42
timestamp 1619729480
transform 1 0 14520 0 -1 3612
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_43
timestamp 1619729480
transform 1 0 11618 0 -1 3612
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_44
timestamp 1619729480
transform -1 0 3492 0 1 492
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_45
timestamp 1619729480
transform -1 0 590 0 1 492
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_46
timestamp 1619729480
transform 1 0 3374 0 1 646
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_47
timestamp 1619729480
transform 1 0 472 0 1 646
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_48
timestamp 1619729480
transform -1 0 14638 0 -1 3458
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_49
timestamp 1619729480
transform -1 0 11736 0 -1 3458
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_50
timestamp 1619729480
transform 1 0 3374 0 1 1878
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_51
timestamp 1619729480
transform 1 0 472 0 1 1878
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_52
timestamp 1619729480
transform -1 0 14638 0 -1 2226
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_53
timestamp 1619729480
transform -1 0 11736 0 -1 2226
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_54
timestamp 1619729480
transform 1 0 14520 0 -1 2380
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_55
timestamp 1619729480
transform 1 0 11618 0 -1 2380
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_56
timestamp 1619729480
transform -1 0 3492 0 1 1724
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_57
timestamp 1619729480
transform -1 0 590 0 1 1724
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_58
timestamp 1619729480
transform 1 0 3374 0 1 6441
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_59
timestamp 1619729480
transform 1 0 472 0 1 6441
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_60
timestamp 1619729480
transform -1 0 14638 0 -1 5592
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_61
timestamp 1619729480
transform -1 0 11736 0 -1 5592
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_62
timestamp 1619729480
transform 1 0 14520 0 -1 5438
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_63
timestamp 1619729480
transform 1 0 11618 0 -1 5438
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_64
timestamp 1619729480
transform -1 0 3492 0 1 6595
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_65
timestamp 1619729480
transform -1 0 590 0 1 6595
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_66
timestamp 1619729480
transform 1 0 3374 0 1 7365
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_67
timestamp 1619729480
transform 1 0 472 0 1 7365
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_68
timestamp 1619729480
transform -1 0 14638 0 -1 4668
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_69
timestamp 1619729480
transform -1 0 11736 0 -1 4668
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_70
timestamp 1619729480
transform 1 0 14520 0 -1 4514
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_71
timestamp 1619729480
transform 1 0 11618 0 -1 4514
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_72
timestamp 1619729480
transform -1 0 3492 0 1 7519
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_73
timestamp 1619729480
transform -1 0 590 0 1 7519
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_74
timestamp 1619729480
transform 1 0 3374 0 1 6749
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_75
timestamp 1619729480
transform 1 0 472 0 1 6749
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_76
timestamp 1619729480
transform -1 0 14638 0 -1 5284
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_77
timestamp 1619729480
transform -1 0 11736 0 -1 5284
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_78
timestamp 1619729480
transform 1 0 3374 0 1 7057
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_79
timestamp 1619729480
transform 1 0 472 0 1 7057
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_80
timestamp 1619729480
transform -1 0 14638 0 -1 4976
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_81
timestamp 1619729480
transform -1 0 11736 0 -1 4976
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_82
timestamp 1619729480
transform 1 0 3374 0 1 1570
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_83
timestamp 1619729480
transform 1 0 472 0 1 1570
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_84
timestamp 1619729480
transform -1 0 14638 0 -1 2534
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_85
timestamp 1619729480
transform -1 0 11736 0 -1 2534
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_86
timestamp 1619729480
transform 1 0 3374 0 1 954
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_87
timestamp 1619729480
transform 1 0 472 0 1 954
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_88
timestamp 1619729480
transform -1 0 14638 0 -1 3150
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_89
timestamp 1619729480
transform -1 0 11736 0 -1 3150
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_90
timestamp 1619729480
transform 1 0 14520 0 -1 3304
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_91
timestamp 1619729480
transform 1 0 11618 0 -1 3304
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_92
timestamp 1619729480
transform -1 0 3492 0 1 800
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_93
timestamp 1619729480
transform -1 0 590 0 1 800
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_94
timestamp 1619729480
transform 1 0 3374 0 1 338
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_95
timestamp 1619729480
transform 1 0 472 0 1 338
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_96
timestamp 1619729480
transform -1 0 14638 0 -1 3766
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_97
timestamp 1619729480
transform -1 0 11736 0 -1 3766
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_98
timestamp 1619729480
transform 1 0 3374 0 1 6133
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_99
timestamp 1619729480
transform 1 0 472 0 1 6133
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_100
timestamp 1619729480
transform -1 0 14638 0 -1 5900
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_101
timestamp 1619729480
transform -1 0 11736 0 -1 5900
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_102
timestamp 1619729480
transform 1 0 12876 0 -1 1628
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_103
timestamp 1619729480
transform -1 0 12994 0 -1 858
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_104
timestamp 1619729480
transform 1 0 12876 0 -1 704
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_105
timestamp 1619729480
transform 1 0 12876 0 -1 1012
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_106
timestamp 1619729480
transform 1 0 12876 0 -1 1936
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_107
timestamp 1619729480
transform -1 0 12994 0 -1 1782
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_108
timestamp 1619729480
transform 1 0 12876 0 -1 1320
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_109
timestamp 1619729480
transform -1 0 12994 0 -1 1166
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_110
timestamp 1619729480
transform -1 0 12994 0 -1 550
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_111
timestamp 1619729480
transform 1 0 12876 0 -1 396
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_112
timestamp 1619729480
transform -1 0 12994 0 -1 242
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_113
timestamp 1619729480
transform -1 0 12994 0 -1 6191
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_114
timestamp 1619729480
transform 1 0 12876 0 -1 6807
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_115
timestamp 1619729480
transform -1 0 12994 0 -1 7269
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_116
timestamp 1619729480
transform 1 0 12876 0 -1 6499
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_117
timestamp 1619729480
transform -1 0 12994 0 -1 6653
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_118
timestamp 1619729480
transform -1 0 12994 0 -1 7577
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808729  sky130_fd_pr__dfl1__example_55959141808729_119
timestamp 1619729480
transform 1 0 12876 0 -1 7423
box 0 0 1 1
use sky130_fd_pr__pfet_01v8__example_55959141808763  sky130_fd_pr__pfet_01v8__example_55959141808763_0
timestamp 1619729480
transform 1 0 525 0 1 4287
box -28 0 10244 675
use sky130_fd_pr__nfet_01v8__example_55959141808762  sky130_fd_pr__nfet_01v8__example_55959141808762_0
timestamp 1619729480
transform 1 0 545 0 1 2321
box -28 0 10244 675
use sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761  sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761_0
timestamp 1619729480
transform 1 0 5906 0 1 1881
box 0 5 92 17
use sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761  sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761_1
timestamp 1619729480
transform 1 0 10894 0 1 1419
box 0 5 92 17
use sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760  sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760_0
timestamp 1619729480
transform 0 -1 596 1 0 1631
box 0 5 92 17
use sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760  sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760_1
timestamp 1619729480
transform 0 1 11612 1 0 5136
box 0 5 92 17
use sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759  sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759_0
timestamp 1619729480
transform 0 -1 3114 1 0 1317
box 0 5 92 17
use sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759  sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759_1
timestamp 1619729480
transform 0 -1 4826 1 0 1009
box 0 5 92 17
use sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759  sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759_2
timestamp 1619729480
transform 0 -1 5682 1 0 701
box 0 5 92 17
use sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759  sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759_3
timestamp 1619729480
transform 0 -1 6538 1 0 393
box 0 5 92 17
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758_0
timestamp 1619729480
transform 0 1 11612 1 0 4520
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758_1
timestamp 1619729480
transform 0 1 11612 1 0 4828
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758_2
timestamp 1619729480
transform 0 -1 596 1 0 1328
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758_3
timestamp 1619729480
transform 0 -1 596 1 0 1020
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758_4
timestamp 1619729480
transform 0 -1 596 1 0 713
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758_5
timestamp 1619729480
transform 0 -1 596 1 0 405
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758_6
timestamp 1619729480
transform 0 1 11612 1 0 5444
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758_7
timestamp 1619729480
transform 0 1 11612 1 0 5752
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_0
timestamp 1619729480
transform 1 0 3307 0 1 7830
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_1
timestamp 1619729480
transform 1 0 14453 0 -1 4357
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_2
timestamp 1619729480
transform 1 0 3307 0 1 7214
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_3
timestamp 1619729480
transform 1 0 3307 0 1 6906
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_4
timestamp 1619729480
transform 1 0 3307 0 1 6290
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_5
timestamp 1619729480
transform 1 0 14453 0 -1 2839
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_6
timestamp 1619729480
transform 1 0 3307 0 1 1419
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_7
timestamp 1619729480
transform 1 0 3307 0 1 1111
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_8
timestamp 1619729480
transform 1 0 3307 0 1 187
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_9
timestamp 1619729480
transform 1 0 3307 0 1 495
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_10
timestamp 1619729480
transform 1 0 14453 0 -1 3455
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_11
timestamp 1619729480
transform 1 0 14453 0 -1 2223
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_12
timestamp 1619729480
transform 1 0 3307 0 1 1727
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_13
timestamp 1619729480
transform 1 0 14453 0 -1 5589
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_14
timestamp 1619729480
transform 1 0 3307 0 1 6598
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_15
timestamp 1619729480
transform 1 0 14453 0 -1 4665
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_16
timestamp 1619729480
transform 1 0 3307 0 1 7522
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_17
timestamp 1619729480
transform 1 0 14453 0 -1 5281
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_18
timestamp 1619729480
transform 1 0 14453 0 -1 4973
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_19
timestamp 1619729480
transform 1 0 14453 0 -1 2531
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_20
timestamp 1619729480
transform 1 0 14453 0 -1 3147
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_21
timestamp 1619729480
transform 1 0 3307 0 1 803
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_22
timestamp 1619729480
transform 1 0 14453 0 -1 3763
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_23
timestamp 1619729480
transform 1 0 14453 0 -1 5897
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_24
timestamp 1619729480
transform -1 0 14356 0 -1 5897
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_25
timestamp 1619729480
transform 1 0 10902 0 1 1727
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_26
timestamp 1619729480
transform 1 0 10902 0 1 1111
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_27
timestamp 1619729480
transform 1 0 10902 0 1 803
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_28
timestamp 1619729480
transform 1 0 10902 0 1 495
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757_29
timestamp 1619729480
transform 1 0 10902 0 1 187
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756_0
timestamp 1619729480
transform 0 -1 1402 1 0 1933
box 0 10 84 15
use sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756  sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756_1
timestamp 1619729480
transform 0 -1 2258 1 0 1625
box 0 10 84 15
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_0
timestamp 1619729480
transform -1 0 12884 0 1 7806
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_1
timestamp 1619729480
transform 1 0 3484 0 1 7652
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_2
timestamp 1619729480
transform -1 0 12884 0 1 7190
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_3
timestamp 1619729480
transform -1 0 12884 0 1 6882
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_4
timestamp 1619729480
transform -1 0 12884 0 1 6266
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_5
timestamp 1619729480
transform 1 0 3484 0 1 1241
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_6
timestamp 1619729480
transform -1 0 12884 0 1 1395
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_7
timestamp 1619729480
transform -1 0 12884 0 1 1087
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_8
timestamp 1619729480
transform -1 0 12884 0 1 163
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_9
timestamp 1619729480
transform -1 0 12884 0 1 471
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_10
timestamp 1619729480
transform 1 0 3484 0 1 625
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_11
timestamp 1619729480
transform 1 0 3484 0 1 1857
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_12
timestamp 1619729480
transform -1 0 12884 0 1 1703
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_13
timestamp 1619729480
transform 1 0 3484 0 1 6420
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_14
timestamp 1619729480
transform -1 0 12884 0 1 6574
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_15
timestamp 1619729480
transform 1 0 3484 0 1 7344
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_16
timestamp 1619729480
transform -1 0 12884 0 1 7498
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_17
timestamp 1619729480
transform 1 0 3484 0 1 6728
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_18
timestamp 1619729480
transform 1 0 3484 0 1 7036
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_19
timestamp 1619729480
transform 1 0 3484 0 1 1549
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_20
timestamp 1619729480
transform 1 0 3484 0 1 933
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_21
timestamp 1619729480
transform -1 0 12884 0 1 779
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_22
timestamp 1619729480
transform 1 0 3484 0 1 317
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808755  sky130_fd_pr__res_generic_nd__example_55959141808755_23
timestamp 1619729480
transform 1 0 3484 0 1 6112
box 7 21 9393 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_0
timestamp 1619729480
transform -1 0 3382 0 1 7806
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_1
timestamp 1619729480
transform 1 0 11728 0 -1 4227
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_2
timestamp 1619729480
transform -1 0 14528 0 -1 4381
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_3
timestamp 1619729480
transform 1 0 582 0 1 7652
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_4
timestamp 1619729480
transform -1 0 3382 0 1 7190
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_5
timestamp 1619729480
transform 1 0 11728 0 -1 4843
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_6
timestamp 1619729480
transform -1 0 3382 0 1 6882
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_7
timestamp 1619729480
transform 1 0 11728 0 -1 5151
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_8
timestamp 1619729480
transform -1 0 3382 0 1 6266
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_9
timestamp 1619729480
transform 1 0 11728 0 -1 5767
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_10
timestamp 1619729480
transform -1 0 14528 0 -1 2863
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_11
timestamp 1619729480
transform 1 0 582 0 1 1241
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_12
timestamp 1619729480
transform -1 0 3382 0 1 1395
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_13
timestamp 1619729480
transform 1 0 11728 0 -1 2709
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_14
timestamp 1619729480
transform -1 0 3382 0 1 1087
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_15
timestamp 1619729480
transform 1 0 11728 0 -1 3017
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_16
timestamp 1619729480
transform -1 0 3382 0 1 163
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_17
timestamp 1619729480
transform 1 0 11728 0 -1 3941
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_18
timestamp 1619729480
transform -1 0 3382 0 1 471
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_19
timestamp 1619729480
transform 1 0 11728 0 -1 3633
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_20
timestamp 1619729480
transform -1 0 14528 0 -1 3479
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_21
timestamp 1619729480
transform 1 0 582 0 1 625
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_22
timestamp 1619729480
transform -1 0 14528 0 -1 2247
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_23
timestamp 1619729480
transform 1 0 582 0 1 1857
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_24
timestamp 1619729480
transform -1 0 3382 0 1 1703
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_25
timestamp 1619729480
transform 1 0 11728 0 -1 2401
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_26
timestamp 1619729480
transform -1 0 14528 0 -1 5613
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_27
timestamp 1619729480
transform 1 0 582 0 1 6420
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_28
timestamp 1619729480
transform -1 0 3382 0 1 6574
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_29
timestamp 1619729480
transform 1 0 11728 0 -1 5459
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_30
timestamp 1619729480
transform -1 0 14528 0 -1 4689
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_31
timestamp 1619729480
transform 1 0 582 0 1 7344
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_32
timestamp 1619729480
transform -1 0 3382 0 1 7498
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_33
timestamp 1619729480
transform 1 0 11728 0 -1 4535
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_34
timestamp 1619729480
transform -1 0 14528 0 -1 5305
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_35
timestamp 1619729480
transform 1 0 582 0 1 6728
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_36
timestamp 1619729480
transform -1 0 14528 0 -1 4997
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_37
timestamp 1619729480
transform 1 0 582 0 1 7036
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_38
timestamp 1619729480
transform -1 0 14528 0 -1 2555
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_39
timestamp 1619729480
transform 1 0 582 0 1 1549
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_40
timestamp 1619729480
transform -1 0 14528 0 -1 3171
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_41
timestamp 1619729480
transform 1 0 582 0 1 933
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_42
timestamp 1619729480
transform -1 0 3382 0 1 779
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_43
timestamp 1619729480
transform 1 0 11728 0 -1 3325
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_44
timestamp 1619729480
transform -1 0 14528 0 -1 3787
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_45
timestamp 1619729480
transform 1 0 582 0 1 317
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_46
timestamp 1619729480
transform -1 0 14528 0 -1 5921
box 7 21 2793 22
use sky130_fd_pr__res_generic_nd__example_55959141808754  sky130_fd_pr__res_generic_nd__example_55959141808754_47
timestamp 1619729480
transform 1 0 582 0 1 6112
box 7 21 2793 22
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_0
timestamp 1619729480
transform 1 0 14451 0 -1 4203
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_1
timestamp 1619729480
transform 1 0 3305 0 1 7676
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_2
timestamp 1619729480
transform 1 0 14451 0 -1 4819
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_3
timestamp 1619729480
transform 1 0 14451 0 -1 5127
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_4
timestamp 1619729480
transform 1 0 14451 0 -1 5743
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_5
timestamp 1619729480
transform 1 0 3305 0 1 1265
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_6
timestamp 1619729480
transform 1 0 14451 0 -1 2685
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_7
timestamp 1619729480
transform 1 0 14451 0 -1 2993
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_8
timestamp 1619729480
transform 1 0 14451 0 -1 3917
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_9
timestamp 1619729480
transform 1 0 14451 0 -1 3609
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_10
timestamp 1619729480
transform 1 0 3305 0 1 649
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_11
timestamp 1619729480
transform 1 0 3305 0 1 1881
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_12
timestamp 1619729480
transform 1 0 14451 0 -1 2377
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_13
timestamp 1619729480
transform 1 0 3305 0 1 6444
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_14
timestamp 1619729480
transform 1 0 14451 0 -1 5435
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_15
timestamp 1619729480
transform 1 0 3305 0 1 7368
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_16
timestamp 1619729480
transform 1 0 14451 0 -1 4511
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_17
timestamp 1619729480
transform 1 0 3305 0 1 6752
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_18
timestamp 1619729480
transform 1 0 3305 0 1 7060
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_19
timestamp 1619729480
transform 1 0 3305 0 1 1573
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_20
timestamp 1619729480
transform 1 0 3305 0 1 957
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_21
timestamp 1619729480
transform 1 0 14451 0 -1 3301
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_22
timestamp 1619729480
transform 1 0 3305 0 1 341
box 0 5 92 17
use sky130_fd_io__xres_p_em1c_cdns_55959141808753  sky130_fd_io__xres_p_em1c_cdns_55959141808753_23
timestamp 1619729480
transform 1 0 3305 0 1 6136
box 0 5 92 17
<< labels >>
flabel metal2 s 609 4512 975 5408 0 FreeSans 1000 0 0 0 VCC_IO
flabel metal1 s 13684 8072 13736 8108 0 FreeSans 200 0 0 0 IN
flabel comment s 14150 7937 14150 7937 0 FreeSans 400 0 0 0 OUT
flabel comment s 13708 7937 13708 7937 0 FreeSans 400 0 0 0 IN
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 4992388
string GDS_START 4457654
<< end >>
