magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1260 -1260 1560 4260
<< locali >>
rect 0 2861 300 3000
rect 0 2827 61 2861
rect 95 2827 133 2861
rect 167 2827 205 2861
rect 239 2827 300 2861
rect 0 2765 300 2827
rect 0 2731 61 2765
rect 95 2731 133 2765
rect 167 2731 205 2765
rect 239 2731 300 2765
rect 0 2669 300 2731
rect 0 2635 61 2669
rect 95 2635 133 2669
rect 167 2635 205 2669
rect 239 2635 300 2669
rect 0 2573 300 2635
rect 0 2539 61 2573
rect 95 2539 133 2573
rect 167 2539 205 2573
rect 239 2539 300 2573
rect 0 2477 300 2539
rect 0 2443 61 2477
rect 95 2443 133 2477
rect 167 2443 205 2477
rect 239 2443 300 2477
rect 0 2381 300 2443
rect 0 2347 61 2381
rect 95 2347 133 2381
rect 167 2347 205 2381
rect 239 2347 300 2381
rect 0 2285 300 2347
rect 0 2251 61 2285
rect 95 2251 133 2285
rect 167 2251 205 2285
rect 239 2251 300 2285
rect 0 2189 300 2251
rect 0 2155 61 2189
rect 95 2155 133 2189
rect 167 2155 205 2189
rect 239 2155 300 2189
rect 0 2093 300 2155
rect 0 2059 61 2093
rect 95 2059 133 2093
rect 167 2059 205 2093
rect 239 2059 300 2093
rect 0 1997 300 2059
rect 0 1963 61 1997
rect 95 1963 133 1997
rect 167 1963 205 1997
rect 239 1963 300 1997
rect 0 1901 300 1963
rect 0 1867 61 1901
rect 95 1867 133 1901
rect 167 1867 205 1901
rect 239 1867 300 1901
rect 0 1805 300 1867
rect 0 1771 61 1805
rect 95 1771 133 1805
rect 167 1771 205 1805
rect 239 1771 300 1805
rect 0 1709 300 1771
rect 0 1675 61 1709
rect 95 1675 133 1709
rect 167 1675 205 1709
rect 239 1675 300 1709
rect 0 1613 300 1675
rect 0 1579 61 1613
rect 95 1579 133 1613
rect 167 1579 205 1613
rect 239 1579 300 1613
rect 0 1517 300 1579
rect 0 1483 61 1517
rect 95 1483 133 1517
rect 167 1483 205 1517
rect 239 1483 300 1517
rect 0 1421 300 1483
rect 0 1387 61 1421
rect 95 1387 133 1421
rect 167 1387 205 1421
rect 239 1387 300 1421
rect 0 1325 300 1387
rect 0 1291 61 1325
rect 95 1291 133 1325
rect 167 1291 205 1325
rect 239 1291 300 1325
rect 0 1229 300 1291
rect 0 1195 61 1229
rect 95 1195 133 1229
rect 167 1195 205 1229
rect 239 1195 300 1229
rect 0 1133 300 1195
rect 0 1099 61 1133
rect 95 1099 133 1133
rect 167 1099 205 1133
rect 239 1099 300 1133
rect 0 1037 300 1099
rect 0 1003 61 1037
rect 95 1003 133 1037
rect 167 1003 205 1037
rect 239 1003 300 1037
rect 0 941 300 1003
rect 0 907 61 941
rect 95 907 133 941
rect 167 907 205 941
rect 239 907 300 941
rect 0 845 300 907
rect 0 811 61 845
rect 95 811 133 845
rect 167 811 205 845
rect 239 811 300 845
rect 0 749 300 811
rect 0 715 61 749
rect 95 715 133 749
rect 167 715 205 749
rect 239 715 300 749
rect 0 653 300 715
rect 0 619 61 653
rect 95 619 133 653
rect 167 619 205 653
rect 239 619 300 653
rect 0 557 300 619
rect 0 523 61 557
rect 95 523 133 557
rect 167 523 205 557
rect 239 523 300 557
rect 0 461 300 523
rect 0 427 61 461
rect 95 427 133 461
rect 167 427 205 461
rect 239 427 300 461
rect 0 365 300 427
rect 0 331 61 365
rect 95 331 133 365
rect 167 331 205 365
rect 239 331 300 365
rect 0 269 300 331
rect 0 235 61 269
rect 95 235 133 269
rect 167 235 205 269
rect 239 235 300 269
rect 0 173 300 235
rect 0 139 61 173
rect 95 139 133 173
rect 167 139 205 173
rect 239 139 300 173
rect 0 0 300 139
<< viali >>
rect 61 2827 95 2861
rect 133 2827 167 2861
rect 205 2827 239 2861
rect 61 2731 95 2765
rect 133 2731 167 2765
rect 205 2731 239 2765
rect 61 2635 95 2669
rect 133 2635 167 2669
rect 205 2635 239 2669
rect 61 2539 95 2573
rect 133 2539 167 2573
rect 205 2539 239 2573
rect 61 2443 95 2477
rect 133 2443 167 2477
rect 205 2443 239 2477
rect 61 2347 95 2381
rect 133 2347 167 2381
rect 205 2347 239 2381
rect 61 2251 95 2285
rect 133 2251 167 2285
rect 205 2251 239 2285
rect 61 2155 95 2189
rect 133 2155 167 2189
rect 205 2155 239 2189
rect 61 2059 95 2093
rect 133 2059 167 2093
rect 205 2059 239 2093
rect 61 1963 95 1997
rect 133 1963 167 1997
rect 205 1963 239 1997
rect 61 1867 95 1901
rect 133 1867 167 1901
rect 205 1867 239 1901
rect 61 1771 95 1805
rect 133 1771 167 1805
rect 205 1771 239 1805
rect 61 1675 95 1709
rect 133 1675 167 1709
rect 205 1675 239 1709
rect 61 1579 95 1613
rect 133 1579 167 1613
rect 205 1579 239 1613
rect 61 1483 95 1517
rect 133 1483 167 1517
rect 205 1483 239 1517
rect 61 1387 95 1421
rect 133 1387 167 1421
rect 205 1387 239 1421
rect 61 1291 95 1325
rect 133 1291 167 1325
rect 205 1291 239 1325
rect 61 1195 95 1229
rect 133 1195 167 1229
rect 205 1195 239 1229
rect 61 1099 95 1133
rect 133 1099 167 1133
rect 205 1099 239 1133
rect 61 1003 95 1037
rect 133 1003 167 1037
rect 205 1003 239 1037
rect 61 907 95 941
rect 133 907 167 941
rect 205 907 239 941
rect 61 811 95 845
rect 133 811 167 845
rect 205 811 239 845
rect 61 715 95 749
rect 133 715 167 749
rect 205 715 239 749
rect 61 619 95 653
rect 133 619 167 653
rect 205 619 239 653
rect 61 523 95 557
rect 133 523 167 557
rect 205 523 239 557
rect 61 427 95 461
rect 133 427 167 461
rect 205 427 239 461
rect 61 331 95 365
rect 133 331 167 365
rect 205 331 239 365
rect 61 235 95 269
rect 133 235 167 269
rect 205 235 239 269
rect 61 139 95 173
rect 133 139 167 173
rect 205 139 239 173
<< metal1 >>
tri 0 2940 60 3000 se
rect 60 2940 240 3000
tri 240 2940 300 3000 sw
rect 0 2861 300 2940
rect 0 2827 61 2861
rect 95 2827 133 2861
rect 167 2827 205 2861
rect 239 2827 300 2861
rect 0 2765 300 2827
rect 0 2731 61 2765
rect 95 2731 133 2765
rect 167 2731 205 2765
rect 239 2731 300 2765
rect 0 2669 300 2731
rect 0 2635 61 2669
rect 95 2635 133 2669
rect 167 2635 205 2669
rect 239 2635 300 2669
rect 0 2573 300 2635
rect 0 2539 61 2573
rect 95 2539 133 2573
rect 167 2539 205 2573
rect 239 2539 300 2573
rect 0 2477 300 2539
rect 0 2443 61 2477
rect 95 2443 133 2477
rect 167 2443 205 2477
rect 239 2443 300 2477
rect 0 2381 300 2443
rect 0 2347 61 2381
rect 95 2347 133 2381
rect 167 2347 205 2381
rect 239 2347 300 2381
rect 0 2285 300 2347
rect 0 2251 61 2285
rect 95 2251 133 2285
rect 167 2251 205 2285
rect 239 2251 300 2285
rect 0 2189 300 2251
rect 0 2155 61 2189
rect 95 2155 133 2189
rect 167 2155 205 2189
rect 239 2155 300 2189
rect 0 2093 300 2155
rect 0 2059 61 2093
rect 95 2059 133 2093
rect 167 2059 205 2093
rect 239 2059 300 2093
rect 0 1997 300 2059
rect 0 1963 61 1997
rect 95 1963 133 1997
rect 167 1963 205 1997
rect 239 1963 300 1997
rect 0 1901 300 1963
rect 0 1867 61 1901
rect 95 1867 133 1901
rect 167 1867 205 1901
rect 239 1867 300 1901
rect 0 1805 300 1867
rect 0 1771 61 1805
rect 95 1771 133 1805
rect 167 1771 205 1805
rect 239 1771 300 1805
rect 0 1709 300 1771
rect 0 1675 61 1709
rect 95 1675 133 1709
rect 167 1675 205 1709
rect 239 1675 300 1709
rect 0 1613 300 1675
rect 0 1579 61 1613
rect 95 1579 133 1613
rect 167 1579 205 1613
rect 239 1579 300 1613
rect 0 1517 300 1579
rect 0 1483 61 1517
rect 95 1483 133 1517
rect 167 1483 205 1517
rect 239 1483 300 1517
rect 0 1421 300 1483
rect 0 1387 61 1421
rect 95 1387 133 1421
rect 167 1387 205 1421
rect 239 1387 300 1421
rect 0 1325 300 1387
rect 0 1291 61 1325
rect 95 1291 133 1325
rect 167 1291 205 1325
rect 239 1291 300 1325
rect 0 1229 300 1291
rect 0 1195 61 1229
rect 95 1195 133 1229
rect 167 1195 205 1229
rect 239 1195 300 1229
rect 0 1133 300 1195
rect 0 1099 61 1133
rect 95 1099 133 1133
rect 167 1099 205 1133
rect 239 1099 300 1133
rect 0 1037 300 1099
rect 0 1003 61 1037
rect 95 1003 133 1037
rect 167 1003 205 1037
rect 239 1003 300 1037
rect 0 941 300 1003
rect 0 907 61 941
rect 95 907 133 941
rect 167 907 205 941
rect 239 907 300 941
rect 0 845 300 907
rect 0 811 61 845
rect 95 811 133 845
rect 167 811 205 845
rect 239 811 300 845
rect 0 749 300 811
rect 0 715 61 749
rect 95 715 133 749
rect 167 715 205 749
rect 239 715 300 749
rect 0 653 300 715
rect 0 619 61 653
rect 95 619 133 653
rect 167 619 205 653
rect 239 619 300 653
rect 0 557 300 619
rect 0 523 61 557
rect 95 523 133 557
rect 167 523 205 557
rect 239 523 300 557
rect 0 461 300 523
rect 0 427 61 461
rect 95 427 133 461
rect 167 427 205 461
rect 239 427 300 461
rect 0 365 300 427
rect 0 331 61 365
rect 95 331 133 365
rect 167 331 205 365
rect 239 331 300 365
rect 0 269 300 331
rect 0 235 61 269
rect 95 235 133 269
rect 167 235 205 269
rect 239 235 300 269
rect 0 173 300 235
rect 0 139 61 173
rect 95 139 133 173
rect 167 139 205 173
rect 239 139 300 173
rect 0 60 300 139
tri 0 0 60 60 ne
rect 60 0 240 60
tri 240 0 300 60 nw
use sky130_fd_pr__via_l1m1__example_55959141808683  sky130_fd_pr__via_l1m1__example_55959141808683_0
timestamp 1619729480
transform 1 0 61 0 1 139
box 0 0 1 1
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 9282696
string GDS_START 9269598
<< end >>
