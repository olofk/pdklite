magic
tech sky130A
magscale 1 2
timestamp 1640697850
<< nwell >>
rect 10462 3498 10993 4199
rect 11779 3498 11790 4199
rect 12214 3498 12495 4199
<< locali >>
rect 18233 5175 18284 5209
rect 18318 5175 18369 5209
rect 18199 5137 18403 5175
rect 18233 5103 18284 5137
rect 18318 5103 18369 5137
rect 18199 5065 18403 5103
rect 18233 5031 18284 5065
rect 18318 5031 18369 5065
rect 11176 4232 11242 4282
rect 11176 4198 11194 4232
rect 11228 4198 11242 4232
rect 11278 4263 11312 4301
rect 11527 4301 11540 4335
rect 11574 4301 11593 4335
rect 11527 4282 11593 4301
rect 11347 4236 11413 4282
rect 11176 4160 11242 4198
rect 11176 4126 11194 4160
rect 11228 4126 11242 4160
rect 11347 4202 11366 4236
rect 11400 4202 11413 4236
rect 11540 4263 11574 4282
rect 11347 4164 11413 4202
rect 11630 4198 11664 4236
rect 11779 4248 11824 4282
rect 11745 4210 11824 4248
rect 11779 4180 11824 4210
rect 11930 4226 11964 4264
rect 12011 4210 12045 4248
rect 11347 4130 11366 4164
rect 11400 4130 11413 4164
rect 11176 4074 11242 4126
<< viali >>
rect 18199 5175 18233 5209
rect 18284 5175 18318 5209
rect 18369 5175 18403 5209
rect 18199 5103 18233 5137
rect 18284 5103 18318 5137
rect 18369 5103 18403 5137
rect 18199 5031 18233 5065
rect 18284 5031 18318 5065
rect 18369 5031 18403 5065
rect 11278 4301 11312 4335
rect 11194 4198 11228 4232
rect 11540 4301 11574 4335
rect 11278 4229 11312 4263
rect 11194 4126 11228 4160
rect 11366 4202 11400 4236
rect 11540 4229 11574 4263
rect 11630 4236 11664 4270
rect 11630 4164 11664 4198
rect 11745 4248 11779 4282
rect 11745 4176 11779 4210
rect 11930 4264 11964 4298
rect 11930 4192 11964 4226
rect 12011 4248 12045 4282
rect 12011 4176 12045 4210
rect 11366 4130 11400 4164
<< metal1 >>
rect 10272 11325 10278 11377
rect 10330 11325 10342 11377
rect 10394 11368 14010 11377
tri 14010 11368 14019 11377 sw
rect 10394 11325 14019 11368
tri 14019 11325 14062 11368 sw
tri 13988 11294 14019 11325 ne
rect 14019 11294 14062 11325
tri 14062 11294 14093 11325 sw
tri 14019 11242 14071 11294 ne
rect 14071 11242 15625 11294
rect 15677 11242 15689 11294
rect 15741 11242 15747 11294
rect 8965 6643 8993 6843
rect 17224 6642 17267 6843
rect 11548 6607 11600 6613
rect 11548 6543 11600 6555
tri 11600 6531 11631 6562 nw
rect 11548 6485 11600 6491
rect 3549 6232 3589 6303
rect 3902 6296 3984 6332
rect 8965 5947 8993 6145
rect 17224 5946 17267 6145
rect 8965 5178 8993 5308
rect 16748 5302 16791 5308
rect 16747 5179 16791 5302
rect 16748 5178 16791 5179
rect 18187 5214 18415 5215
rect 18187 5162 18193 5214
rect 18245 5162 18275 5214
rect 18327 5162 18357 5214
rect 18409 5162 18415 5214
rect 8965 4948 8993 5150
rect 16747 4948 16790 5150
rect 18187 5146 18415 5162
rect 18187 5094 18193 5146
rect 18245 5094 18275 5146
rect 18327 5094 18357 5146
rect 18409 5094 18415 5146
rect 18187 5078 18415 5094
rect 18187 5026 18193 5078
rect 18245 5026 18275 5078
rect 18327 5026 18357 5078
rect 18409 5026 18415 5078
rect 18187 5025 18415 5026
rect 11054 4867 11060 4919
rect 11112 4867 11124 4919
rect 11176 4867 11714 4919
rect 11766 4867 11778 4919
rect 11830 4867 11878 4919
rect 4690 4793 4762 4826
rect 11714 4783 11720 4835
rect 11772 4783 11784 4835
rect 11836 4783 11842 4835
rect 14230 4783 14236 4835
rect 14288 4783 14300 4835
rect 14352 4783 14358 4835
rect 7178 4703 7184 4755
rect 7236 4703 7248 4755
rect 7300 4703 7306 4755
rect 11719 4375 11742 4590
rect 11088 4339 11140 4345
tri 10534 4275 10536 4277 se
rect 4734 4217 4764 4275
tri 10531 4272 10534 4275 se
rect 10534 4272 10536 4275
rect 9684 4215 9736 4221
rect 9889 4208 9931 4265
rect 10066 4205 10092 4268
rect 10103 4208 10536 4272
rect 11088 4275 11140 4287
rect 11272 4335 11318 4347
tri 11318 4335 11330 4347 sw
tri 11522 4335 11534 4347 se
rect 11534 4335 11580 4347
rect 11272 4301 11278 4335
rect 11312 4319 11330 4335
tri 11330 4319 11346 4335 sw
tri 11506 4319 11522 4335 se
rect 11522 4319 11540 4335
rect 11312 4301 11540 4319
rect 11574 4301 11580 4335
rect 11272 4291 11580 4301
rect 11915 4304 11970 4310
rect 11272 4282 11347 4291
tri 11347 4282 11356 4291 nw
tri 11485 4282 11494 4291 ne
rect 11494 4282 11580 4291
rect 11739 4282 11785 4294
rect 11272 4270 11335 4282
tri 11335 4270 11347 4282 nw
tri 11494 4270 11506 4282 ne
rect 11506 4270 11580 4282
rect 11272 4263 11328 4270
tri 11328 4263 11335 4270 nw
tri 11506 4263 11513 4270 ne
rect 11513 4263 11580 4270
rect 10103 4205 10143 4208
tri 10143 4205 10146 4208 nw
tri 10493 4205 10496 4208 ne
rect 10496 4205 10536 4208
rect 10103 4198 10136 4205
tri 10136 4198 10143 4205 nw
tri 10496 4198 10503 4205 ne
rect 10503 4198 10536 4205
tri 11075 4198 11088 4211 se
rect 11088 4198 11140 4223
tri 10103 4165 10136 4198 nw
tri 10503 4165 10536 4198 ne
tri 11060 4183 11075 4198 se
rect 11075 4189 11140 4198
rect 11075 4183 11134 4189
tri 11134 4183 11140 4189 nw
rect 11182 4232 11234 4244
rect 11272 4229 11278 4263
rect 11312 4229 11318 4263
tri 11318 4253 11328 4263 nw
tri 11513 4253 11523 4263 ne
rect 11523 4253 11540 4263
tri 11523 4248 11528 4253 ne
rect 11528 4248 11540 4253
rect 11272 4217 11318 4229
rect 11357 4242 11409 4248
tri 11528 4242 11534 4248 ne
tri 10763 4165 10781 4183 se
rect 10781 4165 11115 4183
tri 10762 4164 10763 4165 se
rect 10763 4164 11115 4165
tri 11115 4164 11134 4183 nw
rect 11182 4168 11234 4180
rect 9684 4146 9736 4163
tri 10758 4160 10762 4164 se
rect 10762 4160 11111 4164
tri 11111 4160 11115 4164 nw
rect 5203 4097 5307 4129
tri 5443 4083 5449 4089 ne
rect 5449 4083 5455 4135
rect 5507 4083 5519 4135
rect 5571 4083 5577 4135
rect 7194 4083 7200 4135
rect 7252 4083 7264 4135
rect 7316 4129 7322 4135
rect 7316 4096 7344 4129
rect 7316 4083 7322 4096
rect 9433 4083 9439 4135
rect 9491 4083 9503 4135
rect 9555 4083 9561 4135
tri 10738 4140 10758 4160 se
rect 10758 4142 11093 4160
tri 11093 4142 11111 4160 nw
rect 10758 4140 10786 4142
tri 9736 4126 9750 4140 sw
tri 10724 4126 10738 4140 se
rect 10738 4126 10786 4140
tri 10786 4126 10802 4142 nw
rect 9736 4121 9750 4126
tri 9750 4121 9755 4126 sw
tri 10719 4121 10724 4126 se
rect 10724 4121 10781 4126
tri 10781 4121 10786 4126 nw
rect 9736 4114 9755 4121
tri 9755 4114 9762 4121 sw
tri 10712 4114 10719 4121 se
rect 10719 4114 10774 4121
tri 10774 4114 10781 4121 nw
rect 11534 4229 11540 4248
rect 11574 4229 11580 4263
rect 11534 4217 11580 4229
rect 11622 4276 11674 4282
rect 11357 4176 11409 4190
rect 11622 4210 11674 4224
rect 11739 4248 11745 4282
rect 11779 4248 11785 4282
rect 11739 4210 11785 4248
rect 11739 4176 11745 4210
rect 11779 4176 11785 4210
rect 11967 4252 11970 4304
rect 11915 4238 11970 4252
rect 11967 4186 11970 4238
rect 11915 4180 11970 4186
rect 12002 4288 12054 4294
rect 12002 4222 12054 4236
rect 11622 4152 11674 4158
tri 11728 4152 11739 4163 se
rect 11739 4152 11785 4176
rect 12002 4164 12054 4170
tri 11722 4146 11728 4152 se
rect 11728 4146 11785 4152
rect 11357 4118 11409 4124
tri 11694 4118 11722 4146 se
rect 11722 4143 11785 4146
rect 11722 4118 11739 4143
rect 9736 4110 10770 4114
tri 10770 4110 10774 4114 nw
rect 11182 4110 11234 4116
tri 11686 4110 11694 4118 se
rect 11694 4110 11739 4118
rect 9736 4094 10748 4110
rect 9684 4088 10748 4094
tri 10748 4088 10770 4110 nw
tri 11677 4101 11686 4110 se
rect 11686 4101 11739 4110
rect 9684 4086 10746 4088
tri 10746 4086 10748 4088 nw
rect 11000 4049 11006 4101
rect 11058 4049 11070 4101
rect 11122 4097 11128 4101
tri 11128 4097 11132 4101 sw
tri 11673 4097 11677 4101 se
rect 11677 4097 11739 4101
tri 11739 4097 11785 4143 nw
rect 13615 4140 13667 4146
rect 11122 4091 11132 4097
tri 11132 4091 11138 4097 sw
tri 11667 4091 11673 4097 se
rect 11673 4091 11733 4097
tri 11733 4091 11739 4097 nw
rect 11122 4088 11138 4091
tri 11138 4088 11141 4091 sw
tri 11664 4088 11667 4091 se
rect 11667 4088 11730 4091
tri 11730 4088 11733 4091 nw
tri 13612 4088 13615 4091 se
rect 11122 4086 11141 4088
tri 11141 4086 11143 4088 sw
tri 11662 4086 11664 4088 se
rect 11664 4086 11728 4088
tri 11728 4086 11730 4088 nw
tri 13610 4086 13612 4088 se
rect 13612 4086 13667 4088
rect 11122 4083 11143 4086
tri 11143 4083 11146 4086 sw
tri 11659 4083 11662 4086 se
rect 11662 4083 11725 4086
tri 11725 4083 11728 4086 nw
tri 13607 4083 13610 4086 se
rect 13610 4083 13667 4086
rect 11122 4077 11146 4083
tri 11146 4077 11152 4083 sw
tri 11653 4077 11659 4083 se
rect 11659 4077 11719 4083
tri 11719 4077 11725 4083 nw
tri 13601 4077 13607 4083 se
rect 13607 4077 13667 4083
rect 11122 4070 11712 4077
tri 11712 4070 11719 4077 nw
tri 13594 4070 13601 4077 se
rect 13601 4076 13667 4077
rect 13601 4070 13615 4076
rect 11122 4049 11691 4070
tri 11691 4049 11712 4070 nw
rect 12193 4018 12199 4070
rect 12251 4018 12263 4070
rect 12315 4057 12321 4070
tri 12321 4057 12334 4070 sw
tri 13581 4057 13594 4070 se
rect 13594 4057 13615 4070
rect 12315 4024 13615 4057
rect 12315 4018 13667 4024
rect 16703 3997 16780 4029
rect 9302 3797 9308 3849
rect 9360 3797 9372 3849
rect 9424 3797 9430 3849
rect 9458 3798 9464 3850
rect 9516 3798 9528 3850
rect 9580 3798 9965 3850
rect 10017 3798 10029 3850
rect 10081 3798 10087 3850
rect 10596 3808 10602 3860
rect 10654 3808 10666 3860
rect 10718 3808 11006 3860
rect 11058 3808 11070 3860
rect 11122 3808 11128 3860
rect 11602 3552 11645 3754
rect 11719 3552 11742 3755
rect 12152 3553 12523 3755
<< via1 >>
rect 10278 11325 10330 11377
rect 10342 11325 10394 11377
rect 15625 11242 15677 11294
rect 15689 11242 15741 11294
rect 11548 6555 11600 6607
rect 11548 6491 11600 6543
rect 18193 5209 18245 5214
rect 18193 5175 18199 5209
rect 18199 5175 18233 5209
rect 18233 5175 18245 5209
rect 18193 5162 18245 5175
rect 18275 5209 18327 5214
rect 18275 5175 18284 5209
rect 18284 5175 18318 5209
rect 18318 5175 18327 5209
rect 18275 5162 18327 5175
rect 18357 5209 18409 5214
rect 18357 5175 18369 5209
rect 18369 5175 18403 5209
rect 18403 5175 18409 5209
rect 18357 5162 18409 5175
rect 18193 5137 18245 5146
rect 18193 5103 18199 5137
rect 18199 5103 18233 5137
rect 18233 5103 18245 5137
rect 18193 5094 18245 5103
rect 18275 5137 18327 5146
rect 18275 5103 18284 5137
rect 18284 5103 18318 5137
rect 18318 5103 18327 5137
rect 18275 5094 18327 5103
rect 18357 5137 18409 5146
rect 18357 5103 18369 5137
rect 18369 5103 18403 5137
rect 18403 5103 18409 5137
rect 18357 5094 18409 5103
rect 18193 5065 18245 5078
rect 18193 5031 18199 5065
rect 18199 5031 18233 5065
rect 18233 5031 18245 5065
rect 18193 5026 18245 5031
rect 18275 5065 18327 5078
rect 18275 5031 18284 5065
rect 18284 5031 18318 5065
rect 18318 5031 18327 5065
rect 18275 5026 18327 5031
rect 18357 5065 18409 5078
rect 18357 5031 18369 5065
rect 18369 5031 18403 5065
rect 18403 5031 18409 5065
rect 18357 5026 18409 5031
rect 11060 4867 11112 4919
rect 11124 4867 11176 4919
rect 11714 4867 11766 4919
rect 11778 4867 11830 4919
rect 11720 4783 11772 4835
rect 11784 4783 11836 4835
rect 14236 4783 14288 4835
rect 14300 4783 14352 4835
rect 7184 4703 7236 4755
rect 7248 4703 7300 4755
rect 11088 4287 11140 4339
rect 9684 4163 9736 4215
rect 11088 4223 11140 4275
rect 11915 4298 11967 4304
rect 11182 4198 11194 4232
rect 11194 4198 11228 4232
rect 11228 4198 11234 4232
rect 11357 4236 11409 4242
rect 11182 4180 11234 4198
rect 11182 4160 11234 4168
rect 5455 4083 5507 4135
rect 5519 4083 5571 4135
rect 7200 4083 7252 4135
rect 7264 4083 7316 4135
rect 9439 4083 9491 4135
rect 9503 4083 9555 4135
rect 9684 4094 9736 4146
rect 11182 4126 11194 4160
rect 11194 4126 11228 4160
rect 11228 4126 11234 4160
rect 11182 4116 11234 4126
rect 11357 4202 11366 4236
rect 11366 4202 11400 4236
rect 11400 4202 11409 4236
rect 11622 4270 11674 4276
rect 11622 4236 11630 4270
rect 11630 4236 11664 4270
rect 11664 4236 11674 4270
rect 11622 4224 11674 4236
rect 11357 4190 11409 4202
rect 11357 4164 11409 4176
rect 11357 4130 11366 4164
rect 11366 4130 11400 4164
rect 11400 4130 11409 4164
rect 11622 4198 11674 4210
rect 11622 4164 11630 4198
rect 11630 4164 11664 4198
rect 11664 4164 11674 4198
rect 11622 4158 11674 4164
rect 11915 4264 11930 4298
rect 11930 4264 11964 4298
rect 11964 4264 11967 4298
rect 11915 4252 11967 4264
rect 11915 4226 11967 4238
rect 11915 4192 11930 4226
rect 11930 4192 11964 4226
rect 11964 4192 11967 4226
rect 11915 4186 11967 4192
rect 12002 4282 12054 4288
rect 12002 4248 12011 4282
rect 12011 4248 12045 4282
rect 12045 4248 12054 4282
rect 12002 4236 12054 4248
rect 12002 4210 12054 4222
rect 12002 4176 12011 4210
rect 12011 4176 12045 4210
rect 12045 4176 12054 4210
rect 12002 4170 12054 4176
rect 11357 4124 11409 4130
rect 11006 4049 11058 4101
rect 11070 4049 11122 4101
rect 13615 4088 13667 4140
rect 12199 4018 12251 4070
rect 12263 4018 12315 4070
rect 13615 4024 13667 4076
rect 9308 3797 9360 3849
rect 9372 3797 9424 3849
rect 9464 3798 9516 3850
rect 9528 3798 9580 3850
rect 9965 3798 10017 3850
rect 10029 3798 10081 3850
rect 10602 3808 10654 3860
rect 10666 3808 10718 3860
rect 11006 3808 11058 3860
rect 11070 3808 11122 3860
<< metal2 >>
rect 10272 11325 10278 11377
rect 10330 11325 10342 11377
rect 10394 11325 10400 11377
rect 10272 11294 10334 11325
tri 10334 11294 10365 11325 nw
tri 10198 6972 10272 7046 se
rect 10272 7024 10324 11294
tri 10324 11284 10334 11294 nw
rect 15619 11242 15625 11294
rect 15677 11242 15689 11294
rect 15741 11242 15747 11294
tri 15665 11200 15707 11242 ne
rect 15707 11008 15747 11242
tri 15707 10983 15732 11008 ne
rect 15732 10983 15747 11008
tri 15747 10983 15790 11026 sw
tri 15732 10968 15747 10983 ne
rect 15747 10968 15790 10983
tri 15747 10925 15790 10968 ne
tri 15790 10925 15848 10983 sw
tri 15790 10867 15848 10925 ne
tri 15848 10867 15906 10925 sw
tri 15848 10849 15866 10867 ne
rect 15866 8684 15906 10867
tri 15906 8684 15922 8700 sw
rect 15866 8682 15922 8684
tri 15866 8626 15922 8682 ne
tri 15922 8626 15980 8684 sw
tri 15922 8568 15980 8626 ne
tri 15980 8568 16038 8626 sw
tri 15980 8550 15998 8568 ne
tri 10272 6972 10324 7024 nw
tri 10186 6960 10198 6972 se
rect 10198 6960 10260 6972
tri 10260 6960 10272 6972 nw
rect 6382 6791 6434 6843
rect 6476 6791 6528 6843
tri 10112 6037 10186 6111 se
rect 10186 6089 10238 6960
tri 10238 6938 10260 6960 nw
rect 10622 6791 10674 6843
rect 10716 6791 10768 6843
rect 11316 6791 11368 6843
rect 14776 6791 14828 6843
rect 14870 6791 14922 6843
rect 15470 6791 15522 6843
rect 15564 6791 15616 6843
rect 15998 6775 16038 8568
tri 15998 6744 16029 6775 ne
rect 16029 6744 16038 6775
tri 16038 6744 16087 6793 sw
tri 16029 6735 16038 6744 ne
rect 16038 6735 16840 6744
tri 16038 6704 16069 6735 ne
rect 16069 6704 16840 6735
tri 10186 6037 10238 6089 nw
rect 11548 6607 11600 6613
rect 11548 6543 11600 6555
tri 10077 6002 10112 6037 se
rect 10112 6002 10151 6037
tri 10151 6002 10186 6037 nw
rect 10077 5146 10129 6002
tri 10129 5980 10151 6002 nw
tri 10129 5146 10132 5149 sw
rect 10077 5127 10132 5146
tri 10132 5127 10151 5146 sw
tri 10077 5094 10110 5127 ne
rect 10110 5094 10151 5127
tri 10151 5094 10184 5127 sw
tri 10110 5078 10126 5094 ne
rect 10126 5078 10184 5094
tri 10184 5078 10200 5094 sw
tri 10126 5053 10151 5078 ne
rect 10151 5075 10200 5078
tri 10200 5075 10203 5078 sw
rect 10151 5053 10203 5075
tri 10203 5053 10225 5075 sw
rect 11548 5053 11600 6491
rect 16114 6547 16123 6603
rect 16179 6547 16218 6603
rect 16274 6547 17233 6603
rect 16114 6523 17233 6547
rect 16114 6467 16123 6523
rect 16179 6467 16218 6523
rect 16274 6467 17233 6523
tri 17233 6467 17369 6603 sw
tri 17137 6456 17148 6467 ne
rect 17148 6456 17369 6467
tri 17369 6456 17380 6467 sw
tri 17148 6372 17232 6456 ne
tri 17135 5705 17232 5802 se
rect 17232 5740 17380 6456
rect 17232 5705 17345 5740
tri 17345 5705 17380 5740 nw
tri 11600 5053 11610 5063 sw
tri 10151 5026 10178 5053 ne
rect 10178 5026 10225 5053
tri 10225 5026 10252 5053 sw
rect 11548 5041 11610 5053
tri 11610 5041 11622 5053 sw
tri 11548 5026 11563 5041 ne
rect 11563 5026 11622 5041
tri 11622 5026 11637 5041 sw
tri 10178 5001 10203 5026 ne
rect 10203 5023 10252 5026
tri 10252 5023 10255 5026 sw
rect 5193 4854 5245 4906
rect 9346 4854 9398 4906
tri 10173 4783 10203 4813 se
rect 10203 4791 10255 5023
tri 11563 4967 11622 5026 ne
rect 11622 4989 11637 5026
tri 11637 4989 11674 5026 sw
rect 11054 4867 11060 4919
rect 11112 4867 11124 4919
rect 11176 4867 11182 4919
tri 11054 4835 11086 4867 ne
rect 11086 4835 11150 4867
tri 11150 4835 11182 4867 nw
tri 11086 4833 11088 4835 ne
rect 11088 4833 11148 4835
tri 11148 4833 11150 4835 nw
rect 10203 4783 10247 4791
tri 10247 4783 10255 4791 nw
rect 5488 4755 5542 4783
tri 5542 4755 5570 4783 nw
tri 10145 4755 10173 4783 se
rect 10173 4755 10203 4783
tri 5486 4172 5488 4174 se
rect 5488 4172 5540 4755
tri 5540 4753 5542 4755 nw
rect 7178 4703 7184 4755
rect 7236 4703 7248 4755
rect 7300 4703 7306 4755
tri 10129 4739 10145 4755 se
rect 10145 4739 10203 4755
tri 10203 4739 10247 4783 nw
tri 10093 4703 10129 4739 se
tri 7178 4679 7202 4703 ne
rect 7202 4679 7306 4703
tri 7202 4660 7221 4679 ne
rect 7221 4665 7292 4679
tri 7292 4665 7306 4679 nw
tri 10055 4665 10093 4703 se
rect 10093 4665 10129 4703
tri 10129 4665 10203 4739 nw
rect 7221 4172 7273 4665
tri 7273 4646 7292 4665 nw
tri 10036 4646 10055 4665 se
tri 9981 4591 10036 4646 se
rect 10036 4591 10055 4646
tri 10055 4591 10129 4665 nw
tri 9975 4585 9981 4591 se
rect 9981 4585 10049 4591
tri 10049 4585 10055 4591 nw
tri 9415 4287 9425 4297 se
rect 9425 4287 9625 4297
tri 9625 4287 9635 4297 sw
tri 9404 4276 9415 4287 se
rect 9415 4276 9635 4287
tri 9635 4276 9646 4287 sw
tri 9403 4275 9404 4276 se
rect 9404 4275 9646 4276
tri 9646 4275 9647 4276 sw
tri 9388 4260 9403 4275 se
rect 9403 4260 9647 4275
tri 9647 4260 9662 4275 sw
tri 9351 4223 9388 4260 se
rect 9388 4245 9662 4260
rect 9388 4223 9425 4245
tri 9425 4223 9447 4245 nw
tri 9603 4223 9625 4245 ne
rect 9625 4223 9662 4245
tri 9662 4223 9699 4260 sw
tri 9343 4215 9351 4223 se
rect 9351 4215 9417 4223
tri 9417 4215 9425 4223 nw
tri 9625 4215 9633 4223 ne
rect 9633 4221 9699 4223
tri 9699 4221 9701 4223 sw
rect 9633 4215 9736 4221
tri 9321 4193 9343 4215 se
rect 9343 4193 9395 4215
tri 9395 4193 9417 4215 nw
tri 9633 4193 9655 4215 ne
rect 9655 4193 9684 4215
rect 9321 4186 9388 4193
tri 9388 4186 9395 4193 nw
tri 9655 4186 9662 4193 ne
rect 9662 4186 9684 4193
rect 9321 4184 9386 4186
tri 9386 4184 9388 4186 nw
tri 9662 4184 9664 4186 ne
rect 9664 4184 9684 4186
tri 7273 4172 7285 4184 sw
rect 9321 4172 9374 4184
tri 9374 4172 9386 4184 nw
tri 9664 4172 9676 4184 ne
rect 9676 4172 9684 4184
tri 5477 4163 5486 4172 se
rect 5486 4163 5540 4172
tri 5540 4163 5549 4172 sw
rect 7221 4163 7285 4172
tri 7285 4163 7294 4172 sw
tri 5460 4146 5477 4163 se
rect 5477 4146 5549 4163
tri 5549 4146 5566 4163 sw
tri 7205 4146 7221 4162 se
rect 7221 4146 7294 4163
tri 7294 4146 7311 4163 sw
tri 5449 4135 5460 4146 se
rect 5460 4135 5566 4146
tri 5566 4135 5577 4146 sw
rect 5449 4083 5455 4135
rect 5507 4083 5519 4135
rect 5571 4083 5577 4135
tri 7194 4135 7205 4146 se
rect 7205 4135 7311 4146
tri 7311 4135 7322 4146 sw
rect 7194 4083 7200 4135
rect 7252 4083 7264 4135
rect 7316 4083 7322 4135
rect 8837 3843 8865 3867
rect 9321 3849 9373 4172
tri 9373 4171 9374 4172 nw
tri 9676 4171 9677 4172 ne
rect 9677 4171 9684 4172
tri 9677 4164 9684 4171 ne
rect 9684 4146 9736 4163
rect 9433 4083 9439 4135
rect 9491 4083 9503 4135
rect 9555 4083 9561 4135
rect 9684 4086 9736 4094
rect 9433 4023 9561 4083
tri 9561 4023 9586 4048 sw
rect 9433 4018 9586 4023
tri 9433 4015 9436 4018 ne
rect 9436 4015 9586 4018
tri 9436 3993 9458 4015 ne
rect 9458 3850 9586 4015
rect 9302 3797 9308 3849
rect 9360 3797 9372 3849
rect 9424 3797 9430 3849
rect 9458 3798 9464 3850
rect 9516 3798 9528 3850
rect 9580 3798 9586 3850
tri 9959 3872 9975 3888 se
rect 9975 3872 10027 4585
tri 10027 4563 10049 4585 nw
rect 11088 4345 11140 4833
tri 11140 4825 11148 4833 nw
tri 11140 4345 11216 4421 sw
rect 11088 4339 11286 4345
rect 11140 4322 11286 4339
tri 11286 4322 11309 4345 sw
rect 11140 4304 11309 4322
tri 11309 4304 11327 4322 sw
rect 11140 4294 11327 4304
tri 11327 4294 11337 4304 sw
rect 11140 4293 11337 4294
rect 11140 4287 11161 4293
rect 11088 4276 11161 4287
tri 11161 4276 11178 4293 nw
tri 11264 4276 11281 4293 ne
rect 11281 4276 11337 4293
tri 11337 4276 11355 4294 sw
rect 11622 4276 11674 4989
rect 11708 4867 11714 4919
rect 11766 4867 11778 4919
rect 11830 4905 11871 4919
tri 11871 4905 11885 4919 sw
rect 11830 4867 11885 4905
tri 11851 4835 11883 4867 ne
rect 11883 4835 11885 4867
tri 11885 4835 11955 4905 sw
rect 12675 4854 12727 4906
rect 13475 4854 13527 4906
rect 11714 4783 11720 4835
rect 11772 4783 11784 4835
rect 11836 4783 11842 4835
tri 11883 4833 11885 4835 ne
rect 11885 4833 11955 4835
tri 11955 4833 11957 4835 sw
tri 14083 4833 14085 4835 se
rect 14085 4833 14236 4835
tri 11885 4783 11935 4833 ne
rect 11935 4783 11957 4833
tri 11957 4783 12007 4833 sw
tri 14033 4783 14083 4833 se
rect 14083 4783 14236 4833
rect 14288 4783 14300 4835
rect 14352 4783 14358 4835
tri 11728 4754 11757 4783 ne
rect 11757 4761 11820 4783
tri 11820 4761 11842 4783 nw
tri 11935 4761 11957 4783 ne
rect 11957 4761 12007 4783
tri 12007 4761 12029 4783 sw
tri 14011 4761 14033 4783 se
rect 14033 4761 14063 4783
rect 11757 4545 11809 4761
tri 11809 4750 11820 4761 nw
tri 11957 4750 11968 4761 ne
rect 11968 4750 12029 4761
tri 11968 4739 11979 4750 ne
rect 11979 4739 12029 4750
tri 12029 4739 12051 4761 sw
tri 13989 4739 14011 4761 se
rect 14011 4739 14063 4761
tri 14063 4739 14107 4783 nw
tri 11979 4689 12029 4739 ne
rect 12029 4713 12051 4739
tri 12051 4713 12077 4739 sw
tri 13963 4713 13989 4739 se
rect 13989 4713 14037 4739
tri 14037 4713 14063 4739 nw
rect 12029 4689 12077 4713
tri 12077 4689 12101 4713 sw
tri 13939 4689 13963 4713 se
rect 13963 4689 13989 4713
tri 12029 4665 12053 4689 ne
rect 12053 4665 12101 4689
tri 12101 4665 12125 4689 sw
tri 13915 4665 13939 4689 se
rect 13939 4665 13989 4689
tri 13989 4665 14037 4713 nw
rect 17135 4681 17283 5705
tri 17283 5643 17345 5705 nw
rect 18187 5214 18415 5215
rect 18187 5162 18193 5214
rect 18245 5162 18275 5214
rect 18327 5162 18357 5214
rect 18409 5162 18415 5214
rect 18187 5146 18415 5162
rect 18187 5094 18193 5146
rect 18245 5094 18275 5146
rect 18327 5094 18357 5146
rect 18409 5094 18415 5146
rect 18187 5078 18415 5094
rect 18187 5026 18193 5078
rect 18245 5026 18275 5078
rect 18327 5026 18357 5078
rect 18409 5026 18415 5078
tri 18131 4835 18187 4891 se
rect 18187 4835 18415 5026
tri 18051 4755 18131 4835 se
rect 18131 4755 18335 4835
tri 18335 4755 18415 4835 nw
tri 17999 4703 18051 4755 se
rect 18051 4703 18283 4755
tri 18283 4703 18335 4755 nw
tri 17998 4702 17999 4703 se
rect 17999 4702 18220 4703
tri 17283 4681 17304 4702 sw
tri 17977 4681 17998 4702 se
rect 17998 4681 18220 4702
tri 12053 4617 12101 4665 ne
rect 12101 4639 12125 4665
tri 12125 4639 12151 4665 sw
tri 13889 4639 13915 4665 se
rect 13915 4639 13963 4665
tri 13963 4639 13989 4665 nw
rect 17135 4640 17304 4681
tri 17304 4640 17345 4681 sw
tri 17936 4640 17977 4681 se
rect 17977 4640 18220 4681
tri 18220 4640 18283 4703 nw
tri 17135 4639 17136 4640 ne
rect 17136 4639 17345 4640
rect 12101 4617 12151 4639
tri 12151 4617 12173 4639 sw
tri 13867 4617 13889 4639 se
rect 13889 4617 13915 4639
tri 12101 4591 12127 4617 ne
rect 12127 4591 12173 4617
tri 12173 4591 12199 4617 sw
tri 13841 4591 13867 4617 se
rect 13867 4591 13915 4617
tri 13915 4591 13963 4639 nw
tri 17136 4591 17184 4639 ne
rect 17184 4619 17345 4639
tri 17345 4619 17366 4640 sw
tri 17915 4619 17936 4640 se
rect 17936 4619 18051 4640
rect 17184 4591 18051 4619
tri 12127 4585 12133 4591 ne
rect 12133 4585 12199 4591
tri 12199 4585 12205 4591 sw
tri 13835 4585 13841 4591 se
rect 13841 4585 13909 4591
tri 13909 4585 13915 4591 nw
tri 17184 4585 17190 4591 ne
rect 17190 4585 18051 4591
tri 12133 4563 12155 4585 ne
rect 12155 4565 12205 4585
tri 12205 4565 12225 4585 sw
tri 13815 4565 13835 4585 se
rect 13835 4565 13889 4585
tri 13889 4565 13909 4585 nw
tri 17190 4565 17210 4585 ne
rect 17210 4565 18051 4585
rect 12155 4563 12225 4565
tri 12225 4563 12227 4565 sw
tri 13813 4563 13815 4565 se
rect 13815 4563 13887 4565
tri 13887 4563 13889 4565 nw
tri 17210 4563 17212 4565 ne
rect 17212 4563 18051 4565
tri 12155 4548 12170 4563 ne
rect 12170 4548 12227 4563
tri 11809 4545 11812 4548 sw
tri 12170 4545 12173 4548 ne
rect 12173 4545 12227 4548
tri 12227 4545 12245 4563 sw
rect 11757 4538 11812 4545
tri 11812 4538 11819 4545 sw
tri 12173 4538 12180 4545 ne
rect 12180 4538 12245 4545
rect 11757 4526 11819 4538
tri 11757 4464 11819 4526 ne
tri 11819 4525 11832 4538 sw
tri 12180 4525 12193 4538 ne
rect 11819 4464 11832 4525
tri 11832 4464 11893 4525 sw
tri 11819 4421 11862 4464 ne
rect 11862 4421 11893 4464
tri 11893 4421 11936 4464 sw
tri 11862 4390 11893 4421 ne
rect 11893 4390 11936 4421
tri 11936 4390 11967 4421 sw
tri 11893 4368 11915 4390 ne
rect 11088 4275 11140 4276
tri 11140 4255 11161 4276 nw
tri 11281 4255 11302 4276 ne
rect 11302 4255 11355 4276
tri 11302 4248 11309 4255 ne
rect 11309 4248 11355 4255
tri 11355 4248 11383 4276 sw
tri 11309 4242 11315 4248 ne
rect 11315 4242 11409 4248
tri 11315 4238 11319 4242 ne
rect 11319 4238 11357 4242
rect 11088 4217 11140 4223
rect 11182 4232 11234 4238
tri 11319 4217 11340 4238 ne
rect 11340 4217 11357 4238
tri 11340 4200 11357 4217 ne
rect 11182 4168 11234 4180
rect 11357 4176 11409 4190
rect 11622 4210 11674 4224
rect 11915 4304 11967 4390
rect 11915 4238 11967 4252
rect 11915 4180 11967 4186
rect 12002 4288 12054 4294
rect 12002 4222 12054 4236
rect 11622 4146 11674 4158
rect 11357 4118 11409 4124
rect 11000 4049 11006 4101
rect 11058 4049 11070 4101
rect 11122 4049 11128 4101
tri 11042 4018 11073 4049 ne
rect 11073 4018 11128 4049
tri 11073 4015 11076 4018 ne
tri 11040 3900 11076 3936 se
rect 11076 3900 11128 4018
tri 10648 3888 10660 3900 sw
tri 11028 3888 11040 3900 se
rect 11040 3888 11128 3900
tri 10027 3872 10043 3888 sw
rect 10648 3872 10660 3888
tri 10660 3872 10676 3888 sw
tri 11012 3872 11028 3888 se
rect 11028 3872 11128 3888
rect 9959 3860 10043 3872
tri 10043 3860 10055 3872 sw
rect 10648 3860 10676 3872
tri 10676 3860 10688 3872 sw
tri 11000 3860 11012 3872 se
rect 11012 3860 11128 3872
rect 9959 3850 10055 3860
tri 10055 3850 10065 3860 sw
rect 9959 3798 9965 3850
rect 10017 3798 10029 3850
rect 10081 3798 10087 3850
rect 10596 3808 10602 3860
rect 10654 3808 10666 3860
rect 10718 3808 10724 3860
rect 11000 3808 11006 3860
rect 11058 3808 11070 3860
rect 11122 3808 11128 3860
rect 10648 3798 10678 3808
tri 10678 3798 10688 3808 nw
rect 10648 3797 10677 3798
tri 10677 3797 10678 3798 nw
tri 10648 3768 10677 3797 nw
rect 11182 3725 11234 4116
tri 11928 3917 12002 3991 se
rect 12002 3969 12054 4170
rect 12193 4088 12245 4538
tri 13741 4491 13813 4563 se
rect 13813 4491 13815 4563
tri 13815 4491 13887 4563 nw
tri 17212 4491 17284 4563 ne
rect 17284 4491 18051 4563
tri 13667 4417 13741 4491 se
rect 13741 4471 13795 4491
tri 13795 4471 13815 4491 nw
tri 17284 4471 17304 4491 ne
rect 17304 4471 18051 4491
tri 18051 4471 18220 4640 nw
tri 13741 4417 13795 4471 nw
tri 13615 4365 13667 4417 se
rect 13615 4140 13667 4365
tri 13667 4343 13741 4417 nw
tri 12245 4088 12261 4104 sw
rect 12193 4076 12261 4088
tri 12261 4076 12273 4088 sw
rect 13615 4076 13667 4088
rect 12193 4070 12273 4076
tri 12273 4070 12279 4076 sw
rect 12193 4018 12199 4070
rect 12251 4018 12263 4070
rect 12315 4018 12321 4070
rect 13615 4018 13667 4024
tri 12002 3917 12054 3969 nw
tri 11871 3860 11928 3917 se
tri 11854 3843 11871 3860 se
rect 11871 3843 11928 3860
tri 11928 3843 12002 3917 nw
tri 11780 3769 11854 3843 se
tri 11854 3769 11928 3843 nw
tri 11775 3764 11780 3769 se
rect 11780 3764 11810 3769
tri 11234 3725 11273 3764 sw
tri 11736 3725 11775 3764 se
rect 11775 3725 11810 3764
tri 11810 3725 11854 3769 nw
rect 11182 3673 11758 3725
tri 11758 3673 11810 3725 nw
rect 11182 3634 11234 3673
tri 11234 3634 11273 3673 nw
<< via2 >>
rect 16123 6547 16179 6603
rect 16218 6547 16274 6603
rect 16123 6467 16179 6523
rect 16218 6467 16274 6523
<< metal3 >>
rect 16118 6603 16279 6608
rect 16118 6547 16123 6603
rect 16179 6547 16218 6603
rect 16274 6547 16279 6603
rect 16118 6523 16279 6547
rect 16118 6467 16123 6523
rect 16179 6467 16218 6523
rect 16274 6467 16279 6523
rect 16118 6462 16279 6467
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1640697850
transform -1 0 11562 0 -1 4614
box -42 24 569 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1640697850
transform 1 0 11380 0 -1 4614
box -46 24 399 1116
use sky130_fd_io__gpiov2_ctl_lsbank  sky130_fd_io__gpiov2_ctl_lsbank_0
timestamp 1640697850
transform -1 0 19429 0 -1 6852
box 883 -1325 16008 3354
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1640697850
transform -1 0 12214 0 -1 4614
box 0 24 534 1116
use sky130_fd_io__com_ctl_hldv2  sky130_fd_io__com_ctl_hldv2_0
timestamp 1640697850
transform -1 0 12986 0 -1 8050
box 417 1201 9109 4552
<< labels >>
flabel metal2 s 6476 6791 6528 6843 3 FreeSans 520 270 0 0 VTRIP_SEL_H_N
port 1 nsew
flabel metal2 s 13475 4854 13527 4906 3 FreeSans 520 90 0 0 DM[0]
port 2 nsew
flabel metal2 s 9346 4854 9398 4906 3 FreeSans 520 90 0 0 DM[2]
port 3 nsew
flabel metal2 s 14776 6791 14828 6843 3 FreeSans 520 270 0 0 DM_H[0]
port 4 nsew
flabel metal2 s 15564 6791 15616 6843 3 FreeSans 520 270 0 0 DM_H[1]
port 5 nsew
flabel metal2 s 8837 3843 8865 3867 3 FreeSans 520 180 0 0 HLD_OVR
port 6 nsew
flabel metal2 s 10622 6791 10674 6843 3 FreeSans 520 270 0 0 DM_H[2]
port 7 nsew
flabel metal2 s 14870 6791 14922 6843 3 FreeSans 520 270 0 0 DM_H_N[0]
port 8 nsew
flabel metal2 s 15470 6791 15522 6843 3 FreeSans 520 270 0 0 DM_H_N[1]
port 9 nsew
flabel metal2 s 10716 6791 10768 6843 3 FreeSans 520 270 0 0 DM_H_N[2]
port 10 nsew
flabel metal2 s 12675 4854 12727 4906 3 FreeSans 520 90 0 0 INP_DIS
port 11 nsew
flabel metal2 s 11316 6791 11368 6843 3 FreeSans 520 270 0 0 INP_DIS_H_N
port 12 nsew
flabel metal2 s 6382 6791 6434 6843 3 FreeSans 520 270 0 0 VTRIP_SEL_H
port 13 nsew
flabel metal2 s 5193 4854 5245 4906 3 FreeSans 520 90 0 0 VTRIP_SEL
port 14 nsew
flabel metal1 s 16748 5178 16791 5308 0 FreeSans 400 0 0 0 VPWR
port 15 nsew
flabel metal1 s 9889 4208 9931 4265 0 FreeSans 400 0 0 0 HLD_H_N
port 16 nsew
flabel metal1 s 5203 4097 5307 4129 3 FreeSans 520 0 0 0 OD_I_H
port 17 nsew
flabel metal1 s 11632 4190 11660 4259 3 FreeSans 520 0 0 0 INP_STARTUP_EN_H
port 18 nsew
flabel metal1 s 3902 6296 3984 6332 3 FreeSans 520 90 0 0 IB_MODE_SEL_H_N
port 19 nsew
flabel metal1 s 3549 6232 3589 6303 3 FreeSans 520 0 0 0 IB_MODE_SEL_H
port 20 nsew
flabel metal1 s 4690 4793 4762 4826 3 FreeSans 520 0 0 0 IB_MODE_SEL
port 21 nsew
flabel metal1 s 16703 3997 16780 4029 3 FreeSans 520 180 0 0 DM[1]
port 22 nsew
flabel metal1 s 11191 4138 11228 4206 3 FreeSans 520 0 0 0 ENABLE_INP_H
port 23 nsew
flabel metal1 s 16747 4948 16790 5150 3 FreeSans 520 180 0 0 VCC_IO
port 24 nsew
flabel metal1 s 11602 3552 11645 3754 3 FreeSans 520 180 0 0 VCC_IO
port 24 nsew
flabel metal1 s 7222 4096 7344 4129 3 FreeSans 520 180 0 0 HLD_I_H_N
port 25 nsew
flabel metal1 s 10066 4205 10092 4268 3 FreeSans 520 180 0 0 ENABLE_H
port 26 nsew
flabel metal1 s 17224 5946 17267 6145 3 FreeSans 520 180 0 0 VGND
port 27 nsew
flabel metal1 s 4734 4217 4764 4275 3 FreeSans 520 180 0 0 HLD_I_OVR_H
port 28 nsew
flabel metal1 s 16747 5179 16790 5302 3 FreeSans 520 180 0 0 VPWR
port 15 nsew
flabel metal1 s 17224 6642 17267 6843 3 FreeSans 520 180 0 0 VPWR
port 15 nsew
flabel metal1 s 16768 5240 16768 5240 3 FreeSans 520 180 0 0 VPWR
port 15 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 8072420
string GDS_START 8052884
<< end >>
