magic
tech sky130A
magscale 1 2
timestamp 1640697977
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 1 157 187 203
rect 1250 157 1436 203
rect 1 21 1436 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 178 47 208 131
rect 268 47 298 131
rect 352 47 382 131
rect 436 47 466 131
rect 520 47 550 131
rect 708 47 738 131
rect 792 47 822 131
rect 876 47 906 131
rect 965 47 995 131
rect 1061 47 1091 131
rect 1133 47 1163 131
rect 1229 47 1259 131
rect 1328 47 1358 177
<< scpmoshvt >>
rect 79 297 109 497
rect 178 413 208 497
rect 268 413 298 497
rect 352 413 382 497
rect 436 413 466 497
rect 520 413 550 497
rect 708 413 738 497
rect 792 413 822 497
rect 876 413 906 497
rect 965 413 995 497
rect 1061 413 1091 497
rect 1133 413 1163 497
rect 1229 413 1259 497
rect 1328 297 1358 497
<< ndiff >>
rect 27 129 79 177
rect 27 95 35 129
rect 69 95 79 129
rect 27 47 79 95
rect 109 131 161 177
rect 1276 131 1328 177
rect 109 93 178 131
rect 109 59 119 93
rect 153 59 178 93
rect 109 47 178 59
rect 208 47 268 131
rect 298 106 352 131
rect 298 72 308 106
rect 342 72 352 106
rect 298 47 352 72
rect 382 106 436 131
rect 382 72 392 106
rect 426 72 436 106
rect 382 47 436 72
rect 466 89 520 131
rect 466 55 476 89
rect 510 55 520 89
rect 466 47 520 55
rect 550 106 602 131
rect 550 72 560 106
rect 594 72 602 106
rect 550 47 602 72
rect 656 98 708 131
rect 656 64 664 98
rect 698 64 708 98
rect 656 47 708 64
rect 738 106 792 131
rect 738 72 748 106
rect 782 72 792 106
rect 738 47 792 72
rect 822 89 876 131
rect 822 55 832 89
rect 866 55 876 89
rect 822 47 876 55
rect 906 106 965 131
rect 906 72 916 106
rect 950 72 965 106
rect 906 47 965 72
rect 995 101 1061 131
rect 995 67 1017 101
rect 1051 67 1061 101
rect 995 47 1061 67
rect 1091 47 1133 131
rect 1163 47 1229 131
rect 1259 89 1328 131
rect 1259 55 1269 89
rect 1303 55 1328 89
rect 1259 47 1328 55
rect 1358 129 1410 177
rect 1358 95 1368 129
rect 1402 95 1410 129
rect 1358 47 1410 95
<< pdiff >>
rect 27 466 79 497
rect 27 432 35 466
rect 69 432 79 466
rect 27 372 79 432
rect 27 338 35 372
rect 69 338 79 372
rect 27 297 79 338
rect 109 481 178 497
rect 109 447 119 481
rect 153 447 178 481
rect 109 413 178 447
rect 208 413 268 497
rect 298 472 352 497
rect 298 438 308 472
rect 342 438 352 472
rect 298 413 352 438
rect 382 472 436 497
rect 382 438 392 472
rect 426 438 436 472
rect 382 413 436 438
rect 466 489 520 497
rect 466 455 476 489
rect 510 455 520 489
rect 466 413 520 455
rect 550 472 602 497
rect 550 438 560 472
rect 594 438 602 472
rect 550 413 602 438
rect 656 485 708 497
rect 656 451 664 485
rect 698 451 708 485
rect 656 413 708 451
rect 738 472 792 497
rect 738 438 748 472
rect 782 438 792 472
rect 738 413 792 438
rect 822 489 876 497
rect 822 455 832 489
rect 866 455 876 489
rect 822 413 876 455
rect 906 472 965 497
rect 906 438 916 472
rect 950 438 965 472
rect 906 413 965 438
rect 995 477 1061 497
rect 995 443 1017 477
rect 1051 443 1061 477
rect 995 413 1061 443
rect 1091 413 1133 497
rect 1163 413 1229 497
rect 1259 489 1328 497
rect 1259 455 1284 489
rect 1318 455 1328 489
rect 1259 413 1328 455
rect 109 297 161 413
rect 1276 297 1328 413
rect 1358 459 1410 497
rect 1358 425 1368 459
rect 1402 425 1410 459
rect 1358 369 1410 425
rect 1358 335 1368 369
rect 1402 335 1410 369
rect 1358 297 1410 335
<< ndiffc >>
rect 35 95 69 129
rect 119 59 153 93
rect 308 72 342 106
rect 392 72 426 106
rect 476 55 510 89
rect 560 72 594 106
rect 664 64 698 98
rect 748 72 782 106
rect 832 55 866 89
rect 916 72 950 106
rect 1017 67 1051 101
rect 1269 55 1303 89
rect 1368 95 1402 129
<< pdiffc >>
rect 35 432 69 466
rect 35 338 69 372
rect 119 447 153 481
rect 308 438 342 472
rect 392 438 426 472
rect 476 455 510 489
rect 560 438 594 472
rect 664 451 698 485
rect 748 438 782 472
rect 832 455 866 489
rect 916 438 950 472
rect 1017 443 1051 477
rect 1284 455 1318 489
rect 1368 425 1402 459
rect 1368 335 1402 369
<< poly >>
rect 79 497 109 523
rect 178 497 208 523
rect 268 497 298 523
rect 352 497 382 523
rect 436 497 466 523
rect 520 497 550 523
rect 708 497 738 523
rect 792 497 822 523
rect 876 497 906 523
rect 965 497 995 523
rect 1061 497 1091 523
rect 1133 497 1163 523
rect 1229 497 1259 523
rect 1328 497 1358 523
rect 79 265 109 297
rect 178 265 208 413
rect 268 376 298 413
rect 250 360 304 376
rect 250 326 260 360
rect 294 326 304 360
rect 250 310 304 326
rect 76 249 130 265
rect 76 215 86 249
rect 120 215 130 249
rect 76 199 130 215
rect 172 249 226 265
rect 172 215 182 249
rect 216 215 226 249
rect 172 199 226 215
rect 79 177 109 199
rect 178 131 208 199
rect 268 131 298 310
rect 352 271 382 413
rect 436 272 466 413
rect 520 398 550 413
rect 708 398 738 413
rect 520 368 738 398
rect 663 337 727 368
rect 792 353 822 413
rect 663 303 673 337
rect 707 303 727 337
rect 663 287 727 303
rect 780 337 834 353
rect 780 303 790 337
rect 824 303 834 337
rect 780 287 834 303
rect 340 255 394 271
rect 340 221 350 255
rect 384 221 394 255
rect 340 205 394 221
rect 436 256 490 272
rect 436 222 446 256
rect 480 222 490 256
rect 436 206 490 222
rect 352 131 382 205
rect 436 131 466 206
rect 697 191 727 287
rect 697 176 738 191
rect 793 176 823 287
rect 876 241 906 413
rect 965 241 995 413
rect 1061 369 1091 413
rect 1037 353 1091 369
rect 1037 319 1047 353
rect 1081 319 1091 353
rect 1037 303 1091 319
rect 520 146 738 176
rect 520 131 550 146
rect 708 131 738 146
rect 792 146 823 176
rect 865 225 919 241
rect 865 191 875 225
rect 909 191 919 225
rect 865 175 919 191
rect 965 225 1019 241
rect 965 191 975 225
rect 1009 191 1019 225
rect 965 175 1019 191
rect 792 131 822 146
rect 876 131 906 175
rect 965 131 995 175
rect 1061 131 1091 303
rect 1133 369 1163 413
rect 1133 353 1187 369
rect 1133 319 1143 353
rect 1177 319 1187 353
rect 1133 303 1187 319
rect 1133 131 1163 303
rect 1229 257 1259 413
rect 1328 265 1358 297
rect 1205 241 1259 257
rect 1205 207 1215 241
rect 1249 207 1259 241
rect 1205 191 1259 207
rect 1304 249 1358 265
rect 1304 215 1314 249
rect 1348 215 1358 249
rect 1304 199 1358 215
rect 1229 131 1259 191
rect 1328 177 1358 199
rect 79 21 109 47
rect 178 21 208 47
rect 268 21 298 47
rect 352 21 382 47
rect 436 21 466 47
rect 520 21 550 47
rect 708 21 738 47
rect 792 21 822 47
rect 876 21 906 47
rect 965 21 995 47
rect 1061 21 1091 47
rect 1133 21 1163 47
rect 1229 21 1259 47
rect 1328 21 1358 47
<< polycont >>
rect 260 326 294 360
rect 86 215 120 249
rect 182 215 216 249
rect 673 303 707 337
rect 790 303 824 337
rect 350 221 384 255
rect 446 222 480 256
rect 1047 319 1081 353
rect 875 191 909 225
rect 975 191 1009 225
rect 1143 319 1177 353
rect 1215 207 1249 241
rect 1314 215 1348 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 17 466 69 493
rect 17 432 35 466
rect 17 372 69 432
rect 103 481 153 527
rect 103 447 119 481
rect 103 430 153 447
rect 187 472 342 493
rect 187 438 308 472
rect 187 413 342 438
rect 392 472 426 493
rect 460 489 526 527
rect 460 455 476 489
rect 510 455 526 489
rect 560 472 607 493
rect 392 421 426 438
rect 594 438 607 472
rect 648 485 714 527
rect 648 451 664 485
rect 698 451 714 485
rect 748 472 782 493
rect 560 421 607 438
rect 187 389 221 413
rect 17 338 35 372
rect 17 297 69 338
rect 103 325 221 389
rect 392 387 607 421
rect 816 489 882 527
rect 816 455 832 489
rect 866 455 882 489
rect 916 472 950 493
rect 748 421 782 438
rect 916 421 950 438
rect 1017 477 1234 493
rect 1051 443 1234 477
rect 1268 489 1334 527
rect 1268 455 1284 489
rect 1318 455 1334 489
rect 1368 459 1448 493
rect 1017 425 1234 443
rect 748 387 950 421
rect 1200 421 1234 425
rect 1402 425 1448 459
rect 260 360 340 376
rect 294 326 340 360
rect 1031 353 1081 391
rect 1200 387 1333 421
rect 17 166 52 297
rect 103 265 137 325
rect 260 323 340 326
rect 260 289 306 323
rect 374 319 592 353
rect 86 249 137 265
rect 120 215 137 249
rect 86 199 137 215
rect 182 255 216 265
rect 374 255 408 319
rect 182 249 214 255
rect 334 221 350 255
rect 384 221 408 255
rect 446 256 524 272
rect 480 255 524 256
rect 480 222 490 255
rect 446 221 490 222
rect 216 215 248 221
rect 182 199 248 215
rect 446 206 524 221
rect 558 250 592 319
rect 640 337 712 353
rect 1031 337 1047 353
rect 640 303 673 337
rect 707 323 712 337
rect 640 289 678 303
rect 640 287 712 289
rect 757 303 790 337
rect 824 319 1047 337
rect 824 303 1081 319
rect 1127 323 1143 353
rect 757 250 791 303
rect 1127 289 1138 323
rect 1177 319 1211 353
rect 1172 289 1211 319
rect 1299 265 1333 387
rect 1368 369 1448 425
rect 1402 335 1448 369
rect 1368 297 1448 335
rect 17 129 69 166
rect 17 95 35 129
rect 103 161 137 199
rect 558 193 791 250
rect 850 221 862 255
rect 896 225 925 255
rect 1177 241 1230 255
rect 850 191 875 221
rect 909 191 925 225
rect 959 191 975 225
rect 1009 191 1092 225
rect 1177 207 1215 241
rect 1264 221 1265 255
rect 1249 207 1265 221
rect 1299 249 1348 265
rect 1299 215 1314 249
rect 993 187 1092 191
rect 294 161 306 187
rect 103 153 306 161
rect 340 153 342 187
rect 103 127 342 153
rect 17 51 69 95
rect 222 106 342 127
rect 103 59 119 93
rect 153 59 169 93
rect 103 17 169 59
rect 222 72 308 106
rect 222 51 342 72
rect 392 123 594 157
rect 392 106 426 123
rect 560 106 594 123
rect 392 51 426 72
rect 460 55 476 89
rect 510 55 526 89
rect 460 17 526 55
rect 748 123 950 157
rect 993 153 1046 187
rect 1080 153 1092 187
rect 1299 199 1348 215
rect 1299 157 1333 199
rect 1382 162 1448 297
rect 748 106 782 123
rect 560 51 594 72
rect 648 64 664 98
rect 698 64 714 98
rect 648 17 714 64
rect 916 106 950 123
rect 1185 123 1333 157
rect 1368 129 1448 162
rect 748 51 782 72
rect 816 55 832 89
rect 866 55 882 89
rect 816 17 882 55
rect 916 51 950 72
rect 1017 101 1051 119
rect 1185 101 1219 123
rect 1051 67 1219 101
rect 1402 95 1448 129
rect 1017 51 1219 67
rect 1253 55 1269 89
rect 1303 55 1319 89
rect 1253 17 1319 55
rect 1368 51 1448 95
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 306 289 340 323
rect 214 249 248 255
rect 214 221 216 249
rect 216 221 248 249
rect 490 221 524 255
rect 678 303 707 323
rect 707 303 712 323
rect 678 289 712 303
rect 1138 319 1143 323
rect 1143 319 1172 323
rect 1138 289 1172 319
rect 862 225 896 255
rect 1230 241 1264 255
rect 862 221 875 225
rect 875 221 896 225
rect 1230 221 1249 241
rect 1249 221 1264 241
rect 306 153 340 187
rect 1046 153 1080 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 294 323 352 329
rect 294 289 306 323
rect 340 320 352 323
rect 666 323 724 329
rect 666 320 678 323
rect 340 292 678 320
rect 340 289 352 292
rect 294 283 352 289
rect 666 289 678 292
rect 712 320 724 323
rect 1126 323 1184 329
rect 1126 320 1138 323
rect 712 292 1138 320
rect 712 289 724 292
rect 666 283 724 289
rect 1126 289 1138 292
rect 1172 289 1184 323
rect 1126 283 1184 289
rect 202 255 260 261
rect 202 221 214 255
rect 248 252 260 255
rect 478 255 536 261
rect 478 252 490 255
rect 248 224 490 252
rect 248 221 260 224
rect 202 215 260 221
rect 478 221 490 224
rect 524 252 536 255
rect 850 255 908 261
rect 850 252 862 255
rect 524 224 862 252
rect 524 221 536 224
rect 478 215 536 221
rect 850 221 862 224
rect 896 252 908 255
rect 1218 255 1276 261
rect 1218 252 1230 255
rect 896 224 1230 252
rect 896 221 908 224
rect 850 215 908 221
rect 1218 221 1230 224
rect 1264 221 1276 255
rect 1218 215 1276 221
rect 294 187 352 193
rect 294 153 306 187
rect 340 184 352 187
rect 1034 187 1092 193
rect 1034 184 1046 187
rect 340 156 1046 184
rect 340 153 352 156
rect 294 147 352 153
rect 1034 153 1046 156
rect 1080 153 1092 187
rect 1034 147 1092 153
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel locali s 30 425 64 459 0 FreeSans 200 0 0 0 COUT
port 8 nsew signal output
flabel locali s 30 357 64 391 0 FreeSans 200 0 0 0 COUT
port 8 nsew signal output
flabel locali s 30 85 64 119 0 FreeSans 200 0 0 0 COUT
port 8 nsew signal output
flabel locali s 1046 357 1080 391 0 FreeSans 200 0 0 0 CIN
port 3 nsew signal input
flabel locali s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel locali s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 1414 85 1448 119 0 FreeSans 200 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1414 153 1448 187 0 FreeSans 200 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1414 221 1448 255 0 FreeSans 200 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1414 289 1448 323 0 FreeSans 200 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1414 357 1448 391 0 FreeSans 200 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1414 425 1448 459 0 FreeSans 200 0 0 0 SUM
port 9 nsew signal output
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 306 289 340 323 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 fa_1
rlabel locali s 446 206 524 272 1 A
port 1 nsew signal input
rlabel locali s 850 191 925 255 1 A
port 1 nsew signal input
rlabel locali s 1177 207 1265 255 1 A
port 1 nsew signal input
rlabel metal1 s 1218 252 1276 261 1 A
port 1 nsew signal input
rlabel metal1 s 1218 215 1276 224 1 A
port 1 nsew signal input
rlabel metal1 s 850 252 908 261 1 A
port 1 nsew signal input
rlabel metal1 s 850 215 908 224 1 A
port 1 nsew signal input
rlabel metal1 s 478 252 536 261 1 A
port 1 nsew signal input
rlabel metal1 s 478 215 536 224 1 A
port 1 nsew signal input
rlabel metal1 s 202 252 260 261 1 A
port 1 nsew signal input
rlabel metal1 s 202 224 1276 252 1 A
port 1 nsew signal input
rlabel metal1 s 202 215 260 224 1 A
port 1 nsew signal input
rlabel locali s 640 287 712 353 1 B
port 2 nsew signal input
rlabel locali s 1127 289 1211 353 1 B
port 2 nsew signal input
rlabel metal1 s 1126 320 1184 329 1 B
port 2 nsew signal input
rlabel metal1 s 1126 283 1184 292 1 B
port 2 nsew signal input
rlabel metal1 s 666 320 724 329 1 B
port 2 nsew signal input
rlabel metal1 s 666 283 724 292 1 B
port 2 nsew signal input
rlabel metal1 s 294 320 352 329 1 B
port 2 nsew signal input
rlabel metal1 s 294 292 1184 320 1 B
port 2 nsew signal input
rlabel metal1 s 294 283 352 292 1 B
port 2 nsew signal input
rlabel metal1 s 0 -48 1472 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1472 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 2064582
string GDS_START 2051632
string path 0.000 0.000 36.800 0.000 
<< end >>
