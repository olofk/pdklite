magic
tech sky130A
magscale 1 2
timestamp 1640697850
<< nwell >>
rect 56 1378 843 1486
rect 56 1320 1033 1378
rect 23 884 1033 1320
<< pwell >>
rect 183 522 973 774
rect 1194 732 2240 1314
rect 1417 340 2268 389
rect 657 137 2268 340
rect 657 46 1987 137
rect 146 37 1987 46
rect 146 -40 1366 37
<< mvnmos >>
rect 736 114 836 314
rect 892 114 992 314
rect 1048 114 1148 314
rect 1204 114 1304 314
rect 1496 63 1596 363
rect 1652 63 1752 363
rect 1808 63 1908 363
rect 2089 163 2189 363
<< mvpmos >>
rect 206 1159 356 1259
rect 544 1159 694 1259
rect 817 1159 967 1259
rect 206 1003 356 1103
rect 544 1003 694 1103
rect 817 1003 967 1103
<< mvnnmos >>
rect 1273 1088 1453 1288
rect 1509 1088 1689 1288
rect 1745 1088 1925 1288
rect 1981 1088 2161 1288
rect 1273 758 1453 958
rect 1509 758 1689 958
rect 1745 758 1925 958
rect 1981 758 2161 958
<< nmoslvt >>
rect 262 548 292 748
rect 348 548 378 748
rect 434 548 464 748
rect 520 548 550 748
rect 606 548 636 748
rect 692 548 722 748
rect 778 548 808 748
rect 864 548 894 748
<< ndiff >>
rect 209 736 262 748
rect 209 702 217 736
rect 251 702 262 736
rect 209 668 262 702
rect 209 634 217 668
rect 251 634 262 668
rect 209 600 262 634
rect 209 566 217 600
rect 251 566 262 600
rect 209 548 262 566
rect 292 736 348 748
rect 292 702 303 736
rect 337 702 348 736
rect 292 668 348 702
rect 292 634 303 668
rect 337 634 348 668
rect 292 600 348 634
rect 292 566 303 600
rect 337 566 348 600
rect 292 548 348 566
rect 378 736 434 748
rect 378 702 389 736
rect 423 702 434 736
rect 378 668 434 702
rect 378 634 389 668
rect 423 634 434 668
rect 378 600 434 634
rect 378 566 389 600
rect 423 566 434 600
rect 378 548 434 566
rect 464 736 520 748
rect 464 702 475 736
rect 509 702 520 736
rect 464 668 520 702
rect 464 634 475 668
rect 509 634 520 668
rect 464 600 520 634
rect 464 566 475 600
rect 509 566 520 600
rect 464 548 520 566
rect 550 736 606 748
rect 550 702 561 736
rect 595 702 606 736
rect 550 668 606 702
rect 550 634 561 668
rect 595 634 606 668
rect 550 600 606 634
rect 550 566 561 600
rect 595 566 606 600
rect 550 548 606 566
rect 636 736 692 748
rect 636 702 647 736
rect 681 702 692 736
rect 636 668 692 702
rect 636 634 647 668
rect 681 634 692 668
rect 636 600 692 634
rect 636 566 647 600
rect 681 566 692 600
rect 636 548 692 566
rect 722 736 778 748
rect 722 702 733 736
rect 767 702 778 736
rect 722 668 778 702
rect 722 634 733 668
rect 767 634 778 668
rect 722 600 778 634
rect 722 566 733 600
rect 767 566 778 600
rect 722 548 778 566
rect 808 736 864 748
rect 808 702 819 736
rect 853 702 864 736
rect 808 668 864 702
rect 808 634 819 668
rect 853 634 864 668
rect 808 600 864 634
rect 808 566 819 600
rect 853 566 864 600
rect 808 548 864 566
rect 894 736 947 748
rect 894 702 905 736
rect 939 702 947 736
rect 894 668 947 702
rect 894 634 905 668
rect 939 634 947 668
rect 894 600 947 634
rect 894 566 905 600
rect 939 566 947 600
rect 894 548 947 566
<< mvndiff >>
rect 1220 1276 1273 1288
rect 1220 1242 1228 1276
rect 1262 1242 1273 1276
rect 1220 1208 1273 1242
rect 1220 1174 1228 1208
rect 1262 1174 1273 1208
rect 1220 1140 1273 1174
rect 1220 1106 1228 1140
rect 1262 1106 1273 1140
rect 1220 1088 1273 1106
rect 1453 1276 1509 1288
rect 1453 1242 1464 1276
rect 1498 1242 1509 1276
rect 1453 1208 1509 1242
rect 1453 1174 1464 1208
rect 1498 1174 1509 1208
rect 1453 1140 1509 1174
rect 1453 1106 1464 1140
rect 1498 1106 1509 1140
rect 1453 1088 1509 1106
rect 1689 1276 1745 1288
rect 1689 1242 1700 1276
rect 1734 1242 1745 1276
rect 1689 1208 1745 1242
rect 1689 1174 1700 1208
rect 1734 1174 1745 1208
rect 1689 1140 1745 1174
rect 1689 1106 1700 1140
rect 1734 1106 1745 1140
rect 1689 1088 1745 1106
rect 1925 1276 1981 1288
rect 1925 1242 1936 1276
rect 1970 1242 1981 1276
rect 1925 1208 1981 1242
rect 1925 1174 1936 1208
rect 1970 1174 1981 1208
rect 1925 1140 1981 1174
rect 1925 1106 1936 1140
rect 1970 1106 1981 1140
rect 1925 1088 1981 1106
rect 2161 1276 2214 1288
rect 2161 1242 2172 1276
rect 2206 1242 2214 1276
rect 2161 1208 2214 1242
rect 2161 1174 2172 1208
rect 2206 1174 2214 1208
rect 2161 1140 2214 1174
rect 2161 1106 2172 1140
rect 2206 1106 2214 1140
rect 2161 1088 2214 1106
rect 1220 940 1273 958
rect 1220 906 1228 940
rect 1262 906 1273 940
rect 1220 872 1273 906
rect 1220 838 1228 872
rect 1262 838 1273 872
rect 1220 804 1273 838
rect 1220 770 1228 804
rect 1262 770 1273 804
rect 1220 758 1273 770
rect 1453 940 1509 958
rect 1453 906 1464 940
rect 1498 906 1509 940
rect 1453 872 1509 906
rect 1453 838 1464 872
rect 1498 838 1509 872
rect 1453 804 1509 838
rect 1453 770 1464 804
rect 1498 770 1509 804
rect 1453 758 1509 770
rect 1689 940 1745 958
rect 1689 906 1700 940
rect 1734 906 1745 940
rect 1689 872 1745 906
rect 1689 838 1700 872
rect 1734 838 1745 872
rect 1689 804 1745 838
rect 1689 770 1700 804
rect 1734 770 1745 804
rect 1689 758 1745 770
rect 1925 940 1981 958
rect 1925 906 1936 940
rect 1970 906 1981 940
rect 1925 872 1981 906
rect 1925 838 1936 872
rect 1970 838 1981 872
rect 1925 804 1981 838
rect 1925 770 1936 804
rect 1970 770 1981 804
rect 1925 758 1981 770
rect 2161 940 2214 958
rect 2161 906 2172 940
rect 2206 906 2214 940
rect 2161 872 2214 906
rect 2161 838 2172 872
rect 2206 838 2214 872
rect 2161 804 2214 838
rect 2161 770 2172 804
rect 2206 770 2214 804
rect 2161 758 2214 770
rect 1443 351 1496 363
rect 1443 317 1451 351
rect 1485 317 1496 351
rect 683 296 736 314
rect 683 262 691 296
rect 725 262 736 296
rect 683 228 736 262
rect 683 194 691 228
rect 725 194 736 228
rect 683 160 736 194
rect 683 126 691 160
rect 725 126 736 160
rect 683 114 736 126
rect 836 296 892 314
rect 836 262 847 296
rect 881 262 892 296
rect 836 228 892 262
rect 836 194 847 228
rect 881 194 892 228
rect 836 160 892 194
rect 836 126 847 160
rect 881 126 892 160
rect 836 114 892 126
rect 992 296 1048 314
rect 992 262 1003 296
rect 1037 262 1048 296
rect 992 228 1048 262
rect 992 194 1003 228
rect 1037 194 1048 228
rect 992 160 1048 194
rect 992 126 1003 160
rect 1037 126 1048 160
rect 992 114 1048 126
rect 1148 296 1204 314
rect 1148 262 1159 296
rect 1193 262 1204 296
rect 1148 228 1204 262
rect 1148 194 1159 228
rect 1193 194 1204 228
rect 1148 160 1204 194
rect 1148 126 1159 160
rect 1193 126 1204 160
rect 1148 114 1204 126
rect 1304 296 1357 314
rect 1304 262 1315 296
rect 1349 262 1357 296
rect 1304 228 1357 262
rect 1304 194 1315 228
rect 1349 194 1357 228
rect 1304 160 1357 194
rect 1304 126 1315 160
rect 1349 126 1357 160
rect 1304 114 1357 126
rect 1443 283 1496 317
rect 1443 249 1451 283
rect 1485 249 1496 283
rect 1443 215 1496 249
rect 1443 181 1451 215
rect 1485 181 1496 215
rect 1443 147 1496 181
rect 1443 113 1451 147
rect 1485 113 1496 147
rect 1443 63 1496 113
rect 1596 351 1652 363
rect 1596 317 1607 351
rect 1641 317 1652 351
rect 1596 283 1652 317
rect 1596 249 1607 283
rect 1641 249 1652 283
rect 1596 215 1652 249
rect 1596 181 1607 215
rect 1641 181 1652 215
rect 1596 147 1652 181
rect 1596 113 1607 147
rect 1641 113 1652 147
rect 1596 63 1652 113
rect 1752 351 1808 363
rect 1752 317 1763 351
rect 1797 317 1808 351
rect 1752 283 1808 317
rect 1752 249 1763 283
rect 1797 249 1808 283
rect 1752 215 1808 249
rect 1752 181 1763 215
rect 1797 181 1808 215
rect 1752 147 1808 181
rect 1752 113 1763 147
rect 1797 113 1808 147
rect 1752 63 1808 113
rect 1908 351 1961 363
rect 1908 317 1919 351
rect 1953 317 1961 351
rect 1908 283 1961 317
rect 1908 249 1919 283
rect 1953 249 1961 283
rect 1908 215 1961 249
rect 1908 181 1919 215
rect 1953 181 1961 215
rect 1908 147 1961 181
rect 2036 351 2089 363
rect 2036 317 2044 351
rect 2078 317 2089 351
rect 2036 283 2089 317
rect 2036 249 2044 283
rect 2078 249 2089 283
rect 2036 215 2089 249
rect 2036 181 2044 215
rect 2078 181 2089 215
rect 2036 163 2089 181
rect 2189 351 2242 363
rect 2189 317 2200 351
rect 2234 317 2242 351
rect 2189 283 2242 317
rect 2189 249 2200 283
rect 2234 249 2242 283
rect 2189 215 2242 249
rect 2189 181 2200 215
rect 2234 181 2242 215
rect 2189 163 2242 181
rect 1908 113 1919 147
rect 1953 113 1961 147
rect 1908 63 1961 113
<< mvpdiff >>
rect 206 1304 356 1312
rect 206 1270 218 1304
rect 252 1270 286 1304
rect 320 1270 356 1304
rect 206 1259 356 1270
rect 544 1304 694 1312
rect 544 1270 556 1304
rect 590 1270 624 1304
rect 658 1270 694 1304
rect 544 1259 694 1270
rect 817 1304 967 1312
rect 817 1270 829 1304
rect 863 1270 897 1304
rect 931 1270 967 1304
rect 817 1259 967 1270
rect 206 1148 356 1159
rect 206 1114 218 1148
rect 252 1114 286 1148
rect 320 1114 356 1148
rect 206 1103 356 1114
rect 544 1148 694 1159
rect 544 1114 556 1148
rect 590 1114 624 1148
rect 658 1114 694 1148
rect 544 1103 694 1114
rect 817 1148 967 1159
rect 817 1114 829 1148
rect 863 1114 897 1148
rect 931 1114 967 1148
rect 817 1103 967 1114
rect 206 992 356 1003
rect 206 958 218 992
rect 252 958 286 992
rect 320 958 356 992
rect 206 950 356 958
rect 544 992 694 1003
rect 544 958 556 992
rect 590 958 624 992
rect 658 958 694 992
rect 544 950 694 958
rect 817 992 967 1003
rect 817 958 829 992
rect 863 958 897 992
rect 931 958 967 992
rect 817 950 967 958
<< ndiffc >>
rect 217 702 251 736
rect 217 634 251 668
rect 217 566 251 600
rect 303 702 337 736
rect 303 634 337 668
rect 303 566 337 600
rect 389 702 423 736
rect 389 634 423 668
rect 389 566 423 600
rect 475 702 509 736
rect 475 634 509 668
rect 475 566 509 600
rect 561 702 595 736
rect 561 634 595 668
rect 561 566 595 600
rect 647 702 681 736
rect 647 634 681 668
rect 647 566 681 600
rect 733 702 767 736
rect 733 634 767 668
rect 733 566 767 600
rect 819 702 853 736
rect 819 634 853 668
rect 819 566 853 600
rect 905 702 939 736
rect 905 634 939 668
rect 905 566 939 600
<< mvndiffc >>
rect 1228 1242 1262 1276
rect 1228 1174 1262 1208
rect 1228 1106 1262 1140
rect 1464 1242 1498 1276
rect 1464 1174 1498 1208
rect 1464 1106 1498 1140
rect 1700 1242 1734 1276
rect 1700 1174 1734 1208
rect 1700 1106 1734 1140
rect 1936 1242 1970 1276
rect 1936 1174 1970 1208
rect 1936 1106 1970 1140
rect 2172 1242 2206 1276
rect 2172 1174 2206 1208
rect 2172 1106 2206 1140
rect 1228 906 1262 940
rect 1228 838 1262 872
rect 1228 770 1262 804
rect 1464 906 1498 940
rect 1464 838 1498 872
rect 1464 770 1498 804
rect 1700 906 1734 940
rect 1700 838 1734 872
rect 1700 770 1734 804
rect 1936 906 1970 940
rect 1936 838 1970 872
rect 1936 770 1970 804
rect 2172 906 2206 940
rect 2172 838 2206 872
rect 2172 770 2206 804
rect 1451 317 1485 351
rect 691 262 725 296
rect 691 194 725 228
rect 691 126 725 160
rect 847 262 881 296
rect 847 194 881 228
rect 847 126 881 160
rect 1003 262 1037 296
rect 1003 194 1037 228
rect 1003 126 1037 160
rect 1159 262 1193 296
rect 1159 194 1193 228
rect 1159 126 1193 160
rect 1315 262 1349 296
rect 1315 194 1349 228
rect 1315 126 1349 160
rect 1451 249 1485 283
rect 1451 181 1485 215
rect 1451 113 1485 147
rect 1607 317 1641 351
rect 1607 249 1641 283
rect 1607 181 1641 215
rect 1607 113 1641 147
rect 1763 317 1797 351
rect 1763 249 1797 283
rect 1763 181 1797 215
rect 1763 113 1797 147
rect 1919 317 1953 351
rect 1919 249 1953 283
rect 1919 181 1953 215
rect 2044 317 2078 351
rect 2044 249 2078 283
rect 2044 181 2078 215
rect 2200 317 2234 351
rect 2200 249 2234 283
rect 2200 181 2234 215
rect 1919 113 1953 147
<< mvpdiffc >>
rect 218 1270 252 1304
rect 286 1270 320 1304
rect 556 1270 590 1304
rect 624 1270 658 1304
rect 829 1270 863 1304
rect 897 1270 931 1304
rect 218 1114 252 1148
rect 286 1114 320 1148
rect 556 1114 590 1148
rect 624 1114 658 1148
rect 829 1114 863 1148
rect 897 1114 931 1148
rect 218 958 252 992
rect 286 958 320 992
rect 556 958 590 992
rect 624 958 658 992
rect 829 958 863 992
rect 897 958 931 992
<< psubdiff >>
rect 172 -14 196 0
rect 230 -14 269 0
rect 303 -14 342 0
rect 376 -14 415 0
rect 449 -14 488 0
rect 522 -14 561 0
rect 595 -14 634 0
rect 668 -14 706 0
rect 740 -14 778 0
rect 812 -14 850 0
rect 884 -14 922 0
rect 956 -14 994 0
rect 1028 -14 1066 0
rect 1100 -14 1138 0
rect 1172 -14 1210 0
rect 1244 -14 1282 0
rect 1316 -14 1340 0
<< mvpsubdiff >>
rect 172 0 196 20
rect 230 0 269 20
rect 303 0 342 20
rect 376 0 415 20
rect 449 0 488 20
rect 522 0 561 20
rect 595 0 634 20
rect 668 0 706 20
rect 740 0 778 20
rect 812 0 850 20
rect 884 0 922 20
rect 956 0 994 20
rect 1028 0 1066 20
rect 1100 0 1138 20
rect 1172 0 1210 20
rect 1244 0 1282 20
rect 1316 0 1340 20
<< mvnsubdiff >>
rect 122 1386 146 1420
rect 180 1386 218 1420
rect 252 1386 290 1420
rect 324 1386 362 1420
rect 396 1386 434 1420
rect 468 1386 506 1420
rect 540 1386 577 1420
rect 611 1386 648 1420
rect 682 1386 719 1420
rect 753 1386 777 1420
<< psubdiffcont >>
rect 196 -14 230 0
rect 269 -14 303 0
rect 342 -14 376 0
rect 415 -14 449 0
rect 488 -14 522 0
rect 561 -14 595 0
rect 634 -14 668 0
rect 706 -14 740 0
rect 778 -14 812 0
rect 850 -14 884 0
rect 922 -14 956 0
rect 994 -14 1028 0
rect 1066 -14 1100 0
rect 1138 -14 1172 0
rect 1210 -14 1244 0
rect 1282 -14 1316 0
<< mvpsubdiffcont >>
rect 196 0 230 20
rect 269 0 303 20
rect 342 0 376 20
rect 415 0 449 20
rect 488 0 522 20
rect 561 0 595 20
rect 634 0 668 20
rect 706 0 740 20
rect 778 0 812 20
rect 850 0 884 20
rect 922 0 956 20
rect 994 0 1028 20
rect 1066 0 1100 20
rect 1138 0 1172 20
rect 1210 0 1244 20
rect 1282 0 1316 20
<< mvnsubdiffcont >>
rect 146 1386 180 1420
rect 218 1386 252 1420
rect 290 1386 324 1420
rect 362 1386 396 1420
rect 434 1386 468 1420
rect 506 1386 540 1420
rect 577 1386 611 1420
rect 648 1386 682 1420
rect 719 1386 753 1420
<< poly >>
rect 1273 1288 1453 1320
rect 1509 1288 1689 1320
rect 1745 1288 1925 1320
rect 1981 1288 2161 1320
rect 999 1270 1065 1286
rect 999 1259 1015 1270
rect 108 1243 206 1259
rect 108 1209 124 1243
rect 158 1209 206 1243
rect 108 1159 206 1209
rect 356 1159 388 1259
rect 446 1243 544 1259
rect 446 1209 462 1243
rect 496 1209 544 1243
rect 446 1159 544 1209
rect 694 1159 726 1259
rect 785 1159 817 1259
rect 967 1236 1015 1259
rect 1049 1236 1065 1270
rect 967 1202 1065 1236
rect 967 1168 1015 1202
rect 1049 1168 1065 1202
rect 967 1159 1065 1168
rect 108 1148 174 1159
rect 108 1114 124 1148
rect 158 1114 174 1148
rect 108 1103 174 1114
rect 446 1148 512 1159
rect 446 1114 462 1148
rect 496 1114 512 1148
rect 446 1103 512 1114
rect 999 1152 1065 1159
rect 999 1103 1065 1109
rect 108 1053 206 1103
rect 108 1019 124 1053
rect 158 1019 206 1053
rect 108 1003 206 1019
rect 356 1003 388 1103
rect 446 1053 544 1103
rect 446 1019 462 1053
rect 496 1019 544 1053
rect 446 1003 544 1019
rect 694 1003 726 1103
rect 785 1003 817 1103
rect 967 1093 1065 1103
rect 967 1059 1015 1093
rect 1049 1059 1065 1093
rect 967 1025 1065 1059
rect 967 1003 1015 1025
rect 999 991 1015 1003
rect 1049 991 1065 1025
rect 999 975 1065 991
rect 1273 1056 1453 1088
rect 1509 1056 1689 1088
rect 1745 1056 1925 1088
rect 1981 1056 2161 1088
rect 1273 1040 2161 1056
rect 1273 1006 1289 1040
rect 1323 1006 1357 1040
rect 1391 1006 1425 1040
rect 1459 1006 1493 1040
rect 1527 1006 1561 1040
rect 1595 1006 1629 1040
rect 1663 1006 1697 1040
rect 1731 1006 1766 1040
rect 1800 1006 1835 1040
rect 1869 1006 1904 1040
rect 1938 1006 1973 1040
rect 2007 1006 2042 1040
rect 2076 1006 2111 1040
rect 2145 1006 2161 1040
rect 1273 990 2161 1006
rect 1273 958 1453 990
rect 1509 958 1689 990
rect 1745 958 1925 990
rect 1981 958 2161 990
rect 262 748 292 780
rect 348 748 378 780
rect 434 748 464 780
rect 520 748 550 780
rect 606 748 636 780
rect 692 748 722 780
rect 778 748 808 780
rect 864 748 894 780
rect 1273 726 1453 758
rect 1509 726 1689 758
rect 1745 726 1925 758
rect 1981 726 2161 758
rect 262 516 292 548
rect 348 516 378 548
rect 434 516 464 548
rect 520 516 550 548
rect 262 500 550 516
rect 262 466 278 500
rect 312 466 352 500
rect 386 466 426 500
rect 460 466 500 500
rect 534 466 550 500
rect 262 450 550 466
rect 606 516 636 548
rect 692 516 722 548
rect 778 516 808 548
rect 864 516 894 548
rect 606 500 894 516
rect 606 466 622 500
rect 656 466 696 500
rect 730 466 770 500
rect 804 466 844 500
rect 878 466 894 500
rect 606 450 894 466
rect 1496 517 1596 533
rect 1496 483 1533 517
rect 1567 483 1596 517
rect 1496 449 1596 483
rect 1496 415 1533 449
rect 1567 415 1596 449
rect 736 390 1304 406
rect 736 356 752 390
rect 786 356 823 390
rect 857 356 894 390
rect 928 356 966 390
rect 1000 356 1038 390
rect 1072 356 1110 390
rect 1144 356 1182 390
rect 1216 356 1254 390
rect 1288 356 1304 390
rect 1496 363 1596 415
rect 1652 517 1752 533
rect 1652 483 1689 517
rect 1723 483 1752 517
rect 1652 449 1752 483
rect 1652 415 1689 449
rect 1723 415 1752 449
rect 1652 363 1752 415
rect 1808 517 1908 533
rect 1808 483 1845 517
rect 1879 483 1908 517
rect 1808 449 1908 483
rect 1808 415 1845 449
rect 1879 415 1908 449
rect 1808 363 1908 415
rect 2089 517 2189 533
rect 2089 483 2125 517
rect 2159 483 2189 517
rect 2089 449 2189 483
rect 2089 415 2125 449
rect 2159 415 2189 449
rect 2089 363 2189 415
rect 736 340 1304 356
rect 736 314 836 340
rect 892 314 992 340
rect 1048 314 1148 340
rect 1204 314 1304 340
rect 736 88 836 114
rect 892 88 992 114
rect 1048 88 1148 114
rect 1204 88 1304 114
rect 2089 131 2189 163
rect 1496 31 1596 63
rect 1652 31 1752 63
rect 1808 31 1908 63
<< polycont >>
rect 124 1209 158 1243
rect 462 1209 496 1243
rect 1015 1236 1049 1270
rect 1015 1168 1049 1202
rect 124 1114 158 1148
rect 462 1114 496 1148
rect 124 1019 158 1053
rect 462 1019 496 1053
rect 1015 1059 1049 1093
rect 1015 991 1049 1025
rect 1289 1006 1323 1040
rect 1357 1006 1391 1040
rect 1425 1006 1459 1040
rect 1493 1006 1527 1040
rect 1561 1006 1595 1040
rect 1629 1006 1663 1040
rect 1697 1006 1731 1040
rect 1766 1006 1800 1040
rect 1835 1006 1869 1040
rect 1904 1006 1938 1040
rect 1973 1006 2007 1040
rect 2042 1006 2076 1040
rect 2111 1006 2145 1040
rect 278 466 312 500
rect 352 466 386 500
rect 426 466 460 500
rect 500 466 534 500
rect 622 466 656 500
rect 696 466 730 500
rect 770 466 804 500
rect 844 466 878 500
rect 1533 483 1567 517
rect 1533 415 1567 449
rect 752 356 786 390
rect 823 356 857 390
rect 894 356 928 390
rect 966 356 1000 390
rect 1038 356 1072 390
rect 1110 356 1144 390
rect 1182 356 1216 390
rect 1254 356 1288 390
rect 1689 483 1723 517
rect 1689 415 1723 449
rect 1845 483 1879 517
rect 1845 415 1879 449
rect 2125 483 2159 517
rect 2125 415 2159 449
<< locali >>
rect 122 1386 134 1420
rect 180 1386 207 1420
rect 252 1386 280 1420
rect 324 1386 354 1420
rect 396 1386 428 1420
rect 468 1386 502 1420
rect 540 1386 576 1420
rect 611 1386 648 1420
rect 684 1386 719 1420
rect 758 1386 777 1420
rect 252 1270 286 1304
rect 540 1270 553 1304
rect 590 1270 624 1304
rect 724 1270 829 1304
rect 863 1270 897 1304
rect 931 1270 947 1304
rect 1015 1270 1049 1286
rect 124 1247 158 1259
rect 152 1243 158 1247
rect 118 1209 124 1213
rect 118 1148 158 1209
rect 462 1243 496 1259
rect 724 1236 775 1270
rect 496 1209 775 1236
rect 462 1182 775 1209
rect 462 1164 496 1182
rect 118 1053 158 1114
rect 202 1154 496 1164
rect 202 1148 462 1154
rect 202 1114 218 1148
rect 252 1114 286 1148
rect 320 1114 462 1148
rect 540 1114 552 1148
rect 590 1114 624 1148
rect 661 1114 674 1148
rect 202 1092 496 1114
rect 118 1049 124 1053
rect 152 1015 158 1019
rect 124 1003 158 1015
rect 462 1079 496 1092
rect 724 1080 775 1182
rect 813 1193 830 1227
rect 864 1193 905 1227
rect 939 1193 947 1227
rect 813 1148 947 1193
rect 1015 1220 1049 1236
rect 1228 1276 1262 1292
rect 1015 1202 1137 1220
rect 1049 1168 1137 1202
rect 1015 1152 1137 1168
rect 813 1114 829 1148
rect 863 1114 897 1148
rect 931 1114 947 1148
rect 1015 1093 1049 1109
rect 724 1063 1015 1080
rect 724 1029 929 1063
rect 963 1029 1004 1063
rect 1038 1029 1049 1059
rect 724 1026 1049 1029
rect 462 1003 496 1019
rect 1015 1025 1049 1026
rect 587 992 653 993
rect 252 958 286 992
rect 540 959 553 992
rect 540 958 556 959
rect 590 958 624 992
rect 658 958 674 959
rect 813 958 829 992
rect 863 958 897 992
rect 931 958 947 992
rect 1015 975 1049 991
rect 813 941 947 958
rect 1083 941 1137 1152
rect 1228 1208 1262 1242
rect 1464 1276 1498 1292
rect 1464 1212 1498 1242
rect 1700 1276 1734 1292
rect 1463 1208 1501 1212
rect 1463 1178 1464 1208
rect 1228 1140 1262 1174
rect 1498 1178 1501 1208
rect 1700 1208 1734 1242
rect 1936 1276 1970 1292
rect 1936 1212 1970 1242
rect 2172 1276 2206 1292
rect 1464 1140 1498 1174
rect 1262 1096 1300 1130
rect 1934 1208 1972 1212
rect 1934 1178 1936 1208
rect 1700 1140 1734 1174
rect 1228 1090 1262 1096
rect 1464 1090 1498 1106
rect 1699 1106 1700 1130
rect 1970 1178 1972 1208
rect 2172 1208 2206 1242
rect 1936 1140 1970 1174
rect 1734 1106 1737 1130
rect 1699 1096 1737 1106
rect 2172 1140 2206 1174
rect 1700 1090 1734 1096
rect 1936 1090 1970 1106
rect 2134 1096 2172 1130
rect 2172 1090 2206 1096
rect 1273 1006 1289 1040
rect 1323 1006 1357 1040
rect 1391 1006 1425 1040
rect 1459 1006 1493 1040
rect 1527 1006 1561 1040
rect 1595 1006 1629 1040
rect 1663 1006 1697 1040
rect 1731 1006 1766 1040
rect 1800 1006 1835 1040
rect 1869 1006 1904 1040
rect 1938 1006 1973 1040
rect 2007 1006 2042 1040
rect 2076 1006 2111 1040
rect 2145 1006 2161 1040
rect 813 907 1007 941
rect 1041 907 1082 941
rect 1116 907 1137 941
rect 813 890 1137 907
rect 217 736 251 752
rect 217 668 251 702
rect 217 600 251 620
rect 303 740 337 778
rect 303 668 337 702
rect 303 600 337 634
rect 303 550 337 566
rect 389 736 423 752
rect 389 668 423 702
rect 389 600 423 620
rect 475 740 509 778
rect 475 668 509 702
rect 475 600 509 634
rect 475 550 509 566
rect 561 736 595 752
rect 561 668 595 702
rect 561 600 595 620
rect 647 740 681 778
rect 647 668 681 702
rect 647 600 681 634
rect 647 550 681 566
rect 733 736 767 752
rect 733 668 767 702
rect 733 600 767 620
rect 819 740 853 778
rect 819 668 853 702
rect 819 600 853 634
rect 819 550 853 566
rect 905 736 939 752
rect 905 668 939 702
rect 905 600 939 620
rect 262 466 278 500
rect 324 466 352 500
rect 386 466 397 500
rect 460 466 500 500
rect 538 466 550 500
rect 606 466 622 500
rect 656 466 696 500
rect 762 466 770 500
rect 804 466 834 500
rect 878 466 894 500
rect 1031 486 1137 890
rect 1228 940 1262 956
rect 1464 943 1498 956
rect 1463 940 1501 943
rect 1463 909 1464 940
rect 1228 872 1262 906
rect 1228 804 1262 838
rect 1224 770 1228 795
rect 1498 909 1501 940
rect 1700 940 1734 956
rect 1936 946 1970 956
rect 1927 940 2018 946
rect 1464 872 1498 906
rect 1464 804 1498 838
rect 1224 761 1262 770
rect 1934 906 1936 940
rect 1970 906 1972 940
rect 2006 906 2018 940
rect 1700 872 1734 906
rect 1700 804 1734 838
rect 1228 754 1262 761
rect 1464 754 1498 770
rect 1699 770 1700 795
rect 1927 872 2018 906
rect 1927 838 1936 872
rect 1970 838 2018 872
rect 1927 804 2018 838
rect 1734 770 1737 795
rect 1699 761 1737 770
rect 1927 770 1936 804
rect 1970 770 2018 804
rect 2172 940 2206 956
rect 2172 872 2206 906
rect 2172 804 2206 838
rect 1700 754 1734 761
rect 1927 754 2018 770
rect 2131 761 2169 795
rect 2203 761 2206 770
rect 2172 754 2206 761
rect 1059 452 1100 486
rect 1134 452 1137 486
rect 1533 525 1567 533
rect 1533 453 1567 483
rect 1533 399 1567 415
rect 1689 525 1723 533
rect 1689 453 1723 483
rect 1689 399 1723 415
rect 1845 525 1879 533
rect 1845 453 1879 483
rect 2154 517 2159 533
rect 2120 483 2125 501
rect 2120 463 2159 483
rect 2154 449 2159 463
rect 1845 399 1879 415
rect 2125 399 2159 415
rect 838 390 882 395
rect 916 390 960 395
rect 994 390 1038 395
rect 1072 390 1116 395
rect 1150 390 1194 395
rect 736 356 752 390
rect 786 361 804 390
rect 857 361 882 390
rect 928 361 960 390
rect 786 356 823 361
rect 857 356 894 361
rect 928 356 966 361
rect 1000 356 1038 390
rect 1072 356 1110 390
rect 1150 361 1182 390
rect 1228 361 1254 390
rect 1144 356 1182 361
rect 1216 356 1254 361
rect 1288 356 1304 390
rect 1451 351 1485 367
rect 691 296 725 312
rect 862 296 900 321
rect 881 287 900 296
rect 1003 296 1037 312
rect 691 228 725 262
rect 691 160 725 180
rect 847 228 881 262
rect 847 160 881 194
rect 847 110 881 126
rect 1161 296 1199 321
rect 1193 287 1199 296
rect 1607 351 1641 367
rect 1763 351 1797 367
rect 1315 296 1349 312
rect 1003 228 1037 262
rect 1003 160 1037 180
rect 691 70 725 108
rect 1159 228 1193 262
rect 1159 160 1193 194
rect 1159 110 1193 126
rect 1315 228 1349 262
rect 1315 160 1349 180
rect 1003 70 1037 108
rect 1315 70 1349 108
rect 172 36 350 61
rect 384 36 423 70
rect 457 36 496 70
rect 530 36 569 70
rect 603 36 642 70
rect 676 36 715 70
rect 749 36 788 70
rect 822 36 862 70
rect 896 36 936 70
rect 970 36 1010 70
rect 1044 36 1084 70
rect 1118 36 1158 70
rect 1192 36 1232 70
rect 1266 36 1306 70
rect 1340 61 1349 70
rect 1451 283 1485 317
rect 1641 317 1652 339
rect 1614 305 1652 317
rect 1919 351 1953 367
rect 1451 215 1485 249
rect 1451 147 1485 180
rect 1451 61 1485 108
rect 1607 283 1641 305
rect 1607 215 1641 249
rect 1607 147 1641 181
rect 1607 97 1641 113
rect 1763 283 1797 317
rect 2044 351 2078 367
rect 1953 317 1957 339
rect 1919 305 1957 317
rect 1763 215 1797 249
rect 1763 147 1797 180
rect 1763 61 1797 108
rect 1919 283 1953 305
rect 1919 215 1953 249
rect 1919 147 1953 181
rect 1919 97 1953 113
rect 2044 283 2078 317
rect 2200 351 2234 367
rect 2200 294 2234 317
rect 2216 283 2254 294
rect 2234 260 2254 283
rect 2044 215 2078 249
rect 2044 142 2078 180
rect 2200 215 2234 249
rect 2200 165 2234 181
rect 1340 36 2336 61
rect 172 20 2336 36
rect 172 -14 196 20
rect 230 -14 269 20
rect 303 -14 342 20
rect 376 -14 415 20
rect 449 -14 488 20
rect 522 -14 561 20
rect 595 -14 634 20
rect 668 -14 706 20
rect 740 -14 778 20
rect 812 -14 850 20
rect 884 -14 922 20
rect 956 -14 994 20
rect 1028 -14 1066 20
rect 1100 -14 1138 20
rect 1172 -14 1210 20
rect 1244 -14 1282 20
rect 1316 -14 2336 20
rect 172 -29 2336 -14
<< viali >>
rect 134 1386 146 1420
rect 146 1386 168 1420
rect 207 1386 218 1420
rect 218 1386 241 1420
rect 280 1386 290 1420
rect 290 1386 314 1420
rect 354 1386 362 1420
rect 362 1386 388 1420
rect 428 1386 434 1420
rect 434 1386 462 1420
rect 502 1386 506 1420
rect 506 1386 536 1420
rect 576 1386 577 1420
rect 577 1386 610 1420
rect 650 1386 682 1420
rect 682 1386 684 1420
rect 724 1386 753 1420
rect 753 1386 758 1420
rect 202 1270 218 1304
rect 218 1270 236 1304
rect 302 1270 320 1304
rect 320 1270 336 1304
rect 553 1270 556 1304
rect 556 1270 587 1304
rect 653 1270 658 1304
rect 658 1270 687 1304
rect 118 1243 152 1247
rect 118 1213 124 1243
rect 124 1213 152 1243
rect 118 1114 124 1148
rect 124 1114 152 1148
rect 462 1148 496 1154
rect 462 1120 496 1148
rect 552 1114 556 1148
rect 556 1114 586 1148
rect 627 1114 658 1148
rect 658 1114 661 1148
rect 118 1019 124 1049
rect 124 1019 152 1049
rect 118 1015 152 1019
rect 462 1053 496 1079
rect 462 1045 496 1053
rect 830 1193 864 1227
rect 905 1193 939 1227
rect 929 1029 963 1063
rect 1004 1059 1015 1063
rect 1015 1059 1038 1063
rect 1004 1029 1038 1059
rect 553 992 587 993
rect 653 992 687 993
rect 202 958 218 992
rect 218 958 236 992
rect 302 958 320 992
rect 320 958 336 992
rect 553 959 556 992
rect 556 959 587 992
rect 653 959 658 992
rect 658 959 687 992
rect 1429 1178 1463 1212
rect 1501 1178 1535 1212
rect 1228 1106 1262 1130
rect 1228 1096 1262 1106
rect 1300 1096 1334 1130
rect 1900 1178 1934 1212
rect 1665 1096 1699 1130
rect 1972 1178 2006 1212
rect 1737 1096 1771 1130
rect 2100 1096 2134 1130
rect 2172 1106 2206 1130
rect 2172 1096 2206 1106
rect 1007 907 1041 941
rect 1082 907 1116 941
rect 303 778 337 812
rect 217 634 251 654
rect 217 620 251 634
rect 217 566 251 582
rect 217 548 251 566
rect 475 778 509 812
rect 303 736 337 740
rect 303 706 337 736
rect 389 634 423 654
rect 389 620 423 634
rect 389 566 423 582
rect 389 548 423 566
rect 647 778 681 812
rect 475 736 509 740
rect 475 706 509 736
rect 561 634 595 654
rect 561 620 595 634
rect 561 566 595 582
rect 561 548 595 566
rect 819 778 853 812
rect 647 736 681 740
rect 647 706 681 736
rect 733 634 767 654
rect 733 620 767 634
rect 733 566 767 582
rect 733 548 767 566
rect 819 736 853 740
rect 819 706 853 736
rect 905 634 939 654
rect 905 620 939 634
rect 905 566 939 582
rect 905 548 939 566
rect 290 466 312 500
rect 312 466 324 500
rect 397 466 426 500
rect 426 466 431 500
rect 504 466 534 500
rect 534 466 538 500
rect 622 466 656 500
rect 728 466 730 500
rect 730 466 762 500
rect 834 466 844 500
rect 844 466 868 500
rect 1429 909 1463 943
rect 1190 761 1224 795
rect 1501 909 1535 943
rect 1262 761 1296 795
rect 1900 906 1934 940
rect 1972 906 2006 940
rect 1665 761 1699 795
rect 1737 761 1771 795
rect 2097 761 2131 795
rect 2169 770 2172 795
rect 2172 770 2203 795
rect 2169 761 2203 770
rect 1025 452 1059 486
rect 1100 452 1134 486
rect 1533 517 1567 525
rect 1533 491 1567 517
rect 1533 449 1567 453
rect 1533 419 1567 449
rect 1689 517 1723 525
rect 1689 491 1723 517
rect 1689 449 1723 453
rect 1689 419 1723 449
rect 1845 517 1879 525
rect 1845 491 1879 517
rect 1845 449 1879 453
rect 1845 419 1879 449
rect 2120 517 2154 535
rect 2120 501 2125 517
rect 2125 501 2154 517
rect 2120 449 2154 463
rect 2120 429 2125 449
rect 2125 429 2154 449
rect 804 390 838 395
rect 882 390 916 395
rect 960 390 994 395
rect 1038 390 1072 395
rect 1116 390 1150 395
rect 1194 390 1228 395
rect 804 361 823 390
rect 823 361 838 390
rect 882 361 894 390
rect 894 361 916 390
rect 960 361 966 390
rect 966 361 994 390
rect 1038 361 1072 390
rect 1116 361 1144 390
rect 1144 361 1150 390
rect 1194 361 1216 390
rect 1216 361 1228 390
rect 828 296 862 321
rect 828 287 847 296
rect 847 287 862 296
rect 900 287 934 321
rect 691 194 725 214
rect 691 180 725 194
rect 691 126 725 142
rect 691 108 725 126
rect 1127 296 1161 321
rect 1127 287 1159 296
rect 1159 287 1161 296
rect 1199 287 1233 321
rect 1003 194 1037 214
rect 1003 180 1037 194
rect 1003 126 1037 142
rect 1003 108 1037 126
rect 1315 194 1349 214
rect 1315 180 1349 194
rect 1315 126 1349 142
rect 1315 108 1349 126
rect 350 36 384 70
rect 423 36 457 70
rect 496 36 530 70
rect 569 36 603 70
rect 642 36 676 70
rect 715 36 749 70
rect 788 36 822 70
rect 862 36 896 70
rect 936 36 970 70
rect 1010 36 1044 70
rect 1084 36 1118 70
rect 1158 36 1192 70
rect 1232 36 1266 70
rect 1306 36 1340 70
rect 1580 317 1607 339
rect 1607 317 1614 339
rect 1580 305 1614 317
rect 1652 305 1686 339
rect 1451 181 1485 214
rect 1451 180 1485 181
rect 1451 113 1485 142
rect 1451 108 1485 113
rect 1885 305 1919 339
rect 1957 305 1991 339
rect 1763 181 1797 214
rect 1763 180 1797 181
rect 1763 113 1797 142
rect 1763 108 1797 113
rect 2182 283 2216 294
rect 2182 260 2200 283
rect 2200 260 2216 283
rect 2254 260 2288 294
rect 2044 181 2078 214
rect 2044 180 2078 181
rect 2044 108 2078 142
<< metal1 >>
rect 122 1420 874 1426
rect 122 1386 134 1420
rect 168 1386 207 1420
rect 241 1386 280 1420
rect 314 1386 354 1420
rect 388 1386 428 1420
rect 462 1386 502 1420
rect 536 1386 576 1420
rect 610 1386 650 1420
rect 684 1386 724 1420
rect 758 1386 874 1420
rect 122 1380 874 1386
tri 147 1337 190 1380 ne
rect 190 1352 874 1380
rect 190 1337 806 1352
tri 806 1337 821 1352 nw
rect 190 1310 779 1337
tri 779 1310 806 1337 nw
rect 190 1304 763 1310
rect 190 1270 202 1304
rect 236 1270 302 1304
rect 336 1270 553 1304
rect 587 1270 653 1304
rect 687 1294 763 1304
tri 763 1294 779 1310 nw
rect 687 1270 733 1294
rect 190 1264 733 1270
tri 733 1264 763 1294 nw
tri 1098 1264 1128 1294 se
rect 1128 1288 2258 1294
rect 1128 1264 2206 1288
rect 190 1259 728 1264
tri 728 1259 733 1264 nw
tri 1093 1259 1098 1264 se
rect 1098 1259 2206 1264
rect 112 1247 158 1259
rect 112 1213 118 1247
rect 152 1213 158 1247
rect 112 1148 158 1213
rect 112 1114 118 1148
rect 152 1114 158 1148
rect 112 1049 158 1114
rect 112 1015 118 1049
rect 152 1015 158 1049
rect 112 922 158 1015
rect 190 1236 705 1259
tri 705 1236 728 1259 nw
tri 1070 1236 1093 1259 se
rect 1093 1254 2206 1259
rect 1093 1236 1128 1254
tri 1128 1236 1146 1254 nw
rect 190 1233 702 1236
tri 702 1233 705 1236 nw
tri 1067 1233 1070 1236 se
rect 1070 1233 1110 1236
rect 190 1230 699 1233
tri 699 1230 702 1233 nw
rect 190 1227 368 1230
tri 368 1227 371 1230 nw
rect 818 1227 951 1233
rect 190 992 348 1227
tri 348 1207 368 1227 nw
rect 818 1193 830 1227
rect 864 1193 905 1227
rect 939 1193 951 1227
tri 1052 1218 1067 1233 se
rect 1067 1218 1110 1233
tri 1110 1218 1128 1236 nw
rect 2206 1224 2258 1236
rect 2034 1218 2040 1221
tri 1046 1212 1052 1218 se
rect 1052 1212 1104 1218
tri 1104 1212 1110 1218 nw
tri 1147 1212 1153 1218 se
rect 1153 1212 2040 1218
rect 818 1187 951 1193
tri 1021 1187 1046 1212 se
rect 1046 1187 1070 1212
tri 1012 1178 1021 1187 se
rect 1021 1178 1070 1187
tri 1070 1178 1104 1212 nw
tri 1120 1185 1147 1212 se
rect 1147 1185 1429 1212
rect 1120 1178 1429 1185
rect 1463 1178 1501 1212
rect 1535 1178 1900 1212
rect 1934 1178 1972 1212
rect 2006 1178 2040 1212
tri 1006 1172 1012 1178 se
rect 1012 1172 1064 1178
tri 1064 1172 1070 1178 nw
rect 1120 1172 2040 1178
tri 1000 1166 1006 1172 se
rect 1006 1166 1040 1172
rect 456 1154 502 1166
tri 988 1154 1000 1166 se
rect 1000 1154 1040 1166
rect 456 1120 462 1154
rect 496 1120 502 1154
rect 456 1079 502 1120
rect 540 1148 673 1154
tri 982 1148 988 1154 se
rect 988 1148 1040 1154
tri 1040 1148 1064 1172 nw
rect 1120 1169 1209 1172
tri 1209 1169 1212 1172 nw
rect 2034 1169 2040 1172
rect 2092 1169 2104 1221
rect 2156 1169 2162 1221
rect 1120 1148 1188 1169
tri 1188 1148 1209 1169 nw
rect 2206 1166 2258 1172
rect 540 1114 552 1148
rect 586 1114 627 1148
rect 661 1136 1028 1148
tri 1028 1136 1040 1148 nw
rect 661 1130 1022 1136
tri 1022 1130 1028 1136 nw
rect 661 1114 1000 1130
rect 540 1108 1000 1114
tri 1000 1108 1022 1130 nw
tri 1116 1096 1120 1100 se
rect 1120 1096 1180 1148
tri 1180 1140 1188 1148 nw
tri 1110 1090 1116 1096 se
rect 1116 1090 1180 1096
rect 1216 1130 2218 1136
rect 1216 1096 1228 1130
rect 1262 1096 1300 1130
rect 1334 1096 1665 1130
rect 1699 1096 1737 1130
rect 1771 1096 2100 1130
rect 2134 1096 2172 1130
rect 2206 1096 2218 1130
rect 1216 1090 2218 1096
rect 456 1045 462 1079
rect 496 1074 502 1079
tri 1094 1074 1110 1090 se
rect 1110 1076 1180 1090
rect 1110 1074 1178 1076
tri 1178 1074 1180 1076 nw
tri 2096 1074 2112 1090 ne
rect 2112 1074 2176 1090
rect 496 1063 1160 1074
rect 496 1045 929 1063
rect 456 1029 929 1045
rect 963 1029 1004 1063
rect 1038 1056 1160 1063
tri 1160 1056 1178 1074 nw
tri 2112 1056 2130 1074 ne
rect 1038 1029 1132 1056
rect 456 1028 1132 1029
tri 1132 1028 1160 1056 nw
rect 917 1023 1050 1028
rect 1614 1010 1642 1038
rect 541 993 699 999
rect 541 992 553 993
rect 190 958 202 992
rect 236 958 302 992
rect 336 959 553 992
rect 587 959 653 993
rect 687 959 699 993
rect 336 958 699 959
rect 190 952 348 958
rect 541 953 699 958
tri 1124 947 1126 949 se
rect 1126 947 1547 949
rect 995 946 1547 947
rect 995 943 2018 946
rect 995 941 1429 943
tri 158 922 169 933 sw
rect 112 911 292 922
tri 112 907 116 911 ne
rect 116 907 292 911
tri 116 906 117 907 ne
rect 117 906 292 907
tri 117 901 122 906 ne
rect 122 901 292 906
tri 122 900 123 901 ne
rect 123 900 292 901
tri 123 872 151 900 ne
rect 151 872 292 900
tri 151 870 153 872 ne
rect 153 870 292 872
rect 344 870 356 922
rect 408 870 414 922
rect 995 907 1007 941
rect 1041 907 1082 941
rect 1116 909 1429 941
rect 1463 909 1501 943
rect 1535 940 2018 943
rect 1535 909 1900 940
rect 1116 907 1900 909
rect 995 906 1900 907
rect 1934 906 1972 940
rect 2006 906 2018 940
rect 995 903 2018 906
rect 995 901 1144 903
tri 1144 901 1146 903 nw
rect 1547 900 2018 903
tri 2119 900 2130 911 se
rect 2130 900 2176 1074
tri 2176 1056 2210 1090 nw
tri 567 872 595 900 se
rect 595 872 903 900
tri 903 872 931 900 sw
tri 2091 872 2119 900 se
rect 2119 891 2176 900
rect 2119 872 2157 891
tri 2157 872 2176 891 nw
tri 565 870 567 872 se
rect 567 870 2139 872
tri 529 834 565 870 se
rect 565 854 2139 870
tri 2139 854 2157 872 nw
rect 565 834 595 854
tri 595 834 615 854 nw
tri 883 834 903 854 ne
rect 903 834 2115 854
tri 519 824 529 834 se
rect 529 824 585 834
tri 585 824 595 834 nw
tri 903 830 907 834 ne
rect 907 830 2115 834
tri 2115 830 2139 854 nw
rect 297 812 573 824
tri 573 812 585 824 nw
rect 641 812 859 824
rect 297 778 303 812
rect 337 778 475 812
rect 509 778 539 812
tri 539 778 573 812 nw
rect 641 778 647 812
rect 681 778 819 812
rect 853 801 859 812
tri 859 801 879 821 sw
rect 853 795 2215 801
rect 853 778 1190 795
rect 297 761 522 778
tri 522 761 539 778 nw
rect 641 763 1190 778
rect 297 740 515 761
tri 515 754 522 761 nw
rect 297 706 303 740
rect 337 706 475 740
rect 509 706 515 740
rect 297 694 515 706
rect 641 740 687 763
rect 641 706 647 740
rect 681 706 687 740
rect 641 694 687 706
rect 813 761 1190 763
rect 1224 761 1262 795
rect 1296 761 1665 795
rect 1699 761 1737 795
rect 1771 761 2097 795
rect 2131 761 2169 795
rect 2203 761 2215 795
rect 813 755 2215 761
rect 813 740 859 755
rect 813 706 819 740
rect 853 706 859 740
rect 813 694 859 706
rect 150 654 945 666
rect 150 620 217 654
rect 251 620 389 654
rect 423 620 561 654
rect 595 620 733 654
rect 767 620 905 654
rect 939 620 945 654
rect 150 582 945 620
rect -2220 361 -1967 574
rect 150 548 217 582
rect 251 548 389 582
rect 423 548 561 582
rect 595 548 733 582
rect 767 548 905 582
rect 939 548 945 582
rect 150 536 945 548
rect 2111 541 2163 547
rect 150 535 237 536
tri 237 535 238 536 nw
rect 150 525 227 535
tri 227 525 237 535 nw
rect 1527 525 1885 537
rect 150 506 208 525
tri 208 506 227 525 nw
rect 150 500 202 506
tri 202 500 208 506 nw
rect 267 500 550 506
rect 150 423 196 500
tri 196 494 202 500 nw
rect 267 466 290 500
rect 324 466 397 500
rect 431 466 504 500
rect 538 466 550 500
rect 267 460 550 466
rect 596 500 886 506
rect 596 466 622 500
rect 656 466 728 500
rect 762 466 834 500
rect 868 466 886 500
rect 596 460 886 466
rect 1013 491 1317 492
tri 1317 491 1318 492 sw
rect 1527 491 1533 525
rect 1567 491 1689 525
rect 1723 491 1845 525
rect 1879 491 1885 525
rect 1013 486 1318 491
rect 1013 452 1025 486
rect 1059 452 1100 486
rect 1134 477 1318 486
tri 1318 477 1332 491 sw
rect 1134 463 1332 477
tri 1332 463 1346 477 sw
rect 1134 460 1346 463
tri 1346 460 1349 463 sw
rect 1134 453 1349 460
tri 1349 453 1356 460 sw
rect 1527 453 1885 491
rect 1134 452 1356 453
rect 1013 446 1356 452
tri 1297 443 1300 446 ne
rect 1300 443 1356 446
tri 1356 443 1366 453 sw
tri 196 423 216 443 sw
tri 1300 423 1320 443 ne
rect 1320 423 1366 443
tri 1366 423 1386 443 sw
tri 150 419 154 423 ne
rect 154 419 216 423
tri 216 419 220 423 sw
tri 1320 419 1324 423 ne
rect 1324 419 1386 423
tri 1386 419 1390 423 sw
rect 1527 419 1533 453
rect 1567 419 1689 453
rect 1723 419 1845 453
rect 1879 419 1885 453
tri 154 395 178 419 ne
rect 178 395 220 419
tri 220 395 244 419 sw
tri 1324 411 1332 419 ne
rect 1332 411 1390 419
tri 1390 411 1398 419 sw
tri 1332 401 1342 411 ne
rect 1342 401 1398 411
rect 792 395 1240 401
tri 178 361 212 395 ne
rect 212 361 244 395
tri 244 361 278 395 sw
rect 792 361 804 395
rect 838 361 882 395
rect 916 361 960 395
rect 994 361 1038 395
rect 1072 361 1116 395
rect 1150 361 1194 395
rect 1228 361 1240 395
rect -2145 302 -1967 361
tri 212 357 216 361 ne
rect 216 357 278 361
tri 278 357 282 361 sw
tri 216 339 234 357 ne
rect 234 339 282 357
tri 282 339 300 357 sw
rect 792 355 1240 361
tri 1342 357 1386 401 ne
rect 1386 357 1398 401
tri 1398 357 1452 411 sw
rect 1527 407 1885 419
rect 2111 475 2163 489
rect 2111 417 2163 423
rect 2206 376 2258 382
tri 1386 355 1388 357 ne
rect 1388 355 1452 357
tri 1388 345 1398 355 ne
rect 1398 345 1452 355
tri 1452 345 1464 357 sw
tri 1398 339 1404 345 ne
rect 1404 339 2003 345
tri 234 321 252 339 ne
rect 252 327 300 339
tri 300 327 312 339 sw
tri 1404 327 1416 339 ne
rect 1416 327 1580 339
rect 252 321 1245 327
tri 252 302 271 321 ne
rect 271 302 828 321
rect -2145 292 -1652 302
tri -1652 292 -1642 302 sw
tri -1528 292 -1518 302 se
rect -1518 292 -1312 302
rect -2145 111 -1312 292
tri 271 291 282 302 ne
rect 282 291 828 302
tri 282 287 286 291 ne
rect 286 287 828 291
rect 862 287 900 321
rect 934 287 1127 321
rect 1161 287 1199 321
rect 1233 287 1245 321
tri 1416 305 1438 327 ne
rect 1438 305 1580 327
rect 1614 305 1652 339
rect 1686 305 1885 339
rect 1919 305 1957 339
rect 1991 305 2003 339
tri 1438 299 1444 305 ne
rect 1444 299 2003 305
rect 2206 312 2258 324
tri 286 281 292 287 ne
rect 292 281 1245 287
rect 2170 294 2206 300
rect 2258 294 2300 300
rect 2170 260 2182 294
rect 2288 260 2300 294
rect 2170 254 2300 260
tri 253 214 265 226 se
rect 265 214 2163 226
tri 219 180 253 214 se
rect 253 180 691 214
rect 725 180 1003 214
rect 1037 180 1315 214
rect 1349 180 1451 214
rect 1485 180 1763 214
rect 1797 180 2044 214
rect 2078 180 2163 214
tri 181 142 219 180 se
rect 219 142 2163 180
tri 180 141 181 142 se
rect 181 141 691 142
tri -23 111 7 141 se
rect 7 111 691 141
tri -26 108 -23 111 se
rect -23 108 691 111
rect 725 108 1003 142
rect 1037 108 1315 142
rect 1349 108 1451 142
rect 1485 108 1763 142
rect 1797 108 2044 142
rect 2078 108 2163 142
tri -38 96 -26 108 se
rect -26 96 2163 108
tri -58 76 -38 96 se
rect -38 76 2163 96
tri -64 70 -58 76 se
rect -58 70 2163 76
tri -98 36 -64 70 se
rect -64 36 350 70
rect 384 36 423 70
rect 457 36 496 70
rect 530 36 569 70
rect 603 36 642 70
rect 676 36 715 70
rect 749 36 788 70
rect 822 36 862 70
rect 896 36 936 70
rect 970 36 1010 70
rect 1044 36 1084 70
rect 1118 36 1158 70
rect 1192 36 1232 70
rect 1266 36 1306 70
rect 1340 36 2163 70
tri -104 30 -98 36 se
rect -98 30 2163 36
tri -165 -31 -104 30 se
rect -104 -31 26 30
tri 26 -31 87 30 nw
tri -967 -140 -858 -31 se
rect -858 -140 -83 -31
tri -83 -140 26 -31 nw
rect -1219 -141 -84 -140
tri -84 -141 -83 -140 nw
rect -1219 -193 -1212 -141
rect -1160 -193 -1094 -141
rect -1042 -193 -139 -141
rect -1219 -196 -139 -193
tri -139 -196 -84 -141 nw
rect -1219 -227 -904 -196
rect -1219 -279 -1212 -227
rect -1160 -279 -1094 -227
rect -1042 -279 -904 -227
tri -904 -279 -821 -196 nw
rect -1219 -282 -907 -279
tri -907 -282 -904 -279 nw
rect -1219 -283 -1001 -282
<< via1 >>
rect 2206 1236 2258 1288
rect 2040 1169 2092 1221
rect 2104 1169 2156 1221
rect 2206 1172 2258 1224
rect 292 870 344 922
rect 356 870 408 922
rect 2111 535 2163 541
rect 2111 501 2120 535
rect 2120 501 2154 535
rect 2154 501 2163 535
rect 2111 489 2163 501
rect 2111 463 2163 475
rect 2111 429 2120 463
rect 2120 429 2154 463
rect 2154 429 2163 463
rect 2111 423 2163 429
rect 2206 324 2258 376
rect 2206 294 2258 312
rect 2206 260 2216 294
rect 2216 260 2254 294
rect 2254 260 2258 294
rect -1212 -193 -1160 -141
rect -1094 -193 -1042 -141
rect -1212 -279 -1160 -227
rect -1094 -279 -1042 -227
<< metal2 >>
rect 2206 1288 2258 1294
rect 2206 1224 2258 1236
rect 2034 1169 2040 1221
rect 2092 1169 2104 1221
rect 2156 1169 2163 1221
rect 286 870 292 922
rect 344 870 356 922
rect 408 870 414 922
rect 2111 541 2163 1169
rect 2111 475 2163 489
rect 2111 415 2163 423
rect 2206 376 2258 1172
rect 2206 312 2258 324
rect 2206 254 2258 260
rect -1218 -193 -1212 -141
rect -1160 -142 -1094 -141
rect -1218 -198 -1208 -193
rect -1152 -198 -1101 -142
rect -1042 -193 -1036 -141
rect -1045 -198 -1036 -193
rect -1218 -226 -1036 -198
rect -1218 -227 -1208 -226
rect -1218 -279 -1212 -227
rect -1217 -282 -1208 -279
rect -1152 -282 -1101 -226
rect -1045 -227 -1036 -226
rect -1042 -279 -1036 -227
rect -1045 -282 -1036 -279
<< via2 >>
rect -1208 -193 -1160 -142
rect -1160 -193 -1152 -142
rect -1208 -198 -1152 -193
rect -1101 -193 -1094 -142
rect -1094 -193 -1045 -142
rect -1101 -198 -1045 -193
rect -1208 -227 -1152 -226
rect -1208 -279 -1160 -227
rect -1160 -279 -1152 -227
rect -1208 -282 -1152 -279
rect -1101 -227 -1045 -226
rect -1101 -279 -1094 -227
rect -1094 -279 -1045 -227
rect -1101 -282 -1045 -279
<< metal3 >>
rect -1213 -142 -1040 -137
rect -1213 -198 -1208 -142
rect -1152 -198 -1101 -142
rect -1045 -198 -1040 -142
rect -1213 -226 -1040 -198
rect -1213 -282 -1208 -226
rect -1152 -282 -1101 -226
rect -1045 -282 -1040 -226
rect -1213 -287 -1040 -282
use sky130_fd_pr__nfet_01v8__example_55959141808468  sky130_fd_pr__nfet_01v8__example_55959141808468_0
timestamp 1640697850
transform -1 0 2161 0 1 758
box -28 0 916 97
use sky130_fd_pr__nfet_01v8__example_55959141808467  sky130_fd_pr__nfet_01v8__example_55959141808467_0
timestamp 1640697850
transform -1 0 894 0 -1 748
box -28 0 316 97
use sky130_fd_pr__nfet_01v8__example_55959141808466  sky130_fd_pr__nfet_01v8__example_55959141808466_0
timestamp 1640697850
transform -1 0 550 0 -1 748
box -28 0 316 97
use sky130_fd_pr__nfet_01v8__example_55959141808465  sky130_fd_pr__nfet_01v8__example_55959141808465_0
timestamp 1640697850
transform 1 0 2089 0 -1 363
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808464  sky130_fd_pr__nfet_01v8__example_55959141808464_0
timestamp 1640697850
transform -1 0 2161 0 -1 1288
box -28 0 916 97
use sky130_fd_pr__nfet_01v8__example_55959141808463  sky130_fd_pr__nfet_01v8__example_55959141808463_0
timestamp 1640697850
transform 1 0 736 0 1 114
box -28 0 596 97
use sky130_fd_pr__nfet_01v8__example_55959141808461  sky130_fd_pr__nfet_01v8__example_55959141808461_0
timestamp 1640697850
transform 1 0 1496 0 -1 363
box -28 0 440 131
use sky130_fd_pr__pfet_01v8__example_55959141808460  sky130_fd_pr__pfet_01v8__example_55959141808460_0
timestamp 1640697850
transform 0 1 817 1 0 1159
box -28 0 128 63
use sky130_fd_pr__pfet_01v8__example_55959141808460  sky130_fd_pr__pfet_01v8__example_55959141808460_1
timestamp 1640697850
transform 0 1 817 1 0 1003
box -28 0 128 63
use sky130_fd_pr__pfet_01v8__example_55959141808460  sky130_fd_pr__pfet_01v8__example_55959141808460_2
timestamp 1640697850
transform 0 1 544 1 0 1159
box -28 0 128 63
use sky130_fd_pr__pfet_01v8__example_55959141808460  sky130_fd_pr__pfet_01v8__example_55959141808460_3
timestamp 1640697850
transform 0 1 544 1 0 1003
box -28 0 128 63
use sky130_fd_pr__pfet_01v8__example_55959141808458  sky130_fd_pr__pfet_01v8__example_55959141808458_0
timestamp 1640697850
transform 0 1 206 -1 0 1259
box -28 0 284 63
<< labels >>
flabel comment s 741 1066 741 1066 0 FreeSans 600 0 0 0 FBK_N
flabel metal1 s 771 472 799 500 3 FreeSans 280 0 0 0 IN_B
port 1 nsew
flabel metal1 s 2181 263 2209 291 3 FreeSans 280 0 0 0 OUT_H
port 2 nsew
flabel metal1 s 127 1006 155 1034 3 FreeSans 280 0 0 0 RST_H_N
port 3 nsew
flabel metal1 s 463 1341 491 1369 3 FreeSans 280 0 0 0 VPWR_HV
port 4 nsew
flabel metal1 s 1980 157 2008 185 3 FreeSans 280 0 0 0 VGND
port 5 nsew
flabel metal1 s 966 357 994 385 3 FreeSans 280 180 0 0 RST_H_N
port 3 nsew
flabel metal1 s 1668 455 1696 483 3 FreeSans 280 0 0 0 RST_H
port 6 nsew
flabel metal1 s 422 471 450 499 3 FreeSans 280 0 0 0 IN
port 7 nsew
flabel metal1 s 1614 1010 1642 1038 3 FreeSans 280 0 0 0 VPWR_LV
port 8 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 48718928
string GDS_START 48688374
<< end >>
