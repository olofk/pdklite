magic
tech sky130A
magscale 1 2
timestamp 1619729575
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 371 323 405 493
rect 539 323 573 493
rect 707 323 741 493
rect 875 323 909 493
rect 371 289 909 323
rect 28 215 248 255
rect 858 181 909 289
rect 371 147 909 181
rect 371 51 405 147
rect 539 51 573 147
rect 707 51 741 147
rect 875 51 909 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 19 323 85 493
rect 119 367 153 527
rect 187 323 253 493
rect 287 367 321 527
rect 439 367 505 527
rect 607 367 673 527
rect 775 367 841 527
rect 19 289 319 323
rect 943 297 1009 527
rect 284 249 319 289
rect 284 215 809 249
rect 284 181 319 215
rect 35 147 319 181
rect 35 51 69 147
rect 103 17 169 113
rect 203 52 237 147
rect 271 17 337 113
rect 439 17 505 113
rect 607 17 673 113
rect 775 17 841 113
rect 943 17 1009 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 28 215 248 255 6 A
port 1 nsew signal input
rlabel locali s 875 323 909 493 6 X
port 6 nsew signal output
rlabel locali s 875 51 909 147 6 X
port 6 nsew signal output
rlabel locali s 858 181 909 289 6 X
port 6 nsew signal output
rlabel locali s 707 323 741 493 6 X
port 6 nsew signal output
rlabel locali s 707 51 741 147 6 X
port 6 nsew signal output
rlabel locali s 539 323 573 493 6 X
port 6 nsew signal output
rlabel locali s 539 51 573 147 6 X
port 6 nsew signal output
rlabel locali s 371 323 405 493 6 X
port 6 nsew signal output
rlabel locali s 371 289 909 323 6 X
port 6 nsew signal output
rlabel locali s 371 147 909 181 6 X
port 6 nsew signal output
rlabel locali s 371 51 405 147 6 X
port 6 nsew signal output
rlabel metal1 s 0 -48 1104 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2351516
string GDS_START 2342684
<< end >>
