magic
tech sky130A
magscale 1 2
timestamp 1619729575
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 88 153 158 327
rect 196 309 432 343
rect 196 164 252 309
rect 196 130 416 164
rect 214 51 248 130
rect 382 51 416 130
rect 573 199 617 265
rect 669 151 711 265
rect 763 147 829 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 417 69 493
rect 103 451 169 527
rect 282 451 348 527
rect 450 451 516 527
rect 695 451 761 527
rect 927 451 993 527
rect 17 383 980 417
rect 17 117 52 383
rect 476 309 909 343
rect 476 249 510 309
rect 288 215 510 249
rect 17 51 69 117
rect 114 17 180 94
rect 282 17 348 94
rect 476 157 510 215
rect 476 123 593 157
rect 946 199 980 383
rect 559 94 593 123
rect 878 94 993 162
rect 457 17 523 89
rect 559 60 993 94
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel locali s 88 153 158 327 6 A_N
port 1 nsew signal input
rlabel locali s 763 147 829 265 6 B
port 2 nsew signal input
rlabel locali s 669 151 711 265 6 C
port 3 nsew signal input
rlabel locali s 573 199 617 265 6 D
port 4 nsew signal input
rlabel locali s 382 51 416 130 6 X
port 9 nsew signal output
rlabel locali s 214 51 248 130 6 X
port 9 nsew signal output
rlabel locali s 196 309 432 343 6 X
port 9 nsew signal output
rlabel locali s 196 164 252 309 6 X
port 9 nsew signal output
rlabel locali s 196 130 416 164 6 X
port 9 nsew signal output
rlabel metal1 s 0 -48 1012 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1050 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 260114
string GDS_START 252436
<< end >>
