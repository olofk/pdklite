magic
tech sky130A
magscale 1 2
timestamp 1619729571
<< checkpaint >>
rect -1298 -1308 3782 1852
<< nwell >>
rect -38 261 2522 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 80 47 110 175
rect 175 47 205 177
rect 404 49 434 177
rect 488 49 518 177
rect 696 47 726 175
rect 829 49 859 177
rect 1016 47 1046 177
rect 1114 49 1144 177
rect 1313 49 1343 177
rect 1398 49 1428 177
rect 1680 49 1710 177
rect 1768 49 1798 177
rect 1994 49 2024 177
rect 2089 47 2119 177
rect 2277 49 2307 177
rect 2372 47 2402 177
<< scpmoshvt >>
rect 80 297 110 497
rect 180 297 210 497
rect 404 297 434 465
rect 488 297 518 465
rect 705 297 735 465
rect 802 322 832 490
rect 1012 297 1042 497
rect 1114 297 1144 497
rect 1302 297 1332 465
rect 1386 297 1416 465
rect 1690 315 1720 483
rect 1774 315 1804 483
rect 2000 297 2030 497
rect 2084 297 2114 497
rect 2277 297 2307 497
rect 2361 297 2391 497
<< ndiff >>
rect 125 175 175 177
rect 28 161 80 175
rect 28 127 36 161
rect 70 127 80 161
rect 28 93 80 127
rect 28 59 36 93
rect 70 59 80 93
rect 28 47 80 59
rect 110 93 175 175
rect 110 59 126 93
rect 160 59 175 93
rect 110 47 175 59
rect 205 161 404 177
rect 205 127 215 161
rect 249 127 404 161
rect 205 93 404 127
rect 205 59 215 93
rect 249 59 360 93
rect 394 59 404 93
rect 205 49 404 59
rect 434 161 488 177
rect 434 127 444 161
rect 478 127 488 161
rect 434 49 488 127
rect 518 165 586 177
rect 763 175 829 177
rect 518 131 544 165
rect 578 131 586 165
rect 518 49 586 131
rect 640 101 696 175
rect 640 67 648 101
rect 682 67 696 101
rect 205 47 318 49
rect 640 47 696 67
rect 726 169 829 175
rect 726 135 785 169
rect 819 135 829 169
rect 726 49 829 135
rect 859 106 909 177
rect 964 163 1016 177
rect 964 129 972 163
rect 1006 129 1016 163
rect 964 121 1016 129
rect 859 95 911 106
rect 859 61 869 95
rect 903 61 911 95
rect 859 49 911 61
rect 726 47 798 49
rect 965 47 1016 121
rect 1046 161 1114 177
rect 1046 127 1056 161
rect 1090 127 1114 161
rect 1046 93 1114 127
rect 1046 59 1056 93
rect 1090 59 1114 93
rect 1046 49 1114 59
rect 1144 133 1196 177
rect 1144 99 1154 133
rect 1188 99 1196 133
rect 1144 49 1196 99
rect 1261 114 1313 177
rect 1261 80 1269 114
rect 1303 80 1313 114
rect 1261 49 1313 80
rect 1343 169 1398 177
rect 1343 135 1353 169
rect 1387 135 1398 169
rect 1343 49 1398 135
rect 1428 169 1489 177
rect 1428 135 1438 169
rect 1472 135 1489 169
rect 1428 49 1489 135
rect 1589 161 1680 177
rect 1589 127 1604 161
rect 1638 127 1680 161
rect 1589 93 1680 127
rect 1589 59 1604 93
rect 1638 59 1680 93
rect 1589 49 1680 59
rect 1710 153 1768 177
rect 1710 119 1724 153
rect 1758 119 1768 153
rect 1710 49 1768 119
rect 1798 165 1994 177
rect 1798 131 1948 165
rect 1982 131 1994 165
rect 1798 97 1994 131
rect 1798 63 1948 97
rect 1982 63 1994 97
rect 1798 49 1994 63
rect 2024 97 2089 177
rect 2024 63 2040 97
rect 2074 63 2089 97
rect 2024 49 2089 63
rect 1046 47 1096 49
rect 2039 47 2089 49
rect 2119 165 2171 177
rect 2119 131 2129 165
rect 2163 131 2171 165
rect 2119 97 2171 131
rect 2119 63 2129 97
rect 2163 63 2171 97
rect 2119 47 2171 63
rect 2225 127 2277 177
rect 2225 93 2233 127
rect 2267 93 2277 127
rect 2225 49 2277 93
rect 2307 95 2372 177
rect 2307 61 2317 95
rect 2351 61 2372 95
rect 2307 49 2372 61
rect 2322 47 2372 49
rect 2402 163 2457 177
rect 2402 129 2415 163
rect 2449 129 2457 163
rect 2402 95 2457 129
rect 2402 61 2415 95
rect 2449 61 2457 95
rect 2402 47 2457 61
<< pdiff >>
rect 28 479 80 497
rect 28 445 36 479
rect 70 445 80 479
rect 28 411 80 445
rect 28 377 36 411
rect 70 377 80 411
rect 28 343 80 377
rect 28 309 36 343
rect 70 309 80 343
rect 28 297 80 309
rect 110 486 180 497
rect 110 452 120 486
rect 154 452 180 486
rect 110 297 180 452
rect 210 369 260 497
rect 638 493 688 505
rect 332 477 389 489
rect 332 443 344 477
rect 378 465 389 477
rect 378 443 404 465
rect 332 431 404 443
rect 210 350 298 369
rect 210 316 256 350
rect 290 316 298 350
rect 210 297 298 316
rect 354 297 404 431
rect 434 341 488 465
rect 434 307 444 341
rect 478 307 488 341
rect 434 297 488 307
rect 518 409 570 465
rect 518 375 528 409
rect 562 375 570 409
rect 518 297 570 375
rect 638 459 646 493
rect 680 465 688 493
rect 752 465 802 490
rect 680 459 705 465
rect 638 341 705 459
rect 638 307 654 341
rect 688 307 705 341
rect 638 297 705 307
rect 735 357 802 465
rect 735 323 745 357
rect 779 323 802 357
rect 735 322 802 323
rect 832 403 888 490
rect 832 369 842 403
rect 876 369 888 403
rect 832 322 888 369
rect 960 345 1012 497
rect 735 297 787 322
rect 960 311 968 345
rect 1002 311 1012 345
rect 960 297 1012 311
rect 1042 481 1114 497
rect 1042 447 1070 481
rect 1104 447 1114 481
rect 1042 297 1114 447
rect 1144 465 1271 497
rect 1634 475 1690 483
rect 1144 413 1302 465
rect 1144 379 1258 413
rect 1292 379 1302 413
rect 1144 345 1302 379
rect 1144 311 1154 345
rect 1188 311 1302 345
rect 1144 297 1302 311
rect 1332 341 1386 465
rect 1332 307 1342 341
rect 1376 307 1386 341
rect 1332 297 1386 307
rect 1416 409 1524 465
rect 1416 375 1478 409
rect 1512 375 1524 409
rect 1416 341 1524 375
rect 1416 307 1478 341
rect 1512 307 1524 341
rect 1634 441 1646 475
rect 1680 441 1690 475
rect 1634 407 1690 441
rect 1634 373 1646 407
rect 1680 373 1690 407
rect 1634 315 1690 373
rect 1720 425 1774 483
rect 1720 391 1730 425
rect 1764 391 1774 425
rect 1720 357 1774 391
rect 1720 323 1730 357
rect 1764 323 1774 357
rect 1720 315 1774 323
rect 1804 425 1876 483
rect 1804 391 1830 425
rect 1864 391 1876 425
rect 1804 357 1876 391
rect 1804 323 1830 357
rect 1864 323 1876 357
rect 1804 315 1876 323
rect 1930 477 2000 497
rect 1930 443 1940 477
rect 1974 443 2000 477
rect 1930 389 2000 443
rect 1930 355 1954 389
rect 1988 355 2000 389
rect 1416 297 1524 307
rect 1930 297 2000 355
rect 2030 489 2084 497
rect 2030 455 2040 489
rect 2074 455 2084 489
rect 2030 297 2084 455
rect 2114 477 2171 497
rect 2114 443 2125 477
rect 2159 443 2171 477
rect 2114 409 2171 443
rect 2114 375 2125 409
rect 2159 375 2171 409
rect 2114 341 2171 375
rect 2114 307 2125 341
rect 2159 307 2171 341
rect 2114 297 2171 307
rect 2225 480 2277 497
rect 2225 446 2233 480
rect 2267 446 2277 480
rect 2225 412 2277 446
rect 2225 378 2233 412
rect 2267 378 2277 412
rect 2225 344 2277 378
rect 2225 310 2233 344
rect 2267 310 2277 344
rect 2225 297 2277 310
rect 2307 475 2361 497
rect 2307 441 2317 475
rect 2351 441 2361 475
rect 2307 407 2361 441
rect 2307 373 2317 407
rect 2351 373 2361 407
rect 2307 297 2361 373
rect 2391 477 2448 497
rect 2391 443 2402 477
rect 2436 443 2448 477
rect 2391 409 2448 443
rect 2391 375 2402 409
rect 2436 375 2448 409
rect 2391 297 2448 375
<< ndiffc >>
rect 36 127 70 161
rect 36 59 70 93
rect 126 59 160 93
rect 215 127 249 161
rect 215 59 249 93
rect 360 59 394 93
rect 444 127 478 161
rect 544 131 578 165
rect 648 67 682 101
rect 785 135 819 169
rect 972 129 1006 163
rect 869 61 903 95
rect 1056 127 1090 161
rect 1056 59 1090 93
rect 1154 99 1188 133
rect 1269 80 1303 114
rect 1353 135 1387 169
rect 1438 135 1472 169
rect 1604 127 1638 161
rect 1604 59 1638 93
rect 1724 119 1758 153
rect 1948 131 1982 165
rect 1948 63 1982 97
rect 2040 63 2074 97
rect 2129 131 2163 165
rect 2129 63 2163 97
rect 2233 93 2267 127
rect 2317 61 2351 95
rect 2415 129 2449 163
rect 2415 61 2449 95
<< pdiffc >>
rect 36 445 70 479
rect 36 377 70 411
rect 36 309 70 343
rect 120 452 154 486
rect 344 443 378 477
rect 256 316 290 350
rect 444 307 478 341
rect 528 375 562 409
rect 646 459 680 493
rect 654 307 688 341
rect 745 323 779 357
rect 842 369 876 403
rect 968 311 1002 345
rect 1070 447 1104 481
rect 1258 379 1292 413
rect 1154 311 1188 345
rect 1342 307 1376 341
rect 1478 375 1512 409
rect 1478 307 1512 341
rect 1646 441 1680 475
rect 1646 373 1680 407
rect 1730 391 1764 425
rect 1730 323 1764 357
rect 1830 391 1864 425
rect 1830 323 1864 357
rect 1940 443 1974 477
rect 1954 355 1988 389
rect 2040 455 2074 489
rect 2125 443 2159 477
rect 2125 375 2159 409
rect 2125 307 2159 341
rect 2233 446 2267 480
rect 2233 378 2267 412
rect 2233 310 2267 344
rect 2317 441 2351 475
rect 2317 373 2351 407
rect 2402 443 2436 477
rect 2402 375 2436 409
<< poly >>
rect 80 497 110 523
rect 180 497 210 523
rect 404 465 434 491
rect 488 465 518 491
rect 705 465 735 491
rect 802 490 832 516
rect 1012 497 1042 523
rect 1114 497 1144 523
rect 80 265 110 297
rect 180 265 210 297
rect 404 265 434 297
rect 67 249 133 265
rect 67 215 85 249
rect 119 215 133 249
rect 67 199 133 215
rect 175 249 262 265
rect 175 215 218 249
rect 252 215 262 249
rect 175 199 262 215
rect 304 249 434 265
rect 304 215 314 249
rect 348 215 434 249
rect 304 199 434 215
rect 80 175 110 199
rect 175 177 205 199
rect 404 177 434 199
rect 488 265 518 297
rect 705 265 735 297
rect 802 265 832 322
rect 1302 465 1332 491
rect 1386 465 1416 491
rect 1690 483 1720 509
rect 1774 483 1804 509
rect 2000 497 2030 523
rect 2084 497 2114 523
rect 2277 497 2307 523
rect 2361 497 2391 523
rect 1690 300 1720 315
rect 1012 265 1042 297
rect 1114 265 1144 297
rect 1302 265 1332 297
rect 1386 265 1416 297
rect 1601 270 1720 300
rect 1601 265 1710 270
rect 1774 265 1804 315
rect 2000 265 2030 297
rect 2084 265 2114 297
rect 2277 265 2307 297
rect 2361 265 2391 297
rect 488 249 737 265
rect 488 215 545 249
rect 579 215 737 249
rect 488 199 737 215
rect 802 249 1144 265
rect 802 215 853 249
rect 887 215 1144 249
rect 802 199 1144 215
rect 1243 249 1343 265
rect 1243 215 1253 249
rect 1287 215 1343 249
rect 1243 199 1343 215
rect 1386 249 1710 265
rect 1386 215 1575 249
rect 1609 215 1710 249
rect 1386 199 1710 215
rect 1762 249 1822 265
rect 1762 215 1772 249
rect 1806 215 1822 249
rect 1762 199 1822 215
rect 1988 249 2042 265
rect 1988 215 1998 249
rect 2032 215 2042 249
rect 1988 199 2042 215
rect 2084 249 2307 265
rect 2084 215 2138 249
rect 2172 215 2307 249
rect 2084 199 2307 215
rect 2349 249 2403 265
rect 2349 215 2359 249
rect 2393 215 2403 249
rect 2349 199 2403 215
rect 488 177 518 199
rect 696 175 726 199
rect 829 177 859 199
rect 1016 177 1046 199
rect 1114 177 1144 199
rect 1313 177 1343 199
rect 1398 177 1428 199
rect 1680 177 1710 199
rect 1768 177 1798 199
rect 1994 177 2024 199
rect 2089 177 2119 199
rect 2277 177 2307 199
rect 2372 177 2402 199
rect 80 21 110 47
rect 175 21 205 47
rect 404 21 434 49
rect 488 21 518 49
rect 696 21 726 47
rect 829 23 859 49
rect 1016 21 1046 47
rect 1114 23 1144 49
rect 1313 23 1343 49
rect 1398 23 1428 49
rect 1680 23 1710 49
rect 1768 21 1798 49
rect 1994 23 2024 49
rect 2089 21 2119 47
rect 2277 23 2307 49
rect 2372 21 2402 47
<< polycont >>
rect 85 215 119 249
rect 218 215 252 249
rect 314 215 348 249
rect 545 215 579 249
rect 853 215 887 249
rect 1253 215 1287 249
rect 1575 215 1609 249
rect 1772 215 1806 249
rect 1998 215 2032 249
rect 2138 215 2172 249
rect 2359 215 2393 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 17 479 86 493
rect 17 445 36 479
rect 70 445 86 479
rect 17 411 86 445
rect 120 486 154 527
rect 475 477 646 493
rect 120 436 154 452
rect 188 443 344 477
rect 378 459 646 477
rect 680 459 708 493
rect 745 459 1020 493
rect 378 443 509 459
rect 17 377 36 411
rect 70 402 86 411
rect 188 402 222 443
rect 70 377 222 402
rect 17 368 222 377
rect 256 391 528 409
rect 17 343 88 368
rect 17 309 36 343
rect 70 309 88 343
rect 290 375 528 391
rect 562 375 584 409
rect 256 350 290 357
rect 17 300 88 309
rect 122 316 256 334
rect 654 341 688 459
rect 122 300 290 316
rect 393 307 444 341
rect 478 307 494 341
rect 17 161 51 300
rect 122 265 156 300
rect 85 249 156 265
rect 119 215 156 249
rect 190 249 268 255
rect 190 215 218 249
rect 252 215 268 249
rect 302 249 356 265
rect 302 215 314 249
rect 348 215 356 249
rect 85 199 156 215
rect 122 181 156 199
rect 302 187 356 215
rect 122 161 265 181
rect 17 147 36 161
rect 20 127 36 147
rect 70 127 86 161
rect 122 147 215 161
rect 20 93 86 127
rect 199 127 215 147
rect 249 127 265 161
rect 302 153 305 187
rect 339 153 356 187
rect 302 142 356 153
rect 393 255 494 307
rect 393 221 397 255
rect 431 221 494 255
rect 393 161 494 221
rect 528 289 586 323
rect 528 249 620 289
rect 528 215 545 249
rect 579 232 620 249
rect 579 215 595 232
rect 654 185 688 307
rect 745 357 779 459
rect 842 403 876 419
rect 975 413 1020 459
rect 1054 481 1120 527
rect 1054 447 1070 481
rect 1104 447 1120 481
rect 1167 459 1592 493
rect 1167 413 1201 459
rect 975 379 1201 413
rect 1242 413 1444 425
rect 1242 379 1258 413
rect 1292 391 1444 413
rect 1292 379 1308 391
rect 842 351 876 357
rect 1242 345 1276 379
rect 745 264 779 323
rect 940 323 968 345
rect 940 289 954 323
rect 1002 311 1036 345
rect 1129 311 1154 345
rect 1188 311 1276 345
rect 1342 341 1376 357
rect 988 289 1036 311
rect 940 277 1036 289
rect 745 230 819 264
rect 611 181 750 185
rect 393 127 444 161
rect 478 127 494 161
rect 528 165 750 181
rect 528 131 544 165
rect 578 151 750 165
rect 578 147 632 151
rect 578 131 605 147
rect 20 59 36 93
rect 70 59 86 93
rect 20 51 86 59
rect 126 93 160 109
rect 126 17 160 59
rect 199 93 265 127
rect 648 101 682 117
rect 199 59 215 93
rect 249 59 360 93
rect 394 67 648 93
rect 394 59 682 67
rect 199 51 682 59
rect 716 85 750 151
rect 785 169 819 230
rect 785 119 819 135
rect 853 249 903 265
rect 887 215 903 249
rect 853 187 903 215
rect 853 153 862 187
rect 896 153 903 187
rect 853 129 903 153
rect 968 199 1036 277
rect 968 163 1006 199
rect 1162 163 1196 311
rect 1322 307 1342 335
rect 968 129 972 163
rect 968 102 1006 129
rect 1040 127 1056 161
rect 1090 127 1106 161
rect 853 85 869 95
rect 716 61 869 85
rect 903 61 919 95
rect 716 51 919 61
rect 1040 93 1106 127
rect 1040 59 1056 93
rect 1090 59 1106 93
rect 1140 133 1196 163
rect 1230 255 1287 265
rect 1264 249 1287 255
rect 1230 215 1253 221
rect 1230 148 1287 215
rect 1322 185 1376 307
rect 1410 246 1444 391
rect 1478 409 1512 425
rect 1478 341 1512 375
rect 1558 344 1592 459
rect 1646 477 1990 493
rect 1646 475 1940 477
rect 1680 459 1940 475
rect 1924 443 1940 459
rect 1974 443 1990 477
rect 2024 489 2091 527
rect 2024 455 2040 489
rect 2074 455 2091 489
rect 2125 477 2167 493
rect 1646 407 1680 441
rect 1646 357 1680 373
rect 1714 391 1730 425
rect 1764 391 1780 425
rect 1714 357 1780 391
rect 1558 310 1609 344
rect 1714 323 1730 357
rect 1764 323 1780 357
rect 1478 306 1512 307
rect 1478 272 1524 306
rect 1490 258 1524 272
rect 1410 212 1456 246
rect 1490 221 1540 258
rect 1422 185 1456 212
rect 1506 187 1540 221
rect 1575 249 1609 310
rect 1575 199 1609 215
rect 1688 289 1690 323
rect 1724 306 1780 323
rect 1814 391 1830 425
rect 1864 409 1884 425
rect 1864 391 1890 409
rect 1814 357 1856 391
rect 1814 323 1830 357
rect 1864 323 1890 357
rect 1814 306 1890 323
rect 1724 289 1748 306
rect 1322 169 1387 185
rect 1322 151 1353 169
rect 1140 99 1154 133
rect 1188 99 1196 133
rect 1353 119 1387 135
rect 1422 169 1472 185
rect 1422 135 1438 169
rect 1422 119 1472 135
rect 1140 76 1196 99
rect 1253 80 1269 114
rect 1303 85 1319 114
rect 1506 85 1540 153
rect 1303 80 1540 85
rect 1040 17 1106 59
rect 1253 51 1540 80
rect 1587 161 1654 165
rect 1587 127 1604 161
rect 1638 127 1654 161
rect 1587 93 1654 127
rect 1688 153 1722 289
rect 1756 249 1782 255
rect 1756 215 1772 249
rect 1816 221 1822 255
rect 1806 215 1822 221
rect 1756 199 1822 215
rect 1688 119 1724 153
rect 1758 119 1780 153
rect 1587 59 1604 93
rect 1638 85 1654 93
rect 1856 85 1890 306
rect 1638 59 1890 85
rect 1587 51 1890 59
rect 1930 389 1990 443
rect 2159 443 2167 477
rect 2125 409 2167 443
rect 1930 355 1954 389
rect 1988 355 1990 389
rect 1930 307 1990 355
rect 2038 391 2125 409
rect 2072 375 2125 391
rect 2159 375 2167 409
rect 2072 357 2167 375
rect 2038 341 2167 357
rect 2038 307 2125 341
rect 2159 307 2167 341
rect 1930 165 1964 307
rect 2038 291 2167 307
rect 2217 480 2283 493
rect 2217 446 2233 480
rect 2267 446 2283 480
rect 2217 412 2283 446
rect 2217 378 2233 412
rect 2267 378 2283 412
rect 2217 344 2283 378
rect 2317 475 2368 527
rect 2351 441 2368 475
rect 2317 407 2368 441
rect 2351 373 2368 407
rect 2317 357 2368 373
rect 2402 477 2467 493
rect 2436 443 2467 477
rect 2402 409 2467 443
rect 2436 375 2467 409
rect 2402 357 2467 375
rect 2217 310 2233 344
rect 2267 310 2283 344
rect 2217 291 2283 310
rect 2038 265 2072 291
rect 1998 249 2072 265
rect 2032 215 2072 249
rect 2106 249 2195 255
rect 2106 215 2138 249
rect 2172 215 2195 249
rect 1998 199 2072 215
rect 2038 181 2072 199
rect 2233 187 2283 291
rect 2331 289 2338 323
rect 2372 289 2393 323
rect 2331 249 2393 289
rect 2331 215 2359 249
rect 2331 199 2393 215
rect 2038 165 2184 181
rect 1930 131 1948 165
rect 1982 131 2004 165
rect 2038 147 2129 165
rect 1930 97 2004 131
rect 2108 131 2129 147
rect 2163 131 2184 165
rect 1930 63 1948 97
rect 1982 63 2004 97
rect 1930 51 2004 63
rect 2040 97 2074 113
rect 2040 17 2074 63
rect 2108 97 2184 131
rect 2108 63 2129 97
rect 2163 63 2184 97
rect 2108 57 2184 63
rect 2233 153 2246 187
rect 2280 153 2283 187
rect 2427 165 2467 357
rect 2233 136 2283 153
rect 2399 163 2467 165
rect 2233 127 2267 136
rect 2399 129 2415 163
rect 2449 129 2467 163
rect 2233 54 2267 93
rect 2307 95 2365 111
rect 2307 61 2317 95
rect 2351 61 2365 95
rect 2307 17 2365 61
rect 2399 95 2467 129
rect 2399 61 2415 95
rect 2449 61 2467 95
rect 2399 51 2467 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 256 357 290 391
rect 305 153 339 187
rect 397 221 431 255
rect 586 289 620 323
rect 842 369 876 391
rect 842 357 876 369
rect 954 311 968 323
rect 968 311 988 323
rect 954 289 988 311
rect 862 153 896 187
rect 1230 249 1264 255
rect 1230 221 1253 249
rect 1253 221 1264 249
rect 1690 289 1724 323
rect 1856 357 1890 391
rect 1506 153 1540 187
rect 1782 249 1816 255
rect 1782 221 1806 249
rect 1806 221 1816 249
rect 2038 357 2072 391
rect 2338 289 2372 323
rect 2246 153 2280 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
<< metal1 >>
rect 0 561 2484 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 0 496 2484 527
rect 239 391 302 397
rect 239 357 256 391
rect 290 388 302 391
rect 830 391 888 397
rect 830 388 842 391
rect 290 360 842 388
rect 290 357 302 360
rect 239 351 302 357
rect 830 357 842 360
rect 876 357 888 391
rect 830 351 888 357
rect 1839 391 1902 397
rect 1839 357 1856 391
rect 1890 388 1902 391
rect 2026 391 2084 397
rect 2026 388 2038 391
rect 1890 360 2038 388
rect 1890 357 1902 360
rect 1839 351 1902 357
rect 2026 357 2038 360
rect 2072 357 2084 391
rect 2026 351 2084 357
rect 569 323 632 329
rect 569 289 586 323
rect 620 320 632 323
rect 942 323 1000 329
rect 942 320 954 323
rect 620 292 954 320
rect 620 289 632 292
rect 569 283 632 289
rect 942 289 954 292
rect 988 289 1000 323
rect 942 283 1000 289
rect 1678 323 1736 329
rect 1678 289 1690 323
rect 1724 320 1736 323
rect 2326 323 2384 329
rect 2326 320 2338 323
rect 1724 292 2338 320
rect 1724 289 1736 292
rect 1678 283 1736 289
rect 2326 289 2338 292
rect 2372 289 2384 323
rect 2326 283 2384 289
rect 385 255 443 261
rect 385 221 397 255
rect 431 252 443 255
rect 1218 255 1276 261
rect 1218 252 1230 255
rect 431 224 1230 252
rect 431 221 443 224
rect 385 215 443 221
rect 1218 221 1230 224
rect 1264 252 1276 255
rect 1770 255 1828 261
rect 1770 252 1782 255
rect 1264 224 1782 252
rect 1264 221 1276 224
rect 1218 215 1276 221
rect 1770 221 1782 224
rect 1816 221 1828 255
rect 1770 215 1828 221
rect 293 187 351 193
rect 293 153 305 187
rect 339 184 351 187
rect 850 187 908 193
rect 850 184 862 187
rect 339 156 862 184
rect 339 153 351 156
rect 293 147 351 153
rect 850 153 862 156
rect 896 153 908 187
rect 850 147 908 153
rect 1494 187 1552 193
rect 1494 153 1506 187
rect 1540 184 1552 187
rect 2234 187 2292 193
rect 2234 184 2246 187
rect 1540 156 2246 184
rect 1540 153 1552 156
rect 1494 147 1552 153
rect 2234 153 2246 156
rect 2280 153 2292 187
rect 2234 147 2292 153
rect 0 17 2484 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
rect 0 -48 2484 -17
<< labels >>
flabel locali s 1322 289 1356 323 0 FreeSans 300 0 0 0 COUT_N
port 8 nsew signal output
flabel locali s 305 153 339 187 0 FreeSans 300 0 0 0 B
port 2 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 300 180 0 0 A
port 1 nsew signal input
flabel locali s 2430 221 2464 255 0 FreeSans 300 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2150 221 2184 255 0 FreeSans 300 0 0 0 CI
port 3 nsew signal input
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 322 170 322 170 0 FreeSans 300 0 0 0 B
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 fahcon_1
rlabel viali s 862 153 896 187 1 B
port 2 nsew signal input
rlabel locali s 853 129 903 265 1 B
port 2 nsew signal input
rlabel metal1 s 850 184 908 193 1 B
port 2 nsew signal input
rlabel metal1 s 850 147 908 156 1 B
port 2 nsew signal input
rlabel metal1 s 293 184 351 193 1 B
port 2 nsew signal input
rlabel metal1 s 293 156 908 184 1 B
port 2 nsew signal input
rlabel metal1 s 293 147 351 156 1 B
port 2 nsew signal input
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2484 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 2192360
string GDS_START 2173556
string path 0.000 13.600 62.100 13.600 
<< end >>
