magic
tech sky130A
magscale 1 2
timestamp 1640697864
<< obsli1 >>
rect -32 2239 16032 42134
<< obsm1 >>
rect -29 824 16029 42193
<< metal2 >>
rect 297 0 353 480
rect 849 0 905 480
rect 1493 0 1549 480
rect 2137 0 2193 480
rect 2689 0 2745 480
rect 3333 0 3389 480
rect 3977 0 4033 480
rect 4529 0 4585 480
rect 5173 0 5229 480
rect 5817 0 5873 480
rect 6369 0 6425 480
rect 7013 0 7069 480
rect 7657 0 7713 480
rect 8301 0 8357 480
rect 8853 0 8909 480
rect 9497 0 9553 480
rect 10141 0 10197 480
rect 10693 0 10749 480
rect 11337 0 11393 480
rect 11981 0 12037 480
rect 12533 0 12589 480
rect 13177 0 13233 480
rect 13821 0 13877 480
rect 14373 0 14429 480
rect 15017 0 15073 480
rect 15661 0 15717 480
<< obsm2 >>
rect 42 536 15983 42193
rect 42 480 241 536
rect 409 480 793 536
rect 961 480 1437 536
rect 1605 480 2081 536
rect 2249 480 2633 536
rect 2801 480 3277 536
rect 3445 480 3921 536
rect 4089 480 4473 536
rect 4641 480 5117 536
rect 5285 480 5761 536
rect 5929 480 6313 536
rect 6481 480 6957 536
rect 7125 480 7601 536
rect 7769 480 8245 536
rect 8413 480 8797 536
rect 8965 480 9441 536
rect 9609 480 10085 536
rect 10253 480 10637 536
rect 10805 480 11281 536
rect 11449 480 11925 536
rect 12093 480 12477 536
rect 12645 480 13121 536
rect 13289 480 13765 536
rect 13933 480 14317 536
rect 14485 480 14961 536
rect 15129 480 15605 536
rect 15773 480 15983 536
<< obsm3 >>
rect 62 1931 15914 42193
<< metal4 >>
rect 0 37350 254 42193
rect 15746 37350 16000 42193
rect 0 16200 254 21193
rect 15746 16200 16000 21193
rect 0 15010 254 15900
rect 15746 15010 16000 15900
rect 0 13840 254 14730
rect 15746 13840 16000 14730
rect 0 13474 522 13540
rect 0 12818 7288 13414
rect 0 12522 254 12758
rect 9418 13474 16000 13540
rect 7752 12818 16000 13414
rect 0 11866 10429 12462
rect 15746 12522 16000 12758
rect 10893 11866 16000 12462
rect 0 11740 522 11806
rect 9418 11740 16000 11806
rect 0 10510 254 11440
rect 15746 10510 16000 11440
rect 0 9540 254 10230
rect 15746 9540 16000 10230
rect 0 8570 254 9260
rect 15746 8570 16000 9260
rect 0 7360 254 8290
rect 15746 7360 16000 8290
rect 0 6150 254 7080
rect 15746 6150 16000 7080
rect 0 5180 193 5870
rect 15794 5180 16000 5870
rect 0 3970 254 4900
rect 15746 3970 16000 4900
rect 0 2600 254 3690
rect 15746 2600 16000 3690
<< obsm4 >>
rect 334 37270 15666 42193
rect 193 21273 15794 37270
rect 334 16120 15666 21273
rect 193 15980 15794 16120
rect 334 14930 15666 15980
rect 193 14810 15794 14930
rect 334 13760 15666 14810
rect 193 13620 15794 13760
rect 602 13494 9338 13620
rect 7368 12738 7672 13494
rect 334 12542 15666 12738
rect 10509 11886 10813 12542
rect 602 11660 9338 11786
rect 193 11520 15794 11660
rect 334 10430 15666 11520
rect 193 10310 15794 10430
rect 334 9460 15666 10310
rect 193 9340 15794 9460
rect 334 8490 15666 9340
rect 193 8370 15794 8490
rect 334 7280 15666 8370
rect 193 7160 15794 7280
rect 334 6070 15666 7160
rect 193 5950 15794 6070
rect 273 5100 15714 5950
rect 193 4980 15794 5100
rect 334 3890 15666 4980
rect 193 3770 15794 3890
rect 334 2520 15666 3770
rect 193 2300 15794 2520
<< metal5 >>
rect 2240 23105 14760 35595
rect 0 16200 254 21190
rect 0 15030 254 15880
rect 0 13860 254 14710
rect 0 11740 254 13540
rect 0 10530 254 11420
rect 0 9561 254 10210
rect 0 8590 254 9240
rect 0 7380 254 8270
rect 0 6170 254 7060
rect 15746 16200 16000 21190
rect 15746 15030 16000 15880
rect 15746 13860 16000 14710
rect 15746 11740 16000 13540
rect 15746 10530 16000 11420
rect 15746 9561 16000 10210
rect 15746 8590 16000 9240
rect 15746 7380 16000 8270
rect 15746 6170 16000 7060
rect 0 5200 193 5850
rect 15794 5200 16000 5850
rect 0 3990 254 4880
rect 0 2620 254 3670
rect 15746 3990 16000 4880
rect 15746 2620 16000 3670
<< obsm5 >>
rect 0 35915 16000 42193
rect 0 22785 1920 35915
rect 15080 22785 16000 35915
rect 0 21510 16000 22785
rect 574 5850 15426 21510
rect 513 5200 15474 5850
rect 574 2620 15426 5200
<< labels >>
rlabel metal4 s 0 12818 7288 13414 6 AMUXBUS_A
port 28 nsew signal bidirectional
rlabel metal4 s 7752 12818 16000 13414 6 AMUXBUS_A
port 28 nsew signal bidirectional
rlabel metal4 s 0 11866 10429 12462 6 AMUXBUS_B
port 29 nsew signal bidirectional
rlabel metal4 s 10893 11866 16000 12462 6 AMUXBUS_B
port 29 nsew signal bidirectional
rlabel metal2 s 10141 0 10197 480 6 ANALOG_EN
port 22 nsew signal input
rlabel metal2 s 8853 0 8909 480 6 ANALOG_POL
port 26 nsew signal input
rlabel metal2 s 5817 0 5873 480 6 ANALOG_SEL
port 23 nsew signal input
rlabel metal2 s 5173 0 5229 480 6 DM[2]
port 6 nsew signal input
rlabel metal2 s 11337 0 11393 480 6 DM[1]
port 7 nsew signal input
rlabel metal2 s 9497 0 9553 480 6 DM[0]
port 8 nsew signal input
rlabel metal2 s 7013 0 7069 480 6 ENABLE_H
port 13 nsew signal input
rlabel metal2 s 7657 0 7713 480 6 ENABLE_INP_H
port 15 nsew signal input
rlabel metal2 s 2689 0 2745 480 6 ENABLE_VDDA_H
port 14 nsew signal input
rlabel metal2 s 13821 0 13877 480 6 ENABLE_VDDIO
port 24 nsew signal input
rlabel metal2 s 3333 0 3389 480 6 ENABLE_VSWITCH_H
port 25 nsew signal input
rlabel metal2 s 6369 0 6425 480 6 HLD_H_N
port 9 nsew signal input
rlabel metal2 s 4529 0 4585 480 6 HLD_OVR
port 21 nsew signal input
rlabel metal2 s 1493 0 1549 480 6 IB_MODE_SEL
port 12 nsew signal input
rlabel metal2 s 15017 0 15073 480 6 IN
port 10 nsew signal output
rlabel metal2 s 297 0 353 480 6 IN_H
port 1 nsew signal output
rlabel metal2 s 8301 0 8357 480 6 INP_DIS
port 11 nsew signal input
rlabel metal2 s 849 0 905 480 6 OE_N
port 16 nsew signal input
rlabel metal2 s 3977 0 4033 480 6 OUT
port 27 nsew signal input
rlabel metal5 s 2240 23105 14760 35595 6 PAD
port 5 nsew signal bidirectional
rlabel metal2 s 12533 0 12589 480 6 PAD_A_ESD_0_H
port 3 nsew signal bidirectional
rlabel metal2 s 11981 0 12037 480 6 PAD_A_ESD_1_H
port 4 nsew signal bidirectional
rlabel metal2 s 10693 0 10749 480 6 PAD_A_NOESD_H
port 2 nsew signal bidirectional
rlabel metal2 s 13177 0 13233 480 6 SLOW
port 19 nsew signal input
rlabel metal2 s 14373 0 14429 480 6 TIE_HI_ESD
port 17 nsew signal output
rlabel metal2 s 15661 0 15717 480 6 TIE_LO_ESD
port 18 nsew signal output
rlabel metal5 s 0 3990 254 4880 6 VCCD
port 36 nsew power bidirectional
rlabel metal4 s 0 3970 254 4900 6 VCCD
port 36 nsew power bidirectional
rlabel metal5 s 15746 3990 16000 4880 6 VCCD
port 36 nsew power bidirectional
rlabel metal4 s 15746 3970 16000 4900 6 VCCD
port 36 nsew power bidirectional
rlabel metal5 s 0 2620 254 3670 6 VCCHIB
port 34 nsew power bidirectional
rlabel metal4 s 0 2600 254 3690 6 VCCHIB
port 34 nsew power bidirectional
rlabel metal5 s 15746 2620 16000 3670 6 VCCHIB
port 34 nsew power bidirectional
rlabel metal4 s 15746 2600 16000 3690 6 VCCHIB
port 34 nsew power bidirectional
rlabel metal5 s 0 5200 193 5850 6 VDDA
port 31 nsew power bidirectional
rlabel metal4 s 0 5180 193 5870 6 VDDA
port 31 nsew power bidirectional
rlabel metal5 s 15794 5200 16000 5850 6 VDDA
port 31 nsew power bidirectional
rlabel metal4 s 15794 5180 16000 5870 6 VDDA
port 31 nsew power bidirectional
rlabel metal5 s 0 16200 254 21190 6 VDDIO
port 35 nsew power bidirectional
rlabel metal5 s 0 6170 254 7060 6 VDDIO
port 35 nsew power bidirectional
rlabel metal4 s 0 6150 254 7080 6 VDDIO
port 35 nsew power bidirectional
rlabel metal4 s 0 16200 254 21193 6 VDDIO
port 35 nsew power bidirectional
rlabel metal5 s 15746 16200 16000 21190 6 VDDIO
port 35 nsew power bidirectional
rlabel metal5 s 15746 6170 16000 7060 6 VDDIO
port 35 nsew power bidirectional
rlabel metal4 s 15746 6150 16000 7080 6 VDDIO
port 35 nsew power bidirectional
rlabel metal4 s 15746 16200 16000 21193 6 VDDIO
port 35 nsew power bidirectional
rlabel metal5 s 0 15030 254 15880 6 VDDIO_Q
port 33 nsew power bidirectional
rlabel metal4 s 0 15010 254 15900 6 VDDIO_Q
port 33 nsew power bidirectional
rlabel metal5 s 15746 15030 16000 15880 6 VDDIO_Q
port 33 nsew power bidirectional
rlabel metal4 s 15746 15010 16000 15900 6 VDDIO_Q
port 33 nsew power bidirectional
rlabel metal5 s 0 11740 254 13540 6 VSSA
port 30 nsew ground bidirectional
rlabel metal5 s 0 9561 254 10210 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 0 11740 522 11806 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 0 12522 254 12758 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 0 13474 522 13540 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 0 9540 254 10230 6 VSSA
port 30 nsew ground bidirectional
rlabel metal5 s 15746 11740 16000 13540 6 VSSA
port 30 nsew ground bidirectional
rlabel metal5 s 15746 9561 16000 10210 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 15746 12522 16000 12758 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 9418 13474 16000 13540 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 9418 11740 16000 11806 6 VSSA
port 30 nsew ground bidirectional
rlabel metal4 s 15746 9540 16000 10230 6 VSSA
port 30 nsew ground bidirectional
rlabel metal5 s 0 10530 254 11420 6 VSSD
port 38 nsew ground bidirectional
rlabel metal4 s 0 10510 254 11440 6 VSSD
port 38 nsew ground bidirectional
rlabel metal5 s 15746 10530 16000 11420 6 VSSD
port 38 nsew ground bidirectional
rlabel metal4 s 15746 10510 16000 11440 6 VSSD
port 38 nsew ground bidirectional
rlabel metal4 s 0 37350 254 42193 6 VSSIO
port 37 nsew ground bidirectional
rlabel metal5 s 0 7380 254 8270 6 VSSIO
port 37 nsew ground bidirectional
rlabel metal4 s 0 7360 254 8290 6 VSSIO
port 37 nsew ground bidirectional
rlabel metal4 s 15746 37350 16000 42193 6 VSSIO
port 37 nsew ground bidirectional
rlabel metal5 s 15746 7380 16000 8270 6 VSSIO
port 37 nsew ground bidirectional
rlabel metal4 s 15746 7360 16000 8290 6 VSSIO
port 37 nsew ground bidirectional
rlabel metal5 s 0 13860 254 14710 6 VSSIO_Q
port 39 nsew ground bidirectional
rlabel metal4 s 0 13840 254 14730 6 VSSIO_Q
port 39 nsew ground bidirectional
rlabel metal5 s 15746 13860 16000 14710 6 VSSIO_Q
port 39 nsew ground bidirectional
rlabel metal4 s 15746 13840 16000 14730 6 VSSIO_Q
port 39 nsew ground bidirectional
rlabel metal5 s 0 8590 254 9240 6 VSWITCH
port 32 nsew power bidirectional
rlabel metal4 s 0 8570 254 9260 6 VSWITCH
port 32 nsew power bidirectional
rlabel metal5 s 15746 8590 16000 9240 6 VSWITCH
port 32 nsew power bidirectional
rlabel metal4 s 15746 8570 16000 9260 6 VSWITCH
port 32 nsew power bidirectional
rlabel metal2 s 2137 0 2193 480 6 VTRIP_SEL
port 20 nsew signal input
<< properties >>
string LEFclass PAD INOUT
string FIXED_BBOX 0 0 16000 42193
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 8275438
string GDS_START 8250650
<< end >>
