magic
tech sky130A
magscale 1 2
timestamp 1619729575
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 275 333 341 425
rect 275 289 427 333
rect 18 215 162 255
rect 196 215 350 255
rect 384 181 427 289
rect 107 147 427 181
rect 107 145 341 147
rect 107 51 173 145
rect 275 51 341 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 18 333 73 493
rect 107 367 173 527
rect 207 459 435 493
rect 207 333 241 459
rect 18 291 241 333
rect 375 367 435 459
rect 18 17 73 181
rect 207 17 241 111
rect 375 17 433 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 18 215 162 255 6 A
port 1 nsew signal input
rlabel locali s 196 215 350 255 6 B
port 2 nsew signal input
rlabel locali s 384 181 427 289 6 Y
port 7 nsew signal output
rlabel locali s 275 333 341 425 6 Y
port 7 nsew signal output
rlabel locali s 275 289 427 333 6 Y
port 7 nsew signal output
rlabel locali s 275 51 341 145 6 Y
port 7 nsew signal output
rlabel locali s 107 147 427 181 6 Y
port 7 nsew signal output
rlabel locali s 107 145 341 147 6 Y
port 7 nsew signal output
rlabel locali s 107 51 173 145 6 Y
port 7 nsew signal output
rlabel metal1 s 0 -48 460 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3154814
string GDS_START 3150072
<< end >>
