magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1288 -1260 2888 1273
use sky130_fd_pr__hvdfm1sd__example_5595914180893  sky130_fd_pr__hvdfm1sd__example_5595914180893_0
timestamp 1619729480
transform 1 0 1600 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfm1sd__example_55959141808258  sky130_fd_pr__dfm1sd__example_55959141808258_0
timestamp 1619729480
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 1628 13 1628 13 0 FreeSans 300 0 0 0 D
flabel comment s -28 13 -28 13 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 37211922
string GDS_START 37210998
<< end >>
