magic
tech sky130A
timestamp 0
<< properties >>
string LEFclass CORE
string FIXED_BBOX 0 0 48 814
string LEFsymmetry y
string LEFview TRUE
<< end >>
