magic
tech sky130A
magscale 1 2
timestamp 1619729575
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 119 349 153 493
rect 287 349 321 493
rect 455 349 489 493
rect 623 349 657 493
rect 119 315 657 349
rect 119 161 163 315
rect 759 323 1207 333
rect 759 299 1134 323
rect 759 199 793 299
rect 1168 289 1207 323
rect 861 255 895 265
rect 892 221 895 255
rect 861 199 895 221
rect 119 127 657 161
rect 1036 163 1070 265
rect 1134 199 1207 289
rect 1405 233 1439 265
rect 1345 199 1439 233
rect 1592 255 1649 265
rect 1626 221 1649 255
rect 1592 199 1649 221
rect 1345 163 1379 199
rect 1036 129 1379 163
rect 119 51 153 127
rect 287 59 321 127
rect 455 51 489 127
rect 623 59 657 127
rect 1061 85 1178 129
rect 1843 289 1868 323
rect 1843 199 1902 289
<< viali >>
rect 1134 289 1168 323
rect 858 221 892 255
rect 1592 221 1626 255
rect 1868 289 1902 323
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 18 383 85 527
rect 187 383 253 527
rect 355 383 421 527
rect 523 383 589 527
rect 691 451 757 527
rect 791 451 1181 485
rect 1215 435 1249 527
rect 1296 451 1729 485
rect 1763 451 1829 527
rect 1863 417 1897 493
rect 691 367 1645 401
rect 1737 383 1897 417
rect 691 249 725 367
rect 1737 333 1771 383
rect 1863 359 1897 383
rect 197 215 725 249
rect 691 161 725 215
rect 950 161 984 187
rect 691 127 984 161
rect 1269 299 1771 333
rect 1269 199 1303 299
rect 1500 161 1534 187
rect 18 17 85 93
rect 187 17 253 93
rect 355 17 421 93
rect 523 17 589 93
rect 691 17 757 93
rect 791 59 1025 93
rect 1423 127 1534 161
rect 1737 163 1771 299
rect 1737 129 1897 163
rect 1212 17 1278 93
rect 1315 59 1573 93
rect 1763 17 1829 93
rect 1863 59 1897 129
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 1122 323 1180 329
rect 1122 289 1134 323
rect 1168 320 1180 323
rect 1856 323 1914 329
rect 1856 320 1868 323
rect 1168 292 1868 320
rect 1168 289 1180 292
rect 1122 283 1180 289
rect 1856 289 1868 292
rect 1902 289 1914 323
rect 1856 283 1914 289
rect 846 255 904 261
rect 846 221 858 255
rect 892 252 904 255
rect 1580 255 1638 261
rect 1580 252 1592 255
rect 892 224 1592 252
rect 892 221 904 224
rect 846 215 904 221
rect 1580 221 1592 224
rect 1626 221 1638 255
rect 1580 215 1638 221
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< obsm1 >>
rect 938 184 996 193
rect 1488 184 1546 193
rect 938 156 1546 184
rect 938 147 996 156
rect 1488 147 1546 156
<< labels >>
rlabel locali s 1405 233 1439 265 6 A0
port 1 nsew signal input
rlabel locali s 1345 199 1439 233 6 A0
port 1 nsew signal input
rlabel locali s 1345 163 1379 199 6 A0
port 1 nsew signal input
rlabel locali s 1061 85 1178 129 6 A0
port 1 nsew signal input
rlabel locali s 1036 163 1070 265 6 A0
port 1 nsew signal input
rlabel locali s 1036 129 1379 163 6 A0
port 1 nsew signal input
rlabel viali s 858 221 892 255 6 A1
port 2 nsew signal input
rlabel locali s 861 255 895 265 6 A1
port 2 nsew signal input
rlabel locali s 861 199 895 221 6 A1
port 2 nsew signal input
rlabel locali s 858 221 895 255 6 A1
port 2 nsew signal input
rlabel viali s 1592 221 1626 255 6 A1
port 2 nsew signal input
rlabel locali s 1592 199 1649 265 6 A1
port 2 nsew signal input
rlabel metal1 s 1580 252 1638 261 6 A1
port 2 nsew signal input
rlabel metal1 s 1580 215 1638 224 6 A1
port 2 nsew signal input
rlabel metal1 s 846 252 904 261 6 A1
port 2 nsew signal input
rlabel metal1 s 846 224 1638 252 6 A1
port 2 nsew signal input
rlabel metal1 s 846 215 904 224 6 A1
port 2 nsew signal input
rlabel viali s 1134 289 1168 323 6 S
port 3 nsew signal input
rlabel locali s 1134 199 1207 299 6 S
port 3 nsew signal input
rlabel locali s 759 299 1207 333 6 S
port 3 nsew signal input
rlabel locali s 759 199 793 299 6 S
port 3 nsew signal input
rlabel viali s 1868 289 1902 323 6 S
port 3 nsew signal input
rlabel locali s 1843 199 1902 323 6 S
port 3 nsew signal input
rlabel metal1 s 1856 320 1914 329 6 S
port 3 nsew signal input
rlabel metal1 s 1856 283 1914 292 6 S
port 3 nsew signal input
rlabel metal1 s 1122 320 1180 329 6 S
port 3 nsew signal input
rlabel metal1 s 1122 292 1914 320 6 S
port 3 nsew signal input
rlabel metal1 s 1122 283 1180 292 6 S
port 3 nsew signal input
rlabel locali s 623 349 657 493 6 X
port 8 nsew signal output
rlabel locali s 623 59 657 127 6 X
port 8 nsew signal output
rlabel locali s 455 349 489 493 6 X
port 8 nsew signal output
rlabel locali s 455 51 489 127 6 X
port 8 nsew signal output
rlabel locali s 287 349 321 493 6 X
port 8 nsew signal output
rlabel locali s 287 59 321 127 6 X
port 8 nsew signal output
rlabel locali s 119 349 153 493 6 X
port 8 nsew signal output
rlabel locali s 119 315 657 349 6 X
port 8 nsew signal output
rlabel locali s 119 161 163 315 6 X
port 8 nsew signal output
rlabel locali s 119 127 657 161 6 X
port 8 nsew signal output
rlabel locali s 119 51 153 127 6 X
port 8 nsew signal output
rlabel metal1 s 0 -48 1932 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1970 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1679350
string GDS_START 1666690
<< end >>
