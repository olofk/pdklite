magic
tech sky130A
magscale 1 2
timestamp 1640697977
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 643 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 164 47 194 177
rect 354 47 384 177
rect 440 47 470 177
rect 534 47 564 177
<< scpmoshvt >>
rect 79 297 109 497
rect 164 297 194 497
rect 354 297 384 497
rect 440 297 470 497
rect 534 297 564 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 101 164 177
rect 109 67 119 101
rect 153 67 164 101
rect 109 47 164 67
rect 194 93 247 177
rect 194 59 205 93
rect 239 59 247 93
rect 194 47 247 59
rect 301 162 354 177
rect 301 128 309 162
rect 343 128 354 162
rect 301 94 354 128
rect 301 60 309 94
rect 343 60 354 94
rect 301 47 354 60
rect 384 149 440 177
rect 384 115 395 149
rect 429 115 440 149
rect 384 47 440 115
rect 470 93 534 177
rect 470 59 485 93
rect 519 59 534 93
rect 470 47 534 59
rect 564 149 617 177
rect 564 115 575 149
rect 609 115 617 149
rect 564 47 617 115
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 380 79 451
rect 27 346 35 380
rect 69 346 79 380
rect 27 297 79 346
rect 109 477 164 497
rect 109 443 119 477
rect 153 443 164 477
rect 109 379 164 443
rect 109 345 119 379
rect 153 345 164 379
rect 109 297 164 345
rect 194 485 354 497
rect 194 451 205 485
rect 239 451 309 485
rect 343 451 354 485
rect 194 297 354 451
rect 384 477 440 497
rect 384 443 395 477
rect 429 443 440 477
rect 384 401 440 443
rect 384 367 395 401
rect 429 367 440 401
rect 384 297 440 367
rect 470 297 534 497
rect 564 485 617 497
rect 564 451 575 485
rect 609 451 617 485
rect 564 385 617 451
rect 564 351 575 385
rect 609 351 617 385
rect 564 297 617 351
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 67 153 101
rect 205 59 239 93
rect 309 128 343 162
rect 309 60 343 94
rect 395 115 429 149
rect 485 59 519 93
rect 575 115 609 149
<< pdiffc >>
rect 35 451 69 485
rect 35 346 69 380
rect 119 443 153 477
rect 119 345 153 379
rect 205 451 239 485
rect 309 451 343 485
rect 395 443 429 477
rect 395 367 429 401
rect 575 451 609 485
rect 575 351 609 385
<< poly >>
rect 79 497 109 523
rect 164 497 194 523
rect 354 497 384 523
rect 440 497 470 523
rect 534 497 564 523
rect 79 267 109 297
rect 164 267 194 297
rect 79 265 194 267
rect 354 265 384 297
rect 440 265 470 297
rect 534 265 564 297
rect 79 249 255 265
rect 79 215 205 249
rect 239 215 255 249
rect 79 199 255 215
rect 305 249 384 265
rect 305 215 321 249
rect 355 215 384 249
rect 305 199 384 215
rect 426 249 492 265
rect 426 215 442 249
rect 476 215 492 249
rect 426 199 492 215
rect 534 249 622 265
rect 534 215 578 249
rect 612 215 622 249
rect 534 199 622 215
rect 79 177 109 199
rect 164 177 194 199
rect 354 177 384 199
rect 440 177 470 199
rect 534 177 564 199
rect 79 21 109 47
rect 164 21 194 47
rect 354 21 384 47
rect 440 21 470 47
rect 534 21 564 47
<< polycont >>
rect 205 215 239 249
rect 321 215 355 249
rect 442 215 476 249
rect 578 215 612 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 380 69 451
rect 18 346 35 380
rect 18 327 69 346
rect 106 477 155 493
rect 106 443 119 477
rect 153 443 155 477
rect 106 379 155 443
rect 189 485 359 527
rect 189 451 205 485
rect 239 451 309 485
rect 343 451 359 485
rect 189 437 359 451
rect 393 477 445 493
rect 393 443 395 477
rect 429 443 445 477
rect 393 401 445 443
rect 106 345 119 379
rect 153 345 155 379
rect 21 161 69 177
rect 21 127 35 161
rect 21 93 69 127
rect 21 59 35 93
rect 21 17 69 59
rect 106 101 155 345
rect 221 367 395 401
rect 429 367 445 401
rect 559 485 624 527
rect 559 451 575 485
rect 609 451 624 485
rect 221 357 445 367
rect 221 266 255 357
rect 189 249 255 266
rect 189 215 205 249
rect 239 215 255 249
rect 189 168 255 215
rect 289 249 371 323
rect 481 280 522 397
rect 559 385 624 451
rect 559 351 575 385
rect 609 351 624 385
rect 559 330 624 351
rect 289 215 321 249
rect 355 215 371 249
rect 289 202 371 215
rect 405 249 522 280
rect 405 215 442 249
rect 476 215 522 249
rect 405 205 522 215
rect 573 249 625 290
rect 573 215 578 249
rect 612 215 625 249
rect 573 199 625 215
rect 189 162 359 168
rect 189 128 309 162
rect 343 128 359 162
rect 189 127 359 128
rect 106 67 119 101
rect 153 67 155 101
rect 293 94 359 127
rect 106 51 155 67
rect 189 59 205 93
rect 239 59 255 93
rect 189 17 255 59
rect 293 60 309 94
rect 343 60 359 94
rect 393 149 624 165
rect 393 115 395 149
rect 429 127 575 149
rect 429 115 435 127
rect 393 93 435 115
rect 569 115 575 127
rect 609 115 624 149
rect 569 99 624 115
rect 293 51 359 60
rect 469 59 485 93
rect 519 59 535 93
rect 469 17 535 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 580 221 614 255 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 304 289 338 323 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 488 357 522 391 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 120 425 154 459 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o21a_2
rlabel metal1 s 0 -48 644 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 1290992
string GDS_START 1285484
string path 0.000 0.000 3.220 0.000 
<< end >>
