magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1322 -1227 2260 3102
<< nwell >>
rect -37 1716 998 1824
rect -62 1500 998 1716
rect -62 1384 824 1500
<< pwell >>
rect 12 228 158 575
<< mvnmos >>
rect 112 1018 212 1102
rect 112 685 212 769
rect 286 228 386 1228
rect 442 228 542 1228
rect 598 228 698 1228
rect 754 228 854 1228
<< mvpmos >>
rect 57 1450 177 1650
rect 233 1450 353 1650
rect 409 1450 529 1650
rect 585 1450 705 1650
rect 779 1566 879 1650
<< mvndiff >>
rect 233 1158 286 1228
rect 233 1124 241 1158
rect 275 1124 286 1158
rect 233 1102 286 1124
rect 59 1090 112 1102
rect 59 1056 67 1090
rect 101 1056 112 1090
rect 59 1018 112 1056
rect 212 1090 286 1102
rect 212 1056 241 1090
rect 275 1056 286 1090
rect 212 1022 286 1056
rect 212 1018 241 1022
rect 233 988 241 1018
rect 275 988 286 1022
rect 233 954 286 988
rect 233 920 241 954
rect 275 920 286 954
rect 233 886 286 920
rect 233 852 241 886
rect 275 852 286 886
rect 233 818 286 852
rect 233 784 241 818
rect 275 784 286 818
rect 233 769 286 784
rect 59 731 112 769
rect 59 697 67 731
rect 101 697 112 731
rect 59 685 112 697
rect 212 750 286 769
rect 212 716 241 750
rect 275 716 286 750
rect 212 685 286 716
rect 233 682 286 685
rect 233 648 241 682
rect 275 648 286 682
rect 233 614 286 648
rect 233 580 241 614
rect 275 580 286 614
rect 233 546 286 580
rect 233 512 241 546
rect 275 512 286 546
rect 233 478 286 512
rect 233 444 241 478
rect 275 444 286 478
rect 233 410 286 444
rect 233 376 241 410
rect 275 376 286 410
rect 233 342 286 376
rect 233 308 241 342
rect 275 308 286 342
rect 233 274 286 308
rect 233 240 241 274
rect 275 240 286 274
rect 233 228 286 240
rect 386 1158 442 1228
rect 386 1124 397 1158
rect 431 1124 442 1158
rect 386 1090 442 1124
rect 386 1056 397 1090
rect 431 1056 442 1090
rect 386 1022 442 1056
rect 386 988 397 1022
rect 431 988 442 1022
rect 386 954 442 988
rect 386 920 397 954
rect 431 920 442 954
rect 386 886 442 920
rect 386 852 397 886
rect 431 852 442 886
rect 386 818 442 852
rect 386 784 397 818
rect 431 784 442 818
rect 386 750 442 784
rect 386 716 397 750
rect 431 716 442 750
rect 386 682 442 716
rect 386 648 397 682
rect 431 648 442 682
rect 386 614 442 648
rect 386 580 397 614
rect 431 580 442 614
rect 386 546 442 580
rect 386 512 397 546
rect 431 512 442 546
rect 386 478 442 512
rect 386 444 397 478
rect 431 444 442 478
rect 386 410 442 444
rect 386 376 397 410
rect 431 376 442 410
rect 386 342 442 376
rect 386 308 397 342
rect 431 308 442 342
rect 386 274 442 308
rect 386 240 397 274
rect 431 240 442 274
rect 386 228 442 240
rect 542 1158 598 1228
rect 542 1124 553 1158
rect 587 1124 598 1158
rect 542 1090 598 1124
rect 542 1056 553 1090
rect 587 1056 598 1090
rect 542 1022 598 1056
rect 542 988 553 1022
rect 587 988 598 1022
rect 542 954 598 988
rect 542 920 553 954
rect 587 920 598 954
rect 542 886 598 920
rect 542 852 553 886
rect 587 852 598 886
rect 542 818 598 852
rect 542 784 553 818
rect 587 784 598 818
rect 542 750 598 784
rect 542 716 553 750
rect 587 716 598 750
rect 542 682 598 716
rect 542 648 553 682
rect 587 648 598 682
rect 542 614 598 648
rect 542 580 553 614
rect 587 580 598 614
rect 542 546 598 580
rect 542 512 553 546
rect 587 512 598 546
rect 542 478 598 512
rect 542 444 553 478
rect 587 444 598 478
rect 542 410 598 444
rect 542 376 553 410
rect 587 376 598 410
rect 542 342 598 376
rect 542 308 553 342
rect 587 308 598 342
rect 542 274 598 308
rect 542 240 553 274
rect 587 240 598 274
rect 542 228 598 240
rect 698 1158 754 1228
rect 698 1124 709 1158
rect 743 1124 754 1158
rect 698 1090 754 1124
rect 698 1056 709 1090
rect 743 1056 754 1090
rect 698 1022 754 1056
rect 698 988 709 1022
rect 743 988 754 1022
rect 698 954 754 988
rect 698 920 709 954
rect 743 920 754 954
rect 698 886 754 920
rect 698 852 709 886
rect 743 852 754 886
rect 698 818 754 852
rect 698 784 709 818
rect 743 784 754 818
rect 698 750 754 784
rect 698 716 709 750
rect 743 716 754 750
rect 698 682 754 716
rect 698 648 709 682
rect 743 648 754 682
rect 698 614 754 648
rect 698 580 709 614
rect 743 580 754 614
rect 698 546 754 580
rect 698 512 709 546
rect 743 512 754 546
rect 698 478 754 512
rect 698 444 709 478
rect 743 444 754 478
rect 698 410 754 444
rect 698 376 709 410
rect 743 376 754 410
rect 698 342 754 376
rect 698 308 709 342
rect 743 308 754 342
rect 698 274 754 308
rect 698 240 709 274
rect 743 240 754 274
rect 698 228 754 240
rect 854 1158 907 1228
rect 854 1124 865 1158
rect 899 1124 907 1158
rect 854 1090 907 1124
rect 854 1056 865 1090
rect 899 1056 907 1090
rect 854 1022 907 1056
rect 854 988 865 1022
rect 899 988 907 1022
rect 854 954 907 988
rect 854 920 865 954
rect 899 920 907 954
rect 854 886 907 920
rect 854 852 865 886
rect 899 852 907 886
rect 854 818 907 852
rect 854 784 865 818
rect 899 784 907 818
rect 854 750 907 784
rect 854 716 865 750
rect 899 716 907 750
rect 854 682 907 716
rect 854 648 865 682
rect 899 648 907 682
rect 854 614 907 648
rect 854 580 865 614
rect 899 580 907 614
rect 854 546 907 580
rect 854 512 865 546
rect 899 512 907 546
rect 854 478 907 512
rect 854 444 865 478
rect 899 444 907 478
rect 854 410 907 444
rect 854 376 865 410
rect 899 376 907 410
rect 854 342 907 376
rect 854 308 865 342
rect 899 308 907 342
rect 854 274 907 308
rect 854 240 865 274
rect 899 240 907 274
rect 854 228 907 240
<< mvpdiff >>
rect 4 1638 57 1650
rect 4 1604 12 1638
rect 46 1604 57 1638
rect 4 1570 57 1604
rect 4 1536 12 1570
rect 46 1536 57 1570
rect 4 1502 57 1536
rect 4 1468 12 1502
rect 46 1468 57 1502
rect 4 1450 57 1468
rect 177 1638 233 1650
rect 177 1604 188 1638
rect 222 1604 233 1638
rect 177 1570 233 1604
rect 177 1536 188 1570
rect 222 1536 233 1570
rect 177 1502 233 1536
rect 177 1468 188 1502
rect 222 1468 233 1502
rect 177 1450 233 1468
rect 353 1638 409 1650
rect 353 1604 364 1638
rect 398 1604 409 1638
rect 353 1570 409 1604
rect 353 1536 364 1570
rect 398 1536 409 1570
rect 353 1502 409 1536
rect 353 1468 364 1502
rect 398 1468 409 1502
rect 353 1450 409 1468
rect 529 1638 585 1650
rect 529 1604 540 1638
rect 574 1604 585 1638
rect 529 1570 585 1604
rect 529 1536 540 1570
rect 574 1536 585 1570
rect 529 1502 585 1536
rect 529 1468 540 1502
rect 574 1468 585 1502
rect 529 1450 585 1468
rect 705 1638 779 1650
rect 705 1604 716 1638
rect 750 1604 779 1638
rect 705 1570 779 1604
rect 705 1536 716 1570
rect 750 1566 779 1570
rect 879 1638 932 1650
rect 879 1604 890 1638
rect 924 1604 932 1638
rect 879 1566 932 1604
rect 750 1536 758 1566
rect 705 1502 758 1536
rect 705 1468 716 1502
rect 750 1468 758 1502
rect 705 1450 758 1468
<< mvndiffc >>
rect 241 1124 275 1158
rect 67 1056 101 1090
rect 241 1056 275 1090
rect 241 988 275 1022
rect 241 920 275 954
rect 241 852 275 886
rect 241 784 275 818
rect 67 697 101 731
rect 241 716 275 750
rect 241 648 275 682
rect 241 580 275 614
rect 241 512 275 546
rect 241 444 275 478
rect 241 376 275 410
rect 241 308 275 342
rect 241 240 275 274
rect 397 1124 431 1158
rect 397 1056 431 1090
rect 397 988 431 1022
rect 397 920 431 954
rect 397 852 431 886
rect 397 784 431 818
rect 397 716 431 750
rect 397 648 431 682
rect 397 580 431 614
rect 397 512 431 546
rect 397 444 431 478
rect 397 376 431 410
rect 397 308 431 342
rect 397 240 431 274
rect 553 1124 587 1158
rect 553 1056 587 1090
rect 553 988 587 1022
rect 553 920 587 954
rect 553 852 587 886
rect 553 784 587 818
rect 553 716 587 750
rect 553 648 587 682
rect 553 580 587 614
rect 553 512 587 546
rect 553 444 587 478
rect 553 376 587 410
rect 553 308 587 342
rect 553 240 587 274
rect 709 1124 743 1158
rect 709 1056 743 1090
rect 709 988 743 1022
rect 709 920 743 954
rect 709 852 743 886
rect 709 784 743 818
rect 709 716 743 750
rect 709 648 743 682
rect 709 580 743 614
rect 709 512 743 546
rect 709 444 743 478
rect 709 376 743 410
rect 709 308 743 342
rect 709 240 743 274
rect 865 1124 899 1158
rect 865 1056 899 1090
rect 865 988 899 1022
rect 865 920 899 954
rect 865 852 899 886
rect 865 784 899 818
rect 865 716 899 750
rect 865 648 899 682
rect 865 580 899 614
rect 865 512 899 546
rect 865 444 899 478
rect 865 376 899 410
rect 865 308 899 342
rect 865 240 899 274
<< mvpdiffc >>
rect 12 1604 46 1638
rect 12 1536 46 1570
rect 12 1468 46 1502
rect 188 1604 222 1638
rect 188 1536 222 1570
rect 188 1468 222 1502
rect 364 1604 398 1638
rect 364 1536 398 1570
rect 364 1468 398 1502
rect 540 1604 574 1638
rect 540 1536 574 1570
rect 540 1468 574 1502
rect 716 1604 750 1638
rect 716 1536 750 1570
rect 890 1604 924 1638
rect 716 1468 750 1502
<< psubdiff >>
rect 12 551 158 575
rect 46 517 124 551
rect 12 462 158 517
rect 46 428 124 462
rect 12 374 158 428
rect 46 340 124 374
rect 12 286 158 340
rect 46 252 124 286
rect 12 228 158 252
<< mvnsubdiff >>
rect 29 1724 63 1758
rect 97 1724 135 1758
rect 169 1724 207 1758
rect 241 1724 280 1758
rect 314 1724 353 1758
rect 387 1724 426 1758
rect 460 1724 499 1758
rect 533 1724 572 1758
rect 606 1724 645 1758
rect 679 1724 718 1758
rect 752 1724 791 1758
rect 825 1724 864 1758
rect 898 1724 932 1758
<< psubdiffcont >>
rect 12 517 46 551
rect 124 517 158 551
rect 12 428 46 462
rect 124 428 158 462
rect 12 340 46 374
rect 124 340 158 374
rect 12 252 46 286
rect 124 252 158 286
<< mvnsubdiffcont >>
rect 63 1724 97 1758
rect 135 1724 169 1758
rect 207 1724 241 1758
rect 280 1724 314 1758
rect 353 1724 387 1758
rect 426 1724 460 1758
rect 499 1724 533 1758
rect 572 1724 606 1758
rect 645 1724 679 1758
rect 718 1724 752 1758
rect 791 1724 825 1758
rect 864 1724 898 1758
<< poly >>
rect 57 1650 177 1682
rect 233 1650 353 1682
rect 409 1650 529 1682
rect 585 1650 705 1682
rect 779 1650 879 1682
rect 779 1517 879 1566
rect 779 1483 821 1517
rect 855 1483 879 1517
rect 57 1418 177 1450
rect 233 1418 353 1450
rect 57 1402 353 1418
rect 57 1368 73 1402
rect 107 1368 150 1402
rect 184 1368 227 1402
rect 261 1368 303 1402
rect 337 1368 353 1402
rect 57 1352 353 1368
rect 409 1418 529 1450
rect 585 1418 705 1450
rect 409 1402 705 1418
rect 409 1368 425 1402
rect 459 1368 501 1402
rect 535 1368 578 1402
rect 612 1368 655 1402
rect 689 1368 705 1402
rect 779 1449 879 1483
rect 779 1415 821 1449
rect 855 1415 879 1449
rect 779 1399 879 1415
rect 409 1352 705 1368
rect 112 1271 212 1288
rect 112 1237 145 1271
rect 179 1237 212 1271
rect 112 1203 212 1237
rect 286 1228 386 1260
rect 442 1228 542 1260
rect 598 1228 698 1260
rect 754 1228 854 1260
rect 112 1169 145 1203
rect 179 1169 212 1203
rect 112 1102 212 1169
rect 112 986 212 1018
rect 112 919 212 935
rect 112 885 145 919
rect 179 885 212 919
rect 112 851 212 885
rect 112 817 145 851
rect 179 817 212 851
rect 112 769 212 817
rect 112 653 212 685
rect 286 158 386 228
rect 286 124 319 158
rect 353 124 386 158
rect 286 90 386 124
rect 286 56 319 90
rect 353 56 386 90
rect 286 40 386 56
rect 442 158 542 228
rect 442 124 479 158
rect 513 124 542 158
rect 442 90 542 124
rect 442 56 479 90
rect 513 56 542 90
rect 442 40 542 56
rect 598 158 698 228
rect 598 124 629 158
rect 663 124 698 158
rect 598 90 698 124
rect 598 56 629 90
rect 663 56 698 90
rect 598 40 698 56
rect 754 156 854 228
rect 754 122 784 156
rect 818 122 854 156
rect 754 88 854 122
rect 754 54 784 88
rect 818 54 854 88
rect 754 38 854 54
<< polycont >>
rect 821 1483 855 1517
rect 73 1368 107 1402
rect 150 1368 184 1402
rect 227 1368 261 1402
rect 303 1368 337 1402
rect 425 1368 459 1402
rect 501 1368 535 1402
rect 578 1368 612 1402
rect 655 1368 689 1402
rect 821 1415 855 1449
rect 145 1237 179 1271
rect 145 1169 179 1203
rect 145 885 179 919
rect 145 817 179 851
rect 319 124 353 158
rect 319 56 353 90
rect 479 124 513 158
rect 479 56 513 90
rect 629 124 663 158
rect 629 56 663 90
rect 784 122 818 156
rect 784 54 818 88
<< locali >>
rect 29 1724 63 1758
rect 127 1724 135 1758
rect 200 1724 207 1758
rect 273 1724 280 1758
rect 347 1724 353 1758
rect 421 1724 426 1758
rect 460 1724 461 1758
rect 495 1724 499 1758
rect 533 1724 535 1758
rect 569 1724 572 1758
rect 606 1724 609 1758
rect 643 1724 645 1758
rect 679 1724 683 1758
rect 717 1724 718 1758
rect 752 1724 757 1758
rect 825 1724 831 1758
rect 898 1724 932 1758
rect 12 1582 46 1604
rect 12 1510 46 1536
rect 12 1452 46 1468
rect 188 1582 222 1604
rect 188 1510 222 1536
rect 188 1452 222 1468
rect 364 1582 398 1604
rect 364 1510 398 1536
rect 364 1452 398 1468
rect 540 1582 574 1604
rect 540 1510 574 1536
rect 540 1452 574 1468
rect 716 1582 750 1604
rect 890 1582 924 1604
rect 716 1510 750 1536
rect 716 1452 750 1468
rect 801 1522 816 1556
rect 850 1522 856 1556
rect 801 1517 856 1522
rect 801 1484 821 1517
rect 855 1514 856 1517
rect 801 1450 816 1484
rect 855 1483 939 1514
rect 850 1450 939 1483
rect 801 1449 939 1450
rect 801 1415 821 1449
rect 855 1415 939 1449
rect 57 1368 73 1402
rect 107 1368 150 1402
rect 184 1368 227 1402
rect 261 1368 303 1402
rect 337 1368 363 1402
rect 409 1368 425 1402
rect 459 1368 501 1402
rect 535 1368 578 1402
rect 612 1368 655 1402
rect 689 1400 705 1402
rect 689 1368 722 1400
rect 153 1299 191 1333
rect 119 1271 225 1299
rect 119 1237 145 1271
rect 179 1237 225 1271
rect 119 1205 225 1237
rect 119 1203 203 1205
rect 119 1169 145 1203
rect 179 1169 203 1203
rect 309 1181 363 1368
rect 424 1356 722 1368
rect 424 1322 478 1356
rect 512 1322 568 1356
rect 602 1322 658 1356
rect 692 1322 722 1356
rect 424 1316 722 1322
rect 801 1282 939 1415
rect 732 1248 770 1282
rect 804 1248 939 1282
rect 698 1229 939 1248
rect 119 1153 203 1169
rect 67 1034 101 1056
rect 137 1093 203 1153
rect 137 1059 143 1093
rect 177 1059 203 1093
rect 137 1021 203 1059
rect 137 987 143 1021
rect 177 987 203 1021
rect 137 986 203 987
rect 241 1158 275 1174
rect 241 1092 275 1124
rect 309 1147 320 1181
rect 354 1147 363 1181
rect 309 1109 363 1147
rect 309 1075 320 1109
rect 354 1075 363 1109
rect 309 1074 363 1075
rect 397 1158 431 1160
rect 397 1122 431 1124
rect 241 1022 275 1056
rect 241 954 275 983
rect 101 919 179 935
rect 101 901 145 919
rect 67 885 145 901
rect 67 863 179 885
rect 101 851 179 863
rect 101 829 145 851
rect 67 817 145 829
rect 67 801 179 817
rect 241 886 275 908
rect 241 818 275 832
rect 241 750 275 756
rect 67 731 101 747
rect 67 643 101 681
rect 241 714 275 716
rect 241 638 275 648
rect 12 557 158 575
rect 46 523 116 557
rect 150 551 158 557
rect 46 517 124 523
rect 12 483 158 517
rect 46 449 116 483
rect 150 462 158 483
rect 46 428 124 449
rect 12 409 158 428
rect 46 375 116 409
rect 150 375 158 409
rect 12 374 158 375
rect 46 340 124 374
rect 12 335 158 340
rect 46 301 116 335
rect 150 301 158 335
rect 12 286 158 301
rect 46 262 124 286
rect 46 228 116 262
rect 150 228 158 252
rect 241 562 275 580
rect 241 486 275 512
rect 241 410 275 444
rect 241 342 275 376
rect 241 274 275 300
rect 397 1050 431 1056
rect 397 978 431 988
rect 397 906 431 920
rect 397 834 431 852
rect 397 762 431 784
rect 397 690 431 716
rect 397 618 431 648
rect 397 546 431 580
rect 397 478 431 512
rect 397 410 431 440
rect 397 342 431 368
rect 397 274 431 296
rect 553 1158 587 1160
rect 553 1122 587 1124
rect 553 1050 587 1056
rect 553 978 587 988
rect 553 906 587 920
rect 553 834 587 852
rect 553 762 587 784
rect 553 690 587 716
rect 553 618 587 648
rect 553 546 587 580
rect 553 478 587 512
rect 553 410 587 440
rect 553 342 587 368
rect 553 274 587 296
rect 709 1158 743 1160
rect 709 1122 743 1124
rect 709 1050 743 1056
rect 709 978 743 988
rect 709 906 743 920
rect 709 834 743 852
rect 709 762 743 784
rect 709 690 743 716
rect 709 618 743 648
rect 709 546 743 580
rect 709 478 743 512
rect 709 410 743 440
rect 709 342 743 368
rect 709 274 743 296
rect 865 1158 899 1160
rect 865 1122 899 1124
rect 865 1050 899 1056
rect 865 978 899 988
rect 865 906 899 920
rect 865 834 899 852
rect 865 762 899 784
rect 865 690 899 716
rect 865 618 899 648
rect 865 546 899 580
rect 865 478 899 512
rect 865 410 899 440
rect 865 342 899 368
rect 865 274 899 296
rect 319 158 320 174
rect 353 124 354 147
rect 319 109 354 124
rect 319 90 320 109
rect 479 158 513 174
rect 479 90 513 124
rect 319 40 353 56
rect 479 40 513 56
rect 629 158 663 174
rect 629 90 663 124
rect 629 40 663 56
rect 784 156 818 172
rect 784 88 818 122
rect 784 38 818 54
<< viali >>
rect 93 1724 97 1758
rect 97 1724 127 1758
rect 166 1724 169 1758
rect 169 1724 200 1758
rect 239 1724 241 1758
rect 241 1724 273 1758
rect 313 1724 314 1758
rect 314 1724 347 1758
rect 387 1724 421 1758
rect 461 1724 495 1758
rect 535 1724 569 1758
rect 609 1724 643 1758
rect 683 1724 717 1758
rect 757 1724 791 1758
rect 831 1724 864 1758
rect 864 1724 865 1758
rect 12 1638 46 1654
rect 12 1620 46 1638
rect 12 1570 46 1582
rect 12 1548 46 1570
rect 12 1502 46 1510
rect 12 1476 46 1502
rect 188 1638 222 1654
rect 188 1620 222 1638
rect 188 1570 222 1582
rect 188 1548 222 1570
rect 188 1502 222 1510
rect 188 1476 222 1502
rect 364 1638 398 1654
rect 364 1620 398 1638
rect 364 1570 398 1582
rect 364 1548 398 1570
rect 364 1502 398 1510
rect 364 1476 398 1502
rect 540 1638 574 1654
rect 540 1620 574 1638
rect 540 1570 574 1582
rect 540 1548 574 1570
rect 540 1502 574 1510
rect 540 1476 574 1502
rect 716 1638 750 1654
rect 716 1620 750 1638
rect 716 1570 750 1582
rect 716 1548 750 1570
rect 890 1638 924 1654
rect 890 1620 924 1638
rect 716 1502 750 1510
rect 716 1476 750 1502
rect 816 1522 850 1556
rect 890 1548 924 1582
rect 816 1483 821 1484
rect 821 1483 850 1484
rect 816 1450 850 1483
rect 119 1299 153 1333
rect 191 1299 225 1333
rect 478 1322 512 1356
rect 568 1322 602 1356
rect 658 1322 692 1356
rect 698 1248 732 1282
rect 770 1248 804 1282
rect 67 1090 101 1106
rect 67 1072 101 1090
rect 67 1000 101 1034
rect 143 1059 177 1093
rect 143 987 177 1021
rect 241 1090 275 1092
rect 241 1058 275 1090
rect 320 1147 354 1181
rect 320 1075 354 1109
rect 397 1160 431 1194
rect 397 1090 431 1122
rect 397 1088 431 1090
rect 241 988 275 1017
rect 241 983 275 988
rect 67 901 101 935
rect 67 829 101 863
rect 241 920 275 942
rect 241 908 275 920
rect 241 852 275 866
rect 241 832 275 852
rect 241 784 275 790
rect 241 756 275 784
rect 67 697 101 715
rect 67 681 101 697
rect 67 609 101 643
rect 241 682 275 714
rect 241 680 275 682
rect 241 614 275 638
rect 241 604 275 614
rect 12 551 46 557
rect 12 523 46 551
rect 116 551 150 557
rect 116 523 124 551
rect 124 523 150 551
rect 12 462 46 483
rect 12 449 46 462
rect 116 462 150 483
rect 116 449 124 462
rect 124 449 150 462
rect 12 375 46 409
rect 116 375 150 409
rect 12 301 46 335
rect 116 301 150 335
rect 12 252 46 262
rect 12 228 46 252
rect 116 252 124 262
rect 124 252 150 262
rect 116 228 150 252
rect 241 546 275 562
rect 241 528 275 546
rect 241 478 275 486
rect 241 452 275 478
rect 241 376 275 410
rect 241 308 275 334
rect 241 300 275 308
rect 241 240 275 258
rect 241 224 275 240
rect 397 1022 431 1050
rect 397 1016 431 1022
rect 397 954 431 978
rect 397 944 431 954
rect 397 886 431 906
rect 397 872 431 886
rect 397 818 431 834
rect 397 800 431 818
rect 397 750 431 762
rect 397 728 431 750
rect 397 682 431 690
rect 397 656 431 682
rect 397 614 431 618
rect 397 584 431 614
rect 397 512 431 546
rect 397 444 431 474
rect 397 440 431 444
rect 397 376 431 402
rect 397 368 431 376
rect 397 308 431 330
rect 397 296 431 308
rect 397 240 431 258
rect 397 224 431 240
rect 553 1160 587 1194
rect 553 1090 587 1122
rect 553 1088 587 1090
rect 553 1022 587 1050
rect 553 1016 587 1022
rect 553 954 587 978
rect 553 944 587 954
rect 553 886 587 906
rect 553 872 587 886
rect 553 818 587 834
rect 553 800 587 818
rect 553 750 587 762
rect 553 728 587 750
rect 553 682 587 690
rect 553 656 587 682
rect 553 614 587 618
rect 553 584 587 614
rect 553 512 587 546
rect 553 444 587 474
rect 553 440 587 444
rect 553 376 587 402
rect 553 368 587 376
rect 553 308 587 330
rect 553 296 587 308
rect 553 240 587 258
rect 553 224 587 240
rect 709 1160 743 1194
rect 709 1090 743 1122
rect 709 1088 743 1090
rect 709 1022 743 1050
rect 709 1016 743 1022
rect 709 954 743 978
rect 709 944 743 954
rect 709 886 743 906
rect 709 872 743 886
rect 709 818 743 834
rect 709 800 743 818
rect 709 750 743 762
rect 709 728 743 750
rect 709 682 743 690
rect 709 656 743 682
rect 709 614 743 618
rect 709 584 743 614
rect 709 512 743 546
rect 709 444 743 474
rect 709 440 743 444
rect 709 376 743 402
rect 709 368 743 376
rect 709 308 743 330
rect 709 296 743 308
rect 709 240 743 258
rect 709 224 743 240
rect 865 1160 899 1194
rect 865 1090 899 1122
rect 865 1088 899 1090
rect 865 1022 899 1050
rect 865 1016 899 1022
rect 865 954 899 978
rect 865 944 899 954
rect 865 886 899 906
rect 865 872 899 886
rect 865 818 899 834
rect 865 800 899 818
rect 865 750 899 762
rect 865 728 899 750
rect 865 682 899 690
rect 865 656 899 682
rect 865 614 899 618
rect 865 584 899 614
rect 865 512 899 546
rect 865 444 899 474
rect 865 440 899 444
rect 865 376 899 402
rect 865 368 899 376
rect 865 308 899 330
rect 865 296 899 308
rect 865 240 899 258
rect 865 224 899 240
rect 320 158 354 181
rect 320 147 353 158
rect 353 147 354 158
rect 320 90 354 109
rect 320 75 353 90
rect 353 75 354 90
<< metal1 >>
rect 6 1758 1000 1842
rect 6 1724 93 1758
rect 127 1724 166 1758
rect 200 1724 239 1758
rect 273 1724 313 1758
rect 347 1724 387 1758
rect 421 1724 461 1758
rect 495 1724 535 1758
rect 569 1724 609 1758
rect 643 1724 683 1758
rect 717 1724 757 1758
rect 791 1724 831 1758
rect 865 1724 1000 1758
rect 6 1714 1000 1724
rect 6 1654 52 1714
tri 52 1680 86 1714 nw
tri 324 1680 358 1714 ne
rect 358 1684 408 1714
tri 408 1684 438 1714 nw
tri 680 1684 710 1714 ne
rect 6 1620 12 1654
rect 46 1620 52 1654
rect 6 1582 52 1620
rect 6 1548 12 1582
rect 46 1548 52 1582
rect 6 1510 52 1548
rect 6 1476 12 1510
rect 46 1476 52 1510
rect 6 1464 52 1476
rect 182 1654 228 1666
rect 182 1620 188 1654
rect 222 1620 228 1654
rect 182 1582 228 1620
rect 182 1548 188 1582
rect 222 1548 228 1582
rect 182 1510 228 1548
rect 358 1654 404 1684
tri 404 1680 408 1684 nw
rect 358 1620 364 1654
rect 398 1620 404 1654
rect 358 1582 404 1620
rect 358 1548 364 1582
rect 398 1548 404 1582
tri 228 1510 234 1516 sw
rect 358 1510 404 1548
rect 182 1476 188 1510
rect 222 1476 234 1510
tri 234 1476 268 1510 sw
rect 358 1476 364 1510
rect 398 1476 404 1510
rect 182 1475 268 1476
tri 268 1475 269 1476 sw
rect 182 1464 269 1475
tri 269 1464 280 1475 sw
rect 358 1464 404 1476
rect 534 1654 580 1666
rect 534 1620 540 1654
rect 574 1620 580 1654
rect 534 1582 580 1620
rect 534 1548 540 1582
rect 574 1548 580 1582
rect 534 1510 580 1548
rect 534 1476 540 1510
rect 574 1476 580 1510
rect 534 1474 580 1476
rect 710 1654 756 1714
tri 756 1684 786 1714 nw
rect 710 1620 716 1654
rect 750 1620 756 1654
rect 710 1582 756 1620
rect 710 1548 716 1582
rect 750 1548 756 1582
rect 884 1654 930 1666
rect 884 1620 890 1654
rect 924 1620 930 1654
rect 884 1582 930 1620
rect 710 1510 756 1548
rect 710 1476 716 1510
rect 750 1476 756 1510
tri 580 1474 581 1475 sw
rect 182 1450 280 1464
tri 280 1450 294 1464 sw
rect 534 1450 581 1474
tri 581 1450 605 1474 sw
rect 710 1464 756 1476
rect 810 1556 856 1568
rect 810 1522 816 1556
rect 850 1522 856 1556
rect 810 1484 856 1522
tri 800 1464 810 1474 se
rect 810 1464 816 1484
tri 786 1450 800 1464 se
rect 800 1450 816 1464
rect 850 1450 856 1484
tri 122 1362 182 1422 se
rect 182 1391 294 1450
tri 294 1391 353 1450 sw
rect 534 1438 605 1450
tri 605 1438 617 1450 sw
tri 774 1438 786 1450 se
rect 786 1438 856 1450
rect 534 1436 617 1438
tri 617 1436 619 1438 sw
tri 772 1436 774 1438 se
rect 774 1436 843 1438
rect 534 1425 843 1436
tri 843 1425 856 1438 nw
rect 884 1548 890 1582
rect 924 1548 930 1582
tri 534 1391 568 1425 ne
rect 568 1391 809 1425
tri 809 1391 843 1425 nw
tri 875 1391 884 1400 se
rect 884 1391 930 1548
rect 182 1362 353 1391
tri 353 1362 382 1391 sw
tri 846 1362 875 1391 se
rect 875 1365 930 1391
rect 875 1362 927 1365
tri 927 1362 930 1365 nw
rect 107 1356 905 1362
rect 107 1333 478 1356
rect 107 1299 119 1333
rect 153 1299 191 1333
rect 225 1322 478 1333
rect 512 1322 568 1356
rect 602 1322 658 1356
rect 692 1322 905 1356
tri 905 1340 927 1362 nw
rect 225 1316 905 1322
rect 225 1299 237 1316
rect 107 1293 237 1299
tri 237 1293 260 1316 nw
tri 834 1293 857 1316 ne
rect 857 1293 905 1316
tri 857 1291 859 1293 ne
tri 272 1282 278 1288 se
rect 278 1282 816 1288
tri 238 1248 272 1282 se
rect 272 1248 698 1282
rect 732 1248 770 1282
rect 804 1248 816 1282
tri 221 1231 238 1248 se
rect 238 1242 816 1248
rect 238 1231 287 1242
tri 287 1231 298 1242 nw
tri 81 1194 118 1231 se
rect 118 1194 250 1231
tri 250 1194 287 1231 nw
rect 391 1194 437 1206
tri 80 1193 81 1194 se
rect 81 1193 249 1194
tri 249 1193 250 1194 nw
tri 68 1181 80 1193 se
rect 80 1185 241 1193
tri 241 1185 249 1193 nw
rect 80 1181 134 1185
tri 134 1181 138 1185 nw
rect 309 1181 363 1193
tri 61 1174 68 1181 se
rect 68 1174 127 1181
tri 127 1174 134 1181 nw
rect 61 1106 107 1174
tri 107 1154 127 1174 nw
rect 61 1072 67 1106
rect 101 1072 107 1106
rect 309 1147 320 1181
rect 354 1147 363 1181
rect 309 1109 363 1147
rect 61 1034 107 1072
rect 61 1000 67 1034
rect 101 1000 107 1034
rect 61 935 107 1000
rect 137 1093 183 1105
rect 137 1059 143 1093
rect 177 1059 183 1093
rect 137 1021 183 1059
rect 137 987 143 1021
rect 177 987 183 1021
rect 137 975 183 987
rect 235 1092 281 1104
rect 235 1058 241 1092
rect 275 1058 281 1092
rect 235 1017 281 1058
rect 235 983 241 1017
rect 275 983 281 1017
rect 61 901 67 935
rect 101 901 107 935
rect 61 863 107 901
rect 61 829 67 863
rect 101 829 107 863
rect 61 817 107 829
rect 235 942 281 983
rect 235 908 241 942
rect 275 908 281 942
rect 235 866 281 908
rect 235 832 241 866
rect 275 832 281 866
rect 235 790 281 832
tri 223 756 235 768 se
rect 235 756 241 790
rect 275 756 281 790
tri 195 728 223 756 se
rect 223 728 281 756
tri 194 727 195 728 se
rect 195 727 281 728
rect 29 715 281 727
rect 29 681 67 715
rect 101 714 281 715
rect 101 681 241 714
rect 29 680 241 681
rect 275 680 281 714
rect 29 643 281 680
rect 29 609 67 643
rect 101 638 281 643
rect 101 609 241 638
rect 29 604 241 609
rect 275 604 281 638
rect 29 569 281 604
rect 6 562 281 569
rect 6 557 241 562
rect 6 523 12 557
rect 46 523 116 557
rect 150 528 241 557
rect 275 528 281 562
rect 150 523 281 528
rect 6 486 281 523
rect 6 483 241 486
rect 6 449 12 483
rect 46 449 116 483
rect 150 452 241 483
rect 275 452 281 486
rect 150 449 281 452
rect 6 410 281 449
rect 6 409 241 410
rect 6 375 12 409
rect 46 375 116 409
rect 150 376 241 409
rect 275 376 281 410
rect 150 375 281 376
rect 6 335 281 375
rect 6 301 12 335
rect 46 301 116 335
rect 150 334 281 335
rect 150 301 241 334
rect 6 300 241 301
rect 275 300 281 334
rect 6 262 281 300
rect 6 228 12 262
rect 46 228 116 262
rect 150 258 281 262
rect 150 228 241 258
rect 6 224 241 228
rect 275 224 281 258
rect 6 216 281 224
rect 29 212 281 216
rect 309 1075 320 1109
rect 354 1075 363 1109
rect 309 181 363 1075
rect 391 1160 397 1194
rect 431 1160 437 1194
rect 391 1122 437 1160
rect 391 1088 397 1122
rect 431 1088 437 1122
rect 391 1050 437 1088
rect 391 1016 397 1050
rect 431 1016 437 1050
rect 391 978 437 1016
rect 391 944 397 978
rect 431 944 437 978
rect 391 906 437 944
rect 391 872 397 906
rect 431 872 437 906
rect 391 834 437 872
rect 391 800 397 834
rect 431 800 437 834
rect 391 762 437 800
rect 391 728 397 762
rect 431 728 437 762
rect 391 690 437 728
rect 391 656 397 690
rect 431 656 437 690
rect 391 618 437 656
rect 391 584 397 618
rect 431 584 437 618
rect 391 546 437 584
rect 391 512 397 546
rect 431 512 437 546
rect 391 474 437 512
rect 391 440 397 474
rect 431 440 437 474
rect 391 402 437 440
rect 391 368 397 402
rect 431 368 437 402
rect 391 330 437 368
rect 391 296 397 330
rect 431 296 437 330
rect 391 258 437 296
rect 391 224 397 258
rect 431 224 437 258
rect 391 212 437 224
rect 547 1194 593 1206
rect 547 1160 553 1194
rect 587 1160 593 1194
rect 547 1122 593 1160
rect 547 1088 553 1122
rect 587 1088 593 1122
rect 547 1050 593 1088
rect 547 1016 553 1050
rect 587 1016 593 1050
rect 547 978 593 1016
rect 547 944 553 978
rect 587 944 593 978
rect 547 906 593 944
rect 547 872 553 906
rect 587 872 593 906
rect 547 834 593 872
rect 547 800 553 834
rect 587 800 593 834
rect 547 762 593 800
rect 547 728 553 762
rect 587 728 593 762
rect 547 690 593 728
rect 547 656 553 690
rect 587 656 593 690
rect 547 618 593 656
rect 547 584 553 618
rect 587 584 593 618
rect 547 546 593 584
rect 547 512 553 546
rect 587 512 593 546
rect 547 474 593 512
rect 547 440 553 474
rect 587 440 593 474
rect 547 402 593 440
rect 547 368 553 402
rect 587 368 593 402
rect 547 330 593 368
rect 547 296 553 330
rect 587 296 593 330
rect 547 258 593 296
rect 547 224 553 258
rect 587 224 593 258
rect 547 212 593 224
rect 703 1194 749 1206
rect 703 1160 709 1194
rect 743 1160 749 1194
rect 703 1122 749 1160
rect 703 1088 709 1122
rect 743 1088 749 1122
rect 703 1050 749 1088
rect 703 1016 709 1050
rect 743 1016 749 1050
rect 703 978 749 1016
rect 703 944 709 978
rect 743 944 749 978
rect 703 906 749 944
rect 703 872 709 906
rect 743 872 749 906
rect 703 834 749 872
rect 703 800 709 834
rect 743 800 749 834
rect 703 762 749 800
rect 703 728 709 762
rect 743 728 749 762
rect 703 690 749 728
rect 703 656 709 690
rect 743 656 749 690
rect 703 618 749 656
rect 703 584 709 618
rect 743 584 749 618
rect 703 546 749 584
rect 703 512 709 546
rect 743 512 749 546
rect 703 474 749 512
rect 703 440 709 474
rect 743 440 749 474
rect 703 402 749 440
rect 703 368 709 402
rect 743 368 749 402
rect 703 330 749 368
rect 703 296 709 330
rect 743 296 749 330
rect 703 258 749 296
rect 703 224 709 258
rect 743 224 749 258
rect 703 212 749 224
rect 859 1194 905 1293
rect 859 1160 865 1194
rect 899 1160 905 1194
rect 859 1122 905 1160
rect 859 1088 865 1122
rect 899 1088 905 1122
rect 859 1050 905 1088
rect 859 1016 865 1050
rect 899 1016 905 1050
rect 859 978 905 1016
rect 859 944 865 978
rect 899 944 905 978
rect 859 906 905 944
rect 859 872 865 906
rect 899 872 905 906
rect 859 834 905 872
rect 859 800 865 834
rect 899 800 905 834
rect 859 762 905 800
rect 859 728 865 762
rect 899 728 905 762
rect 859 690 905 728
rect 859 656 865 690
rect 899 656 905 690
rect 859 618 905 656
rect 859 584 865 618
rect 899 584 905 618
rect 859 546 905 584
rect 859 512 865 546
rect 899 512 905 546
rect 859 474 905 512
rect 859 440 865 474
rect 899 440 905 474
rect 859 402 905 440
rect 859 368 865 402
rect 899 368 905 402
rect 859 330 905 368
rect 859 296 865 330
rect 899 296 905 330
rect 859 258 905 296
rect 859 224 865 258
rect 899 224 905 258
rect 859 212 905 224
rect 309 147 320 181
rect 354 147 363 181
rect 309 109 363 147
rect 309 75 320 109
rect 354 75 363 109
rect 309 33 363 75
use sky130_fd_pr__pfet_01v8__example_55959141808451  sky130_fd_pr__pfet_01v8__example_55959141808451_0
timestamp 1619729480
transform 1 0 779 0 -1 1650
box -46 0 128 29
use sky130_fd_pr__pfet_01v8__example_55959141808450  sky130_fd_pr__pfet_01v8__example_55959141808450_0
timestamp 1619729480
transform -1 0 705 0 -1 1650
box -28 0 324 85
use sky130_fd_pr__pfet_01v8__example_55959141808457  sky130_fd_pr__pfet_01v8__example_55959141808457_0
timestamp 1619729480
transform 1 0 57 0 -1 1650
box -28 0 324 85
use sky130_fd_pr__nfet_01v8__example_55959141808248  sky130_fd_pr__nfet_01v8__example_55959141808248_0
timestamp 1619729480
transform 1 0 754 0 1 228
box -28 0 128 481
use sky130_fd_pr__nfet_01v8__example_55959141808447  sky130_fd_pr__nfet_01v8__example_55959141808447_0
timestamp 1619729480
transform 1 0 442 0 1 228
box -28 0 128 481
use sky130_fd_pr__nfet_01v8__example_55959141808447  sky130_fd_pr__nfet_01v8__example_55959141808447_1
timestamp 1619729480
transform 1 0 598 0 1 228
box -28 0 128 481
use sky130_fd_pr__nfet_01v8__example_55959141808446  sky130_fd_pr__nfet_01v8__example_55959141808446_0
timestamp 1619729480
transform -1 0 212 0 -1 1102
box -46 0 128 29
use sky130_fd_pr__nfet_01v8__example_55959141808445  sky130_fd_pr__nfet_01v8__example_55959141808445_0
timestamp 1619729480
transform 1 0 286 0 1 228
box -28 0 128 481
use sky130_fd_pr__nfet_01v8__example_55959141808585  sky130_fd_pr__nfet_01v8__example_55959141808585_0
timestamp 1619729480
transform -1 0 212 0 1 685
box -25 0 128 42
<< labels >>
flabel metal1 s 871 1285 899 1313 3 FreeSans 280 180 0 0 OUT
flabel metal1 s 227 1732 321 1803 3 FreeSans 520 0 0 0 VPWR
flabel metal1 s 55 427 142 548 3 FreeSans 520 0 0 0 VGND
flabel locali s 788 109 816 137 3 FreeSans 280 270 0 0 IN1
flabel locali s 322 109 350 137 3 FreeSans 280 270 0 0 IN0
flabel locali s 482 109 510 137 3 FreeSans 280 270 0 0 IN3
flabel locali s 634 109 662 137 3 FreeSans 280 270 0 0 IN2
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 18702340
string GDS_START 18687962
<< end >>
