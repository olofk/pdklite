magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1285 -1110 1385 1411
<< labels >>
flabel comment s 125 150 125 150 0 FreeSans 300 0 0 0 D
flabel comment s -25 150 -25 150 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 17444760
string GDS_START 17444120
<< end >>
