* NGSPICE file created from sky130_ef_sc_hvl__fill_8.ext - technology: sky130A

.subckt sky130_ef_sc_hvl__fill_8 VNB VGND VPWR VPB
.ends

