magic
tech sky130A
magscale 1 2
timestamp 1619729573
<< checkpaint >>
rect -1326 -1283 2958 2911
<< nwell >>
rect -66 377 306 1251
rect 706 385 1000 1115
rect 1400 377 1698 1251
<< pwell >>
rect 0 1611 1632 1645
rect 0 -17 1632 17
<< scnmos >>
rect 795 151 825 299
<< scpmoshvt >>
rect 795 855 825 1079
rect 795 421 825 645
rect 881 421 911 645
<< mvnmos >>
rect 87 1337 187 1421
rect 289 1337 389 1487
rect 445 1337 545 1487
rect 601 1337 701 1487
rect 445 1127 545 1277
rect 445 635 545 785
rect 445 425 545 575
rect 87 207 187 291
rect 289 141 389 291
rect 445 141 545 291
<< mvpmos >>
rect 87 1101 187 1185
rect 87 443 187 527
<< ndiff >>
rect 742 287 795 299
rect 742 253 750 287
rect 784 253 795 287
rect 742 197 795 253
rect 742 163 750 197
rect 784 163 795 197
rect 742 151 795 163
rect 825 287 878 299
rect 825 253 836 287
rect 870 253 878 287
rect 825 197 878 253
rect 825 163 836 197
rect 870 163 878 197
rect 825 151 878 163
<< pdiff >>
rect 742 1067 795 1079
rect 742 1033 750 1067
rect 784 1033 795 1067
rect 742 984 795 1033
rect 742 950 750 984
rect 784 950 795 984
rect 742 901 795 950
rect 742 867 750 901
rect 784 867 795 901
rect 742 855 795 867
rect 825 1067 878 1079
rect 825 1033 836 1067
rect 870 1033 878 1067
rect 825 984 878 1033
rect 825 950 836 984
rect 870 950 878 984
rect 825 901 878 950
rect 825 867 836 901
rect 870 867 878 901
rect 825 855 878 867
rect 742 633 795 645
rect 742 599 750 633
rect 784 599 795 633
rect 742 550 795 599
rect 742 516 750 550
rect 784 516 795 550
rect 742 467 795 516
rect 742 433 750 467
rect 784 433 795 467
rect 742 421 795 433
rect 825 633 881 645
rect 825 599 836 633
rect 870 599 881 633
rect 825 550 881 599
rect 825 516 836 550
rect 870 516 881 550
rect 825 467 881 516
rect 825 433 836 467
rect 870 433 881 467
rect 825 421 881 433
rect 911 565 964 645
rect 911 531 922 565
rect 956 531 964 565
rect 911 467 964 531
rect 911 433 922 467
rect 956 433 964 467
rect 911 421 964 433
<< mvndiff >>
rect 202 1475 289 1487
rect 202 1441 244 1475
rect 278 1441 289 1475
rect 202 1421 289 1441
rect 30 1396 87 1421
rect 30 1362 42 1396
rect 76 1362 87 1396
rect 30 1337 87 1362
rect 187 1396 289 1421
rect 187 1362 198 1396
rect 232 1362 289 1396
rect 187 1337 289 1362
rect 389 1475 445 1487
rect 389 1441 400 1475
rect 434 1441 445 1475
rect 389 1383 445 1441
rect 389 1349 400 1383
rect 434 1349 445 1383
rect 389 1337 445 1349
rect 545 1475 601 1487
rect 545 1441 556 1475
rect 590 1441 601 1475
rect 545 1383 601 1441
rect 545 1349 556 1383
rect 590 1349 601 1383
rect 545 1337 601 1349
rect 701 1475 754 1487
rect 701 1441 712 1475
rect 746 1441 754 1475
rect 701 1383 754 1441
rect 701 1349 712 1383
rect 746 1349 754 1383
rect 701 1337 754 1349
rect 392 1265 445 1277
rect 392 1231 400 1265
rect 434 1231 445 1265
rect 392 1173 445 1231
rect 392 1139 400 1173
rect 434 1139 445 1173
rect 392 1127 445 1139
rect 545 1265 598 1277
rect 545 1231 556 1265
rect 590 1231 598 1265
rect 545 1173 598 1231
rect 545 1139 556 1173
rect 590 1139 598 1173
rect 545 1127 598 1139
rect 392 769 445 785
rect 392 735 400 769
rect 434 735 445 769
rect 392 681 445 735
rect 392 647 400 681
rect 434 647 445 681
rect 392 635 445 647
rect 545 769 598 785
rect 545 735 556 769
rect 590 735 598 769
rect 545 681 598 735
rect 545 647 556 681
rect 590 647 598 681
rect 545 635 598 647
rect 392 559 445 575
rect 392 525 400 559
rect 434 525 445 559
rect 392 471 445 525
rect 392 437 400 471
rect 434 437 445 471
rect 392 425 445 437
rect 545 559 598 575
rect 545 525 556 559
rect 590 525 598 559
rect 545 471 598 525
rect 545 437 556 471
rect 590 437 598 471
rect 545 425 598 437
rect 30 266 87 291
rect 30 232 42 266
rect 76 232 87 266
rect 30 207 87 232
rect 187 266 289 291
rect 187 232 198 266
rect 232 232 289 266
rect 187 207 289 232
rect 202 187 289 207
rect 202 153 244 187
rect 278 153 289 187
rect 202 141 289 153
rect 389 275 445 291
rect 389 241 400 275
rect 434 241 445 275
rect 389 187 445 241
rect 389 153 400 187
rect 434 153 445 187
rect 389 141 445 153
rect 545 275 598 291
rect 545 241 556 275
rect 590 241 598 275
rect 545 187 598 241
rect 545 153 556 187
rect 590 153 598 187
rect 545 141 598 153
<< mvpdiff >>
rect 30 1160 87 1185
rect 30 1126 42 1160
rect 76 1126 87 1160
rect 30 1101 87 1126
rect 187 1160 240 1185
rect 187 1126 198 1160
rect 232 1126 240 1160
rect 187 1101 240 1126
rect 30 502 87 527
rect 30 468 42 502
rect 76 468 87 502
rect 30 443 87 468
rect 187 502 240 527
rect 187 468 198 502
rect 232 468 240 502
rect 187 443 240 468
<< ndiffc >>
rect 750 253 784 287
rect 750 163 784 197
rect 836 253 870 287
rect 836 163 870 197
<< pdiffc >>
rect 750 1033 784 1067
rect 750 950 784 984
rect 750 867 784 901
rect 836 1033 870 1067
rect 836 950 870 984
rect 836 867 870 901
rect 750 599 784 633
rect 750 516 784 550
rect 750 433 784 467
rect 836 599 870 633
rect 836 516 870 550
rect 836 433 870 467
rect 922 531 956 565
rect 922 433 956 467
<< mvndiffc >>
rect 244 1441 278 1475
rect 42 1362 76 1396
rect 198 1362 232 1396
rect 400 1441 434 1475
rect 400 1349 434 1383
rect 556 1441 590 1475
rect 556 1349 590 1383
rect 712 1441 746 1475
rect 712 1349 746 1383
rect 400 1231 434 1265
rect 400 1139 434 1173
rect 556 1231 590 1265
rect 556 1139 590 1173
rect 400 735 434 769
rect 400 647 434 681
rect 556 735 590 769
rect 556 647 590 681
rect 400 525 434 559
rect 400 437 434 471
rect 556 525 590 559
rect 556 437 590 471
rect 42 232 76 266
rect 198 232 232 266
rect 244 153 278 187
rect 400 241 434 275
rect 400 153 434 187
rect 556 241 590 275
rect 556 153 590 187
<< mvpdiffc >>
rect 42 1126 76 1160
rect 198 1126 232 1160
rect 42 468 76 502
rect 198 468 232 502
<< nsubdiff >>
rect 742 767 766 801
rect 800 767 836 801
rect 870 767 906 801
rect 940 767 964 801
rect 742 733 964 767
rect 742 699 766 733
rect 800 699 836 733
rect 870 699 906 733
rect 940 699 964 733
<< mvpsubdiff >>
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1632 1645
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 240 831
rect 1466 797 1490 831
rect 1524 797 1567 831
rect 1601 797 1632 831
<< nsubdiffcont >>
rect 766 767 800 801
rect 836 767 870 801
rect 906 767 940 801
rect 766 699 800 733
rect 836 699 870 733
rect 906 699 940 733
<< mvpsubdiffcont >>
rect 31 1611 65 1645
rect 127 1611 161 1645
rect 223 1611 257 1645
rect 319 1611 353 1645
rect 415 1611 449 1645
rect 511 1611 545 1645
rect 607 1611 641 1645
rect 703 1611 737 1645
rect 799 1611 833 1645
rect 895 1611 929 1645
rect 991 1611 1025 1645
rect 1087 1611 1121 1645
rect 1183 1611 1217 1645
rect 1279 1611 1313 1645
rect 1375 1611 1409 1645
rect 1471 1611 1505 1645
rect 1567 1611 1601 1645
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 1490 797 1524 831
rect 1567 797 1601 831
<< poly >>
rect 289 1487 389 1513
rect 445 1487 545 1513
rect 601 1487 701 1513
rect 87 1421 187 1474
rect 87 1185 187 1337
rect 289 1322 389 1337
rect 445 1322 545 1337
rect 601 1322 701 1337
rect 289 1299 701 1322
rect 289 1265 305 1299
rect 339 1292 701 1299
rect 339 1265 355 1292
rect 445 1277 545 1292
rect 289 1231 355 1265
rect 289 1197 305 1231
rect 339 1197 355 1231
rect 289 1181 355 1197
rect 743 1161 877 1177
rect 743 1127 759 1161
rect 793 1127 827 1161
rect 861 1127 877 1161
rect 445 1101 545 1127
rect 743 1111 877 1127
rect 87 1075 187 1101
rect 795 1079 825 1111
rect 126 1040 187 1075
rect 126 1024 260 1040
rect 126 990 142 1024
rect 176 990 210 1024
rect 244 990 260 1024
rect 126 974 260 990
rect 566 903 700 919
rect 566 869 582 903
rect 616 869 650 903
rect 684 869 700 903
rect 566 853 700 869
rect 445 785 545 811
rect 126 609 260 625
rect 126 575 142 609
rect 176 575 210 609
rect 244 575 260 609
rect 445 575 545 635
rect 126 559 260 575
rect 126 553 187 559
rect 87 527 187 553
rect 87 291 187 443
rect 289 431 355 447
rect 289 397 305 431
rect 339 397 355 431
rect 289 396 355 397
rect 445 396 545 425
rect 289 363 545 396
rect 289 329 305 363
rect 339 330 545 363
rect 339 329 389 330
rect 289 291 389 329
rect 445 291 545 330
rect 634 393 700 853
rect 795 829 825 855
rect 795 645 825 671
rect 881 645 911 671
rect 795 393 825 421
rect 881 393 911 421
rect 634 327 911 393
rect 795 299 825 327
rect 87 181 187 207
rect 289 115 389 141
rect 445 115 545 141
rect 795 125 825 151
<< polycont >>
rect 305 1265 339 1299
rect 305 1197 339 1231
rect 759 1127 793 1161
rect 827 1127 861 1161
rect 142 990 176 1024
rect 210 990 244 1024
rect 582 869 616 903
rect 650 869 684 903
rect 142 575 176 609
rect 210 575 244 609
rect 305 397 339 431
rect 305 329 339 363
<< locali >>
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1632 1645
rect 179 1543 297 1549
rect 179 1509 185 1543
rect 219 1509 257 1543
rect 291 1509 297 1543
rect 179 1475 297 1509
rect 506 1543 624 1549
rect 506 1509 512 1543
rect 546 1509 584 1543
rect 618 1509 624 1543
rect 179 1441 244 1475
rect 278 1441 297 1475
rect 34 1396 84 1412
rect 34 1362 42 1396
rect 76 1362 84 1396
rect 34 1315 84 1362
rect 179 1396 297 1441
rect 179 1362 198 1396
rect 232 1362 297 1396
rect 179 1349 297 1362
rect 384 1475 450 1491
rect 384 1441 400 1475
rect 434 1441 450 1475
rect 384 1383 450 1441
rect 384 1349 400 1383
rect 434 1349 450 1383
rect 34 1299 350 1315
rect 34 1265 305 1299
rect 339 1265 350 1299
rect 34 1244 350 1265
rect 190 1231 350 1244
rect 190 1197 305 1231
rect 339 1197 350 1231
rect 26 1160 92 1176
rect 26 1126 42 1160
rect 76 1126 92 1160
rect 26 939 92 1126
rect 190 1160 350 1197
rect 190 1126 198 1160
rect 232 1126 350 1160
rect 190 1110 350 1126
rect 126 1024 260 1040
rect 126 990 142 1024
rect 176 990 210 1024
rect 244 990 260 1024
rect 126 974 260 990
rect 26 933 144 939
rect 26 899 32 933
rect 66 899 104 933
rect 138 899 144 933
rect 26 893 144 899
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 177 831
rect 26 729 144 735
rect 26 695 32 729
rect 66 695 104 729
rect 138 695 144 729
rect 26 689 144 695
rect 26 502 92 689
rect 294 617 350 1110
rect 384 1265 450 1349
rect 384 1231 400 1265
rect 434 1231 450 1265
rect 384 1173 450 1231
rect 384 1139 400 1173
rect 434 1139 450 1173
rect 384 1089 450 1139
rect 506 1475 624 1509
rect 506 1441 556 1475
rect 590 1441 624 1475
rect 506 1383 624 1441
rect 506 1349 556 1383
rect 590 1349 624 1383
rect 506 1265 624 1349
rect 506 1231 556 1265
rect 590 1231 624 1265
rect 506 1173 624 1231
rect 506 1139 556 1173
rect 590 1139 624 1173
rect 696 1475 762 1491
rect 696 1441 712 1475
rect 746 1441 762 1475
rect 696 1383 762 1441
rect 696 1349 712 1383
rect 746 1349 762 1383
rect 696 1169 762 1349
rect 506 1123 624 1139
rect 658 1161 1034 1169
rect 658 1127 759 1161
rect 793 1127 827 1161
rect 861 1127 1034 1161
rect 658 1119 1034 1127
rect 658 1089 708 1119
rect 384 1039 708 1089
rect 742 1067 792 1083
rect 742 1033 750 1067
rect 784 1033 792 1067
rect 742 984 792 1033
rect 742 950 750 984
rect 784 950 792 984
rect 742 919 792 950
rect 126 609 350 617
rect 126 575 142 609
rect 176 575 210 609
rect 244 575 350 609
rect 126 567 350 575
rect 384 903 792 919
rect 384 869 582 903
rect 616 869 650 903
rect 684 901 792 903
rect 684 869 750 901
rect 384 867 750 869
rect 784 867 792 901
rect 384 851 792 867
rect 826 1067 880 1083
rect 826 1033 836 1067
rect 870 1033 880 1067
rect 826 984 880 1033
rect 826 950 836 984
rect 870 950 880 984
rect 826 901 880 950
rect 826 867 836 901
rect 870 867 880 901
rect 384 769 450 851
rect 826 817 880 867
rect 756 801 950 817
rect 384 735 400 769
rect 434 735 450 769
rect 384 681 450 735
rect 384 647 400 681
rect 434 647 450 681
rect 384 559 450 647
rect 384 525 400 559
rect 434 525 450 559
rect 26 468 42 502
rect 76 468 92 502
rect 26 452 92 468
rect 190 502 240 518
rect 190 468 198 502
rect 232 468 240 502
rect 190 379 240 468
rect 384 471 450 525
rect 289 431 350 447
rect 289 397 305 431
rect 339 397 350 431
rect 289 379 350 397
rect 34 363 350 379
rect 34 329 305 363
rect 339 329 350 363
rect 34 313 350 329
rect 384 437 400 471
rect 434 437 450 471
rect 34 266 84 313
rect 34 232 42 266
rect 76 232 84 266
rect 34 216 84 232
rect 179 266 297 279
rect 179 232 198 266
rect 232 232 297 266
rect 179 187 297 232
rect 179 153 244 187
rect 278 153 297 187
rect 179 119 297 153
rect 384 275 450 437
rect 384 241 400 275
rect 434 241 450 275
rect 384 187 450 241
rect 384 153 400 187
rect 434 153 450 187
rect 384 137 450 153
rect 514 769 632 782
rect 514 735 556 769
rect 590 735 632 769
rect 514 681 632 735
rect 756 767 766 801
rect 800 767 836 801
rect 870 767 906 801
rect 940 767 950 801
rect 756 733 950 767
rect 756 699 766 733
rect 800 699 836 733
rect 870 699 906 733
rect 940 699 950 733
rect 756 683 950 699
rect 514 647 556 681
rect 590 647 632 681
rect 826 655 950 683
rect 514 559 632 647
rect 514 525 556 559
rect 590 525 632 559
rect 514 471 632 525
rect 514 437 556 471
rect 590 437 632 471
rect 514 275 632 437
rect 514 241 556 275
rect 590 241 632 275
rect 514 187 632 241
rect 514 153 556 187
rect 590 153 632 187
rect 179 85 185 119
rect 219 85 257 119
rect 291 85 297 119
rect 179 79 297 85
rect 514 119 632 153
rect 697 633 792 649
rect 697 599 750 633
rect 784 599 792 633
rect 697 550 792 599
rect 697 516 750 550
rect 784 516 792 550
rect 697 467 792 516
rect 697 433 750 467
rect 784 433 792 467
rect 697 287 792 433
rect 826 621 832 655
rect 866 633 904 655
rect 870 621 904 633
rect 938 621 950 655
rect 826 599 836 621
rect 870 615 950 621
rect 870 599 880 615
rect 826 550 880 599
rect 984 581 1034 1119
rect 1455 797 1471 831
rect 1524 797 1567 831
rect 1601 797 1632 831
rect 826 516 836 550
rect 870 516 880 550
rect 826 467 880 516
rect 826 433 836 467
rect 870 433 880 467
rect 826 417 880 433
rect 914 565 1034 581
rect 914 531 922 565
rect 956 531 1034 565
rect 914 467 964 531
rect 914 433 922 467
rect 956 433 964 467
rect 914 417 964 433
rect 697 253 750 287
rect 784 253 792 287
rect 697 197 792 253
rect 697 163 750 197
rect 784 163 792 197
rect 697 147 792 163
rect 826 287 944 303
rect 826 253 836 287
rect 870 253 944 287
rect 826 197 944 253
rect 826 163 836 197
rect 870 163 944 197
rect 514 85 520 119
rect 554 85 592 119
rect 626 85 632 119
rect 514 79 632 85
rect 826 119 944 163
rect 826 85 832 119
rect 866 85 904 119
rect 938 85 944 119
rect 826 79 944 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 1611 65 1645
rect 127 1611 161 1645
rect 223 1611 257 1645
rect 319 1611 353 1645
rect 415 1611 449 1645
rect 511 1611 545 1645
rect 607 1611 641 1645
rect 703 1611 737 1645
rect 799 1611 833 1645
rect 895 1611 929 1645
rect 991 1611 1025 1645
rect 1087 1611 1121 1645
rect 1183 1611 1217 1645
rect 1279 1611 1313 1645
rect 1375 1611 1409 1645
rect 1471 1611 1505 1645
rect 1567 1611 1601 1645
rect 185 1509 219 1543
rect 257 1509 291 1543
rect 512 1509 546 1543
rect 584 1509 618 1543
rect 32 899 66 933
rect 104 899 138 933
rect 31 797 65 831
rect 127 797 161 831
rect 32 695 66 729
rect 104 695 138 729
rect 185 85 219 119
rect 257 85 291 119
rect 832 633 866 655
rect 832 621 836 633
rect 836 621 866 633
rect 904 621 938 655
rect 1471 797 1490 831
rect 1490 797 1505 831
rect 1567 797 1601 831
rect 520 85 554 119
rect 592 85 626 119
rect 832 85 866 119
rect 904 85 938 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 1645 1632 1651
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1632 1645
rect 0 1605 1632 1611
rect 0 1543 1632 1577
rect 0 1509 185 1543
rect 219 1509 257 1543
rect 291 1509 512 1543
rect 546 1509 584 1543
rect 618 1509 1632 1543
rect 0 1503 1632 1509
rect 0 933 1632 939
rect 0 899 32 933
rect 66 899 104 933
rect 138 899 1632 933
rect 0 865 1632 899
rect 0 831 1632 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1632 831
rect 0 791 1632 797
rect 0 729 1632 763
rect 0 695 32 729
rect 66 695 104 729
rect 138 695 1632 729
rect 0 689 1632 695
rect 14 655 1618 661
rect 14 621 832 655
rect 866 621 904 655
rect 938 621 1618 655
rect 14 604 1618 621
rect 0 119 1632 125
rect 0 85 185 119
rect 219 85 257 119
rect 291 85 520 119
rect 554 85 592 119
rect 626 85 832 119
rect 866 85 904 119
rect 938 85 1632 119
rect 0 51 1632 85
rect 0 17 1632 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -23 1632 -17
<< labels >>
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 127 982 161 1016 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 982 257 1016 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
rlabel comment s 0 0 0 0 4 lsbuflv2hv_1
flabel comment s 636 470 636 470 0 FreeSans 200 90 0 0 cross2
flabel metal1 s 0 689 1632 763 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 865 1632 939 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 1503 1632 1577 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 51 1632 125 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 0 1632 23 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 14 604 1618 661 0 FreeSans 340 0 0 0 LVPWR
port 2 nsew power bidirectional
flabel metal1 s 0 791 1632 837 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 0 1605 1632 1628 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
<< properties >>
string LEFsite unithvdbl
string LEFclass CORE
string FIXED_BBOX 0 0 1632 1628
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string LEFsymmetry X Y
string GDS_END 297540
string GDS_START 278850
<< end >>
