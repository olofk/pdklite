magic
tech sky130A
magscale 1 2
timestamp 1640697980
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 1 21 551 183
rect 29 -17 63 21
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 17 309 535 527
rect 17 171 259 275
rect 293 205 535 309
rect 17 17 535 171
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel metal1 s 0 -48 552 48 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 489 -17 523 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 397 -17 431 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 305 -17 339 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 213 -17 247 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 121 -17 155 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel viali s 29 -17 63 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 17 17 535 171 6 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 17 171 259 275 6 VGND
port 1 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 2 nsew ground bidirectional
rlabel pwell s 1 21 551 183 6 VNB
port 2 nsew ground bidirectional
rlabel nwell s -38 261 590 582 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 489 527 523 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 397 527 431 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 305 527 339 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 213 527 247 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 121 527 155 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel viali s 29 527 63 561 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 293 205 535 309 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 17 309 535 527 6 VPWR
port 4 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3296048
string GDS_START 3292962
<< end >>
