magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1511 -1250 8782 4971
<< nwell >>
rect 2009 2487 2390 3309
rect 81 513 262 1767
rect 1316 1759 2628 1767
rect 1316 1193 2743 1759
rect 5233 1388 5375 1759
rect 5233 1222 5268 1388
rect 317 1087 2743 1193
rect 2773 1087 5203 1193
rect 1316 521 2743 1087
rect 1316 440 2628 521
<< pwell >>
rect 2095 3677 2311 3711
rect 306 2112 1313 2146
rect 2784 2138 3714 2285
rect 2784 2104 5170 2138
rect 317 117 1247 151
rect 2805 142 5167 176
<< psubdiff >>
rect 2095 3677 2119 3711
rect 2153 3677 2253 3711
rect 2287 3677 2311 3711
<< mvpsubdiff >>
rect 2784 2251 2840 2285
rect 2874 2251 2908 2285
rect 2942 2251 2976 2285
rect 3010 2251 3044 2285
rect 3078 2251 3112 2285
rect 3146 2251 3180 2285
rect 3214 2251 3248 2285
rect 3282 2251 3316 2285
rect 3350 2251 3384 2285
rect 3418 2251 3452 2285
rect 3486 2251 3520 2285
rect 3554 2251 3588 2285
rect 3622 2251 3656 2285
rect 3690 2251 3714 2285
rect 2784 2211 3714 2251
rect 2784 2177 2840 2211
rect 2874 2177 2908 2211
rect 2942 2177 2976 2211
rect 3010 2177 3044 2211
rect 3078 2177 3112 2211
rect 3146 2177 3180 2211
rect 3214 2177 3248 2211
rect 3282 2177 3316 2211
rect 3350 2177 3384 2211
rect 3418 2177 3452 2211
rect 3486 2177 3520 2211
rect 3554 2177 3588 2211
rect 3622 2177 3656 2211
rect 3690 2177 3714 2211
rect 306 2112 371 2146
rect 405 2112 439 2146
rect 473 2112 507 2146
rect 541 2112 575 2146
rect 609 2112 643 2146
rect 677 2112 711 2146
rect 745 2112 779 2146
rect 813 2112 847 2146
rect 881 2112 915 2146
rect 949 2112 983 2146
rect 1017 2112 1051 2146
rect 1085 2112 1119 2146
rect 1153 2112 1187 2146
rect 1221 2112 1255 2146
rect 1289 2112 1313 2146
rect 2784 2138 3714 2177
rect 2784 2104 2868 2138
rect 2902 2104 2936 2138
rect 2970 2104 3004 2138
rect 3038 2104 3072 2138
rect 3106 2104 3140 2138
rect 3174 2104 3208 2138
rect 3242 2104 3276 2138
rect 3310 2104 3344 2138
rect 3378 2104 3412 2138
rect 3446 2104 3480 2138
rect 3514 2104 3548 2138
rect 3582 2104 3616 2138
rect 3650 2104 3684 2138
rect 3718 2104 3752 2138
rect 3786 2104 3820 2138
rect 3854 2104 3888 2138
rect 3922 2104 3956 2138
rect 3990 2104 4024 2138
rect 4058 2104 4092 2138
rect 4126 2104 4160 2138
rect 4194 2104 4228 2138
rect 4262 2104 4296 2138
rect 4330 2104 4364 2138
rect 4398 2104 4432 2138
rect 4466 2104 4500 2138
rect 4534 2104 4568 2138
rect 4602 2104 4636 2138
rect 4670 2104 4704 2138
rect 4738 2104 4772 2138
rect 4806 2104 4840 2138
rect 4874 2104 4908 2138
rect 4942 2104 4976 2138
rect 5010 2104 5044 2138
rect 5078 2104 5112 2138
rect 5146 2104 5170 2138
rect 317 117 373 151
rect 407 117 441 151
rect 475 117 509 151
rect 543 117 577 151
rect 611 117 645 151
rect 679 117 713 151
rect 747 117 781 151
rect 815 117 849 151
rect 883 117 917 151
rect 951 117 985 151
rect 1019 117 1053 151
rect 1087 117 1121 151
rect 1155 117 1189 151
rect 1223 117 1247 151
rect 2805 142 2865 176
rect 2899 142 2933 176
rect 2967 142 3001 176
rect 3035 142 3069 176
rect 3103 142 3137 176
rect 3171 142 3205 176
rect 3239 142 3273 176
rect 3307 142 3341 176
rect 3375 142 3409 176
rect 3443 142 3477 176
rect 3511 142 3545 176
rect 3579 142 3613 176
rect 3647 142 3681 176
rect 3715 142 3749 176
rect 3783 142 3817 176
rect 3851 142 3885 176
rect 3919 142 3953 176
rect 3987 142 4021 176
rect 4055 142 4089 176
rect 4123 142 4157 176
rect 4191 142 4225 176
rect 4259 142 4293 176
rect 4327 142 4361 176
rect 4395 142 4429 176
rect 4463 142 4497 176
rect 4531 142 4565 176
rect 4599 142 4633 176
rect 4667 142 4701 176
rect 4735 142 4769 176
rect 4803 142 4837 176
rect 4871 142 4905 176
rect 4939 142 4973 176
rect 5007 142 5041 176
rect 5075 142 5109 176
rect 5143 142 5167 176
<< mvnsubdiff >>
rect 2075 2621 2099 2655
rect 2133 2621 2183 2655
rect 2217 2621 2266 2655
rect 2300 2621 2324 2655
rect 2075 2587 2324 2621
rect 2075 2553 2099 2587
rect 2133 2553 2183 2587
rect 2217 2553 2266 2587
rect 2300 2553 2324 2587
rect 353 1123 425 1157
rect 459 1123 493 1157
rect 527 1123 561 1157
rect 595 1123 629 1157
rect 663 1123 697 1157
rect 731 1123 765 1157
rect 799 1123 833 1157
rect 867 1123 901 1157
rect 935 1123 969 1157
rect 1003 1123 1037 1157
rect 1071 1123 1105 1157
rect 1139 1123 1173 1157
rect 1207 1123 1241 1157
rect 1275 1123 1309 1157
rect 1343 1123 1377 1157
rect 1411 1123 1515 1157
rect 1549 1123 1583 1157
rect 1617 1123 1651 1157
rect 1685 1123 1719 1157
rect 1753 1123 1787 1157
rect 1821 1123 1855 1157
rect 1889 1123 1923 1157
rect 1957 1123 1991 1157
rect 2025 1123 2059 1157
rect 2093 1123 2127 1157
rect 2161 1123 2195 1157
rect 2229 1123 2263 1157
rect 2297 1123 2331 1157
rect 2365 1123 2399 1157
rect 2433 1123 2467 1157
rect 2501 1123 2532 1157
rect 2809 1123 2865 1157
rect 2899 1123 2933 1157
rect 2967 1123 3001 1157
rect 3035 1123 3069 1157
rect 3103 1123 3137 1157
rect 3171 1123 3205 1157
rect 3239 1123 3273 1157
rect 3307 1123 3341 1157
rect 3375 1123 3409 1157
rect 3443 1123 3477 1157
rect 3511 1123 3545 1157
rect 3579 1123 3613 1157
rect 3647 1123 3681 1157
rect 3715 1123 3749 1157
rect 3783 1123 3817 1157
rect 3851 1123 3885 1157
rect 3919 1123 3953 1157
rect 3987 1123 4021 1157
rect 4055 1123 4089 1157
rect 4123 1123 4157 1157
rect 4191 1123 4225 1157
rect 4259 1123 4293 1157
rect 4327 1123 4361 1157
rect 4395 1123 4429 1157
rect 4463 1123 4497 1157
rect 4531 1123 4565 1157
rect 4599 1123 4633 1157
rect 4667 1123 4701 1157
rect 4735 1123 4769 1157
rect 4803 1123 4837 1157
rect 4871 1123 4905 1157
rect 4939 1123 4973 1157
rect 5007 1123 5041 1157
rect 5075 1123 5109 1157
rect 5143 1123 5167 1157
<< psubdiffcont >>
rect 2119 3677 2153 3711
rect 2253 3677 2287 3711
<< mvpsubdiffcont >>
rect 2840 2251 2874 2285
rect 2908 2251 2942 2285
rect 2976 2251 3010 2285
rect 3044 2251 3078 2285
rect 3112 2251 3146 2285
rect 3180 2251 3214 2285
rect 3248 2251 3282 2285
rect 3316 2251 3350 2285
rect 3384 2251 3418 2285
rect 3452 2251 3486 2285
rect 3520 2251 3554 2285
rect 3588 2251 3622 2285
rect 3656 2251 3690 2285
rect 2840 2177 2874 2211
rect 2908 2177 2942 2211
rect 2976 2177 3010 2211
rect 3044 2177 3078 2211
rect 3112 2177 3146 2211
rect 3180 2177 3214 2211
rect 3248 2177 3282 2211
rect 3316 2177 3350 2211
rect 3384 2177 3418 2211
rect 3452 2177 3486 2211
rect 3520 2177 3554 2211
rect 3588 2177 3622 2211
rect 3656 2177 3690 2211
rect 371 2112 405 2146
rect 439 2112 473 2146
rect 507 2112 541 2146
rect 575 2112 609 2146
rect 643 2112 677 2146
rect 711 2112 745 2146
rect 779 2112 813 2146
rect 847 2112 881 2146
rect 915 2112 949 2146
rect 983 2112 1017 2146
rect 1051 2112 1085 2146
rect 1119 2112 1153 2146
rect 1187 2112 1221 2146
rect 1255 2112 1289 2146
rect 2868 2104 2902 2138
rect 2936 2104 2970 2138
rect 3004 2104 3038 2138
rect 3072 2104 3106 2138
rect 3140 2104 3174 2138
rect 3208 2104 3242 2138
rect 3276 2104 3310 2138
rect 3344 2104 3378 2138
rect 3412 2104 3446 2138
rect 3480 2104 3514 2138
rect 3548 2104 3582 2138
rect 3616 2104 3650 2138
rect 3684 2104 3718 2138
rect 3752 2104 3786 2138
rect 3820 2104 3854 2138
rect 3888 2104 3922 2138
rect 3956 2104 3990 2138
rect 4024 2104 4058 2138
rect 4092 2104 4126 2138
rect 4160 2104 4194 2138
rect 4228 2104 4262 2138
rect 4296 2104 4330 2138
rect 4364 2104 4398 2138
rect 4432 2104 4466 2138
rect 4500 2104 4534 2138
rect 4568 2104 4602 2138
rect 4636 2104 4670 2138
rect 4704 2104 4738 2138
rect 4772 2104 4806 2138
rect 4840 2104 4874 2138
rect 4908 2104 4942 2138
rect 4976 2104 5010 2138
rect 5044 2104 5078 2138
rect 5112 2104 5146 2138
rect 373 117 407 151
rect 441 117 475 151
rect 509 117 543 151
rect 577 117 611 151
rect 645 117 679 151
rect 713 117 747 151
rect 781 117 815 151
rect 849 117 883 151
rect 917 117 951 151
rect 985 117 1019 151
rect 1053 117 1087 151
rect 1121 117 1155 151
rect 1189 117 1223 151
rect 2865 142 2899 176
rect 2933 142 2967 176
rect 3001 142 3035 176
rect 3069 142 3103 176
rect 3137 142 3171 176
rect 3205 142 3239 176
rect 3273 142 3307 176
rect 3341 142 3375 176
rect 3409 142 3443 176
rect 3477 142 3511 176
rect 3545 142 3579 176
rect 3613 142 3647 176
rect 3681 142 3715 176
rect 3749 142 3783 176
rect 3817 142 3851 176
rect 3885 142 3919 176
rect 3953 142 3987 176
rect 4021 142 4055 176
rect 4089 142 4123 176
rect 4157 142 4191 176
rect 4225 142 4259 176
rect 4293 142 4327 176
rect 4361 142 4395 176
rect 4429 142 4463 176
rect 4497 142 4531 176
rect 4565 142 4599 176
rect 4633 142 4667 176
rect 4701 142 4735 176
rect 4769 142 4803 176
rect 4837 142 4871 176
rect 4905 142 4939 176
rect 4973 142 5007 176
rect 5041 142 5075 176
rect 5109 142 5143 176
<< mvnsubdiffcont >>
rect 2099 2621 2133 2655
rect 2183 2621 2217 2655
rect 2266 2621 2300 2655
rect 2099 2553 2133 2587
rect 2183 2553 2217 2587
rect 2266 2553 2300 2587
rect 425 1123 459 1157
rect 493 1123 527 1157
rect 561 1123 595 1157
rect 629 1123 663 1157
rect 697 1123 731 1157
rect 765 1123 799 1157
rect 833 1123 867 1157
rect 901 1123 935 1157
rect 969 1123 1003 1157
rect 1037 1123 1071 1157
rect 1105 1123 1139 1157
rect 1173 1123 1207 1157
rect 1241 1123 1275 1157
rect 1309 1123 1343 1157
rect 1377 1123 1411 1157
rect 1515 1123 1549 1157
rect 1583 1123 1617 1157
rect 1651 1123 1685 1157
rect 1719 1123 1753 1157
rect 1787 1123 1821 1157
rect 1855 1123 1889 1157
rect 1923 1123 1957 1157
rect 1991 1123 2025 1157
rect 2059 1123 2093 1157
rect 2127 1123 2161 1157
rect 2195 1123 2229 1157
rect 2263 1123 2297 1157
rect 2331 1123 2365 1157
rect 2399 1123 2433 1157
rect 2467 1123 2501 1157
rect 2865 1123 2899 1157
rect 2933 1123 2967 1157
rect 3001 1123 3035 1157
rect 3069 1123 3103 1157
rect 3137 1123 3171 1157
rect 3205 1123 3239 1157
rect 3273 1123 3307 1157
rect 3341 1123 3375 1157
rect 3409 1123 3443 1157
rect 3477 1123 3511 1157
rect 3545 1123 3579 1157
rect 3613 1123 3647 1157
rect 3681 1123 3715 1157
rect 3749 1123 3783 1157
rect 3817 1123 3851 1157
rect 3885 1123 3919 1157
rect 3953 1123 3987 1157
rect 4021 1123 4055 1157
rect 4089 1123 4123 1157
rect 4157 1123 4191 1157
rect 4225 1123 4259 1157
rect 4293 1123 4327 1157
rect 4361 1123 4395 1157
rect 4429 1123 4463 1157
rect 4497 1123 4531 1157
rect 4565 1123 4599 1157
rect 4633 1123 4667 1157
rect 4701 1123 4735 1157
rect 4769 1123 4803 1157
rect 4837 1123 4871 1157
rect 4905 1123 4939 1157
rect 4973 1123 5007 1157
rect 5041 1123 5075 1157
rect 5109 1123 5143 1157
<< locali >>
rect 2067 3677 2119 3711
rect 2153 3677 2253 3711
rect 2287 3677 2311 3711
rect 2067 3436 2140 3677
rect 2040 2655 2140 3239
rect 2040 2621 2099 2655
rect 2133 2621 2183 2655
rect 2217 2621 2266 2655
rect 2300 2621 2324 2655
rect 2040 2587 2324 2621
rect 2040 2553 2099 2587
rect 2133 2553 2183 2587
rect 2217 2553 2266 2587
rect 2300 2553 2324 2587
rect 2784 2251 2804 2285
rect 2838 2251 2840 2285
rect 2874 2251 2876 2285
rect 2942 2251 2948 2285
rect 3010 2251 3020 2285
rect 3078 2251 3092 2285
rect 3146 2251 3164 2285
rect 3214 2251 3236 2285
rect 3282 2251 3308 2285
rect 3350 2251 3380 2285
rect 3418 2251 3452 2285
rect 3486 2251 3520 2285
rect 3558 2251 3588 2285
rect 3630 2251 3656 2285
rect 3702 2251 3714 2285
rect 2784 2211 3714 2251
rect 2784 2177 2804 2211
rect 2838 2177 2840 2211
rect 2874 2177 2876 2211
rect 2942 2177 2948 2211
rect 3010 2177 3020 2211
rect 3078 2177 3092 2211
rect 3146 2177 3164 2211
rect 3214 2177 3236 2211
rect 3282 2177 3308 2211
rect 3350 2177 3380 2211
rect 3418 2177 3452 2211
rect 3486 2177 3520 2211
rect 3558 2177 3588 2211
rect 3630 2177 3656 2211
rect 3702 2177 3714 2211
rect 306 2112 331 2146
rect 365 2112 371 2146
rect 437 2112 439 2146
rect 473 2112 475 2146
rect 541 2112 547 2146
rect 609 2112 619 2146
rect 677 2112 691 2146
rect 745 2112 763 2146
rect 813 2112 835 2146
rect 881 2112 907 2146
rect 949 2112 979 2146
rect 1017 2112 1051 2146
rect 1085 2112 1119 2146
rect 1157 2112 1187 2146
rect 1229 2112 1255 2146
rect 1301 2112 1313 2146
rect 2784 2138 3714 2177
rect 2784 2104 2820 2138
rect 2854 2104 2868 2138
rect 2926 2104 2936 2138
rect 2998 2104 3004 2138
rect 3070 2104 3072 2138
rect 3106 2104 3108 2138
rect 3174 2104 3180 2138
rect 3242 2104 3252 2138
rect 3310 2104 3324 2138
rect 3378 2104 3396 2138
rect 3446 2104 3468 2138
rect 3514 2104 3540 2138
rect 3582 2104 3612 2138
rect 3650 2104 3684 2138
rect 3718 2104 3752 2138
rect 3790 2104 3820 2138
rect 3862 2104 3888 2138
rect 3934 2104 3956 2138
rect 4006 2104 4024 2138
rect 4078 2104 4092 2138
rect 4150 2104 4160 2138
rect 4222 2104 4228 2138
rect 4294 2104 4296 2138
rect 4330 2104 4332 2138
rect 4398 2104 4404 2138
rect 4466 2104 4476 2138
rect 4534 2104 4548 2138
rect 4602 2104 4620 2138
rect 4670 2104 4692 2138
rect 4738 2104 4764 2138
rect 4806 2104 4836 2138
rect 4874 2104 4908 2138
rect 4942 2104 4976 2138
rect 5014 2104 5044 2138
rect 5086 2104 5112 2138
rect 5158 2104 5170 2138
rect -54 1778 -20 1816
rect 132 1778 166 1816
rect 685 1773 719 1811
rect 333 1627 367 1665
rect 405 1484 471 1748
rect 580 1699 642 1750
rect 949 1782 983 1820
rect 580 1665 589 1699
rect 623 1665 642 1699
rect 580 1627 642 1665
rect 580 1593 589 1627
rect 623 1593 642 1627
rect 580 1575 642 1593
rect 763 1696 827 1750
rect 1128 1781 1162 1819
rect 1758 1758 1792 1796
rect 3267 1770 3301 1808
rect 3558 1805 3592 1843
rect 4297 1802 4331 1899
rect 763 1662 783 1696
rect 817 1662 827 1696
rect 763 1624 827 1662
rect 2295 1671 2329 1709
rect 2061 1624 2099 1658
rect 2886 1689 2949 1740
rect 2886 1655 2893 1689
rect 2927 1655 2949 1689
rect 763 1590 783 1624
rect 817 1590 827 1624
rect 763 1575 827 1590
rect 2886 1617 2949 1655
rect 2886 1583 2893 1617
rect 2927 1583 2949 1617
rect 2886 1565 2949 1583
rect 3070 1689 3135 1740
rect 4101 1768 4139 1802
rect 4173 1768 4225 1802
rect 4259 1768 4297 1802
rect 4389 1807 4423 1845
rect 5023 1847 5089 1860
rect 5023 1841 5042 1847
rect 5076 1841 5089 1847
rect 5042 1775 5076 1813
rect 3070 1655 3087 1689
rect 3121 1655 3135 1689
rect 3070 1617 3135 1655
rect 3070 1583 3087 1617
rect 3121 1583 3135 1617
rect 3345 1617 3379 1655
rect 3645 1649 3679 1687
rect 3070 1565 3135 1583
rect 3714 1534 3780 1740
rect 3896 1721 3962 1741
rect 3896 1687 3911 1721
rect 3945 1687 3962 1721
rect 3896 1649 3962 1687
rect 3896 1615 3911 1649
rect 3945 1615 3962 1649
rect 3997 1571 4031 1609
rect 4542 1618 4608 1740
rect 4542 1584 4565 1618
rect 4599 1584 4608 1618
rect 4542 1546 4608 1584
rect 3714 1500 3730 1534
rect 3764 1500 3780 1534
rect 4542 1520 4565 1546
rect 4599 1520 4608 1546
rect 4845 1527 4911 1740
rect 4949 1690 4983 1728
rect 210 1405 244 1443
rect 405 1450 421 1484
rect 455 1450 471 1484
rect 405 1412 471 1450
rect 405 1378 421 1412
rect 455 1378 471 1412
rect 1196 1412 1230 1450
rect 2993 1412 3027 1450
rect 3714 1462 3780 1500
rect 3714 1428 3730 1462
rect 3764 1428 3780 1462
rect 3714 1410 3780 1428
rect 4845 1493 4864 1527
rect 4898 1493 4911 1527
rect 4845 1455 4911 1493
rect 4845 1421 4864 1455
rect 4898 1421 4911 1455
rect 4845 1417 4911 1421
rect 353 1123 425 1157
rect 475 1123 493 1157
rect 547 1123 561 1157
rect 619 1123 629 1157
rect 691 1123 697 1157
rect 763 1123 765 1157
rect 799 1123 801 1157
rect 867 1123 873 1157
rect 935 1123 945 1157
rect 1003 1123 1017 1157
rect 1071 1123 1089 1157
rect 1139 1123 1161 1157
rect 1207 1123 1233 1157
rect 1275 1123 1305 1157
rect 1343 1123 1377 1157
rect 1411 1123 1503 1157
rect 1549 1123 1575 1157
rect 1617 1123 1647 1157
rect 1685 1123 1719 1157
rect 1753 1123 1787 1157
rect 1825 1123 1855 1157
rect 1897 1123 1923 1157
rect 1969 1123 1991 1157
rect 2041 1123 2059 1157
rect 2113 1123 2127 1157
rect 2185 1123 2195 1157
rect 2257 1123 2263 1157
rect 2329 1123 2331 1157
rect 2365 1123 2367 1157
rect 2433 1123 2439 1157
rect 2501 1123 2532 1157
rect 2809 1123 2865 1157
rect 2923 1123 2933 1157
rect 2995 1123 3001 1157
rect 3067 1123 3069 1157
rect 3103 1123 3105 1157
rect 3171 1123 3177 1157
rect 3239 1123 3249 1157
rect 3307 1123 3321 1157
rect 3375 1123 3393 1157
rect 3443 1123 3465 1157
rect 3511 1123 3537 1157
rect 3579 1123 3609 1157
rect 3647 1123 3681 1157
rect 3715 1123 3749 1157
rect 3787 1123 3817 1157
rect 3859 1123 3885 1157
rect 3931 1123 3953 1157
rect 4003 1123 4021 1157
rect 4075 1123 4089 1157
rect 4147 1123 4157 1157
rect 4219 1123 4225 1157
rect 4291 1123 4293 1157
rect 4327 1123 4329 1157
rect 4395 1123 4401 1157
rect 4463 1123 4473 1157
rect 4531 1123 4545 1157
rect 4599 1123 4617 1157
rect 4667 1123 4689 1157
rect 4735 1123 4761 1157
rect 4803 1123 4833 1157
rect 4871 1123 4905 1157
rect 4939 1123 4973 1157
rect 5011 1123 5041 1157
rect 5083 1123 5109 1157
rect 5155 1123 5167 1157
rect 4848 925 4914 937
rect 685 824 719 862
rect 4848 891 4860 925
rect 4894 891 4914 925
rect 4848 853 4914 891
rect 2027 757 2065 791
rect 2993 758 3027 796
rect 3242 796 3261 830
rect 3295 796 3308 830
rect 3242 758 3308 796
rect 3242 724 3261 758
rect 3295 724 3308 758
rect 3645 765 3679 803
rect 3715 805 3737 837
rect 3771 805 3781 837
rect 3715 767 3781 805
rect 3715 733 3737 767
rect 3771 733 3781 767
rect 4121 767 4155 805
rect 4848 819 4860 853
rect 4894 819 4914 853
rect 30 681 64 719
rect 579 689 642 707
rect 332 617 366 655
rect 579 655 589 689
rect 623 655 642 689
rect 579 617 642 655
rect 579 583 589 617
rect 623 583 642 617
rect -56 461 -22 499
rect 579 532 642 583
rect 763 689 827 707
rect 763 655 783 689
rect 817 655 827 689
rect 763 617 827 655
rect 763 583 783 617
rect 817 583 827 617
rect 763 532 827 583
rect 1057 651 1075 685
rect 1109 651 1123 685
rect 1057 613 1123 651
rect 1728 650 1762 688
rect 2887 697 2949 715
rect 2887 663 2893 697
rect 2927 663 2949 697
rect 2887 625 2949 663
rect 1057 579 1075 613
rect 1109 579 1123 613
rect 119 461 153 499
rect 421 454 455 492
rect 986 502 1020 540
rect 1057 532 1123 579
rect 2887 591 2893 625
rect 2927 591 2949 625
rect 2887 540 2949 591
rect 3070 697 3134 715
rect 3070 663 3087 697
rect 3121 663 3134 697
rect 3070 625 3134 663
rect 3070 591 3087 625
rect 3121 591 3134 625
rect 3070 540 3134 591
rect 3242 540 3308 724
rect 3345 625 3379 663
rect 3715 540 3781 733
rect 4474 635 4508 673
rect 3559 483 3593 521
rect 4036 483 4070 521
rect 4372 540 4392 559
rect 4209 483 4243 521
rect 4426 540 4438 559
rect 4543 540 4561 559
rect 4392 487 4426 525
rect 4595 540 4609 559
rect 4848 540 4914 819
rect 4949 738 4983 776
rect 4561 487 4595 525
rect 5033 490 5067 528
rect 2257 276 2295 310
rect 317 117 337 151
rect 371 117 373 151
rect 407 117 409 151
rect 475 117 481 151
rect 543 117 553 151
rect 611 117 625 151
rect 679 117 697 151
rect 747 117 769 151
rect 815 117 841 151
rect 883 117 913 151
rect 951 117 985 151
rect 1019 117 1053 151
rect 1091 117 1121 151
rect 1163 117 1189 151
rect 1235 117 1247 151
rect 2805 142 2817 176
rect 2851 142 2865 176
rect 2923 142 2933 176
rect 2995 142 3001 176
rect 3067 142 3069 176
rect 3103 142 3105 176
rect 3171 142 3177 176
rect 3239 142 3249 176
rect 3307 142 3321 176
rect 3375 142 3393 176
rect 3443 142 3465 176
rect 3511 142 3537 176
rect 3579 142 3609 176
rect 3647 142 3681 176
rect 3715 142 3749 176
rect 3787 142 3817 176
rect 3859 142 3885 176
rect 3931 142 3953 176
rect 4003 142 4021 176
rect 4075 142 4089 176
rect 4147 142 4157 176
rect 4219 142 4225 176
rect 4291 142 4293 176
rect 4327 142 4329 176
rect 4395 142 4401 176
rect 4463 142 4473 176
rect 4531 142 4545 176
rect 4599 142 4617 176
rect 4667 142 4689 176
rect 4735 142 4761 176
rect 4803 142 4833 176
rect 4871 142 4905 176
rect 4939 142 4973 176
rect 5011 142 5041 176
rect 5083 142 5109 176
rect 5155 142 5167 176
<< viali >>
rect 2804 2251 2838 2285
rect 2876 2251 2908 2285
rect 2908 2251 2910 2285
rect 2948 2251 2976 2285
rect 2976 2251 2982 2285
rect 3020 2251 3044 2285
rect 3044 2251 3054 2285
rect 3092 2251 3112 2285
rect 3112 2251 3126 2285
rect 3164 2251 3180 2285
rect 3180 2251 3198 2285
rect 3236 2251 3248 2285
rect 3248 2251 3270 2285
rect 3308 2251 3316 2285
rect 3316 2251 3342 2285
rect 3380 2251 3384 2285
rect 3384 2251 3414 2285
rect 3452 2251 3486 2285
rect 3524 2251 3554 2285
rect 3554 2251 3558 2285
rect 3596 2251 3622 2285
rect 3622 2251 3630 2285
rect 3668 2251 3690 2285
rect 3690 2251 3702 2285
rect 2804 2177 2838 2211
rect 2876 2177 2908 2211
rect 2908 2177 2910 2211
rect 2948 2177 2976 2211
rect 2976 2177 2982 2211
rect 3020 2177 3044 2211
rect 3044 2177 3054 2211
rect 3092 2177 3112 2211
rect 3112 2177 3126 2211
rect 3164 2177 3180 2211
rect 3180 2177 3198 2211
rect 3236 2177 3248 2211
rect 3248 2177 3270 2211
rect 3308 2177 3316 2211
rect 3316 2177 3342 2211
rect 3380 2177 3384 2211
rect 3384 2177 3414 2211
rect 3452 2177 3486 2211
rect 3524 2177 3554 2211
rect 3554 2177 3558 2211
rect 3596 2177 3622 2211
rect 3622 2177 3630 2211
rect 3668 2177 3690 2211
rect 3690 2177 3702 2211
rect 331 2112 365 2146
rect 403 2112 405 2146
rect 405 2112 437 2146
rect 475 2112 507 2146
rect 507 2112 509 2146
rect 547 2112 575 2146
rect 575 2112 581 2146
rect 619 2112 643 2146
rect 643 2112 653 2146
rect 691 2112 711 2146
rect 711 2112 725 2146
rect 763 2112 779 2146
rect 779 2112 797 2146
rect 835 2112 847 2146
rect 847 2112 869 2146
rect 907 2112 915 2146
rect 915 2112 941 2146
rect 979 2112 983 2146
rect 983 2112 1013 2146
rect 1051 2112 1085 2146
rect 1123 2112 1153 2146
rect 1153 2112 1157 2146
rect 1195 2112 1221 2146
rect 1221 2112 1229 2146
rect 1267 2112 1289 2146
rect 1289 2112 1301 2146
rect 2820 2104 2854 2138
rect 2892 2104 2902 2138
rect 2902 2104 2926 2138
rect 2964 2104 2970 2138
rect 2970 2104 2998 2138
rect 3036 2104 3038 2138
rect 3038 2104 3070 2138
rect 3108 2104 3140 2138
rect 3140 2104 3142 2138
rect 3180 2104 3208 2138
rect 3208 2104 3214 2138
rect 3252 2104 3276 2138
rect 3276 2104 3286 2138
rect 3324 2104 3344 2138
rect 3344 2104 3358 2138
rect 3396 2104 3412 2138
rect 3412 2104 3430 2138
rect 3468 2104 3480 2138
rect 3480 2104 3502 2138
rect 3540 2104 3548 2138
rect 3548 2104 3574 2138
rect 3612 2104 3616 2138
rect 3616 2104 3646 2138
rect 3684 2104 3718 2138
rect 3756 2104 3786 2138
rect 3786 2104 3790 2138
rect 3828 2104 3854 2138
rect 3854 2104 3862 2138
rect 3900 2104 3922 2138
rect 3922 2104 3934 2138
rect 3972 2104 3990 2138
rect 3990 2104 4006 2138
rect 4044 2104 4058 2138
rect 4058 2104 4078 2138
rect 4116 2104 4126 2138
rect 4126 2104 4150 2138
rect 4188 2104 4194 2138
rect 4194 2104 4222 2138
rect 4260 2104 4262 2138
rect 4262 2104 4294 2138
rect 4332 2104 4364 2138
rect 4364 2104 4366 2138
rect 4404 2104 4432 2138
rect 4432 2104 4438 2138
rect 4476 2104 4500 2138
rect 4500 2104 4510 2138
rect 4548 2104 4568 2138
rect 4568 2104 4582 2138
rect 4620 2104 4636 2138
rect 4636 2104 4654 2138
rect 4692 2104 4704 2138
rect 4704 2104 4726 2138
rect 4764 2104 4772 2138
rect 4772 2104 4798 2138
rect 4836 2104 4840 2138
rect 4840 2104 4870 2138
rect 4908 2104 4942 2138
rect 4980 2104 5010 2138
rect 5010 2104 5014 2138
rect 5052 2104 5078 2138
rect 5078 2104 5086 2138
rect 5124 2104 5146 2138
rect 5146 2104 5158 2138
rect -54 1816 -20 1850
rect -54 1744 -20 1778
rect 132 1816 166 1850
rect 132 1744 166 1778
rect 685 1811 719 1845
rect 333 1665 367 1699
rect 333 1593 367 1627
rect 685 1739 719 1773
rect 949 1820 983 1854
rect 589 1665 623 1699
rect 589 1593 623 1627
rect 949 1748 983 1782
rect 1128 1819 1162 1853
rect 3558 1843 3592 1877
rect 1128 1747 1162 1781
rect 1758 1796 1792 1830
rect 1758 1724 1792 1758
rect 3267 1808 3301 1842
rect 3558 1771 3592 1805
rect 783 1662 817 1696
rect 2295 1709 2329 1743
rect 2027 1624 2061 1658
rect 2099 1624 2133 1658
rect 2295 1637 2329 1671
rect 2893 1655 2927 1689
rect 783 1590 817 1624
rect 2893 1583 2927 1617
rect 3267 1736 3301 1770
rect 4067 1768 4101 1802
rect 4139 1768 4173 1802
rect 4225 1768 4259 1802
rect 4297 1768 4331 1802
rect 4389 1845 4423 1879
rect 4389 1773 4423 1807
rect 5042 1813 5076 1847
rect 3087 1655 3121 1689
rect 3087 1583 3121 1617
rect 3345 1655 3379 1689
rect 3345 1583 3379 1617
rect 3645 1687 3679 1721
rect 3645 1615 3679 1649
rect 3911 1687 3945 1721
rect 3911 1615 3945 1649
rect 3997 1609 4031 1643
rect 3997 1537 4031 1571
rect 4565 1584 4599 1618
rect 3730 1500 3764 1534
rect 4565 1512 4599 1546
rect 4949 1728 4983 1762
rect 5042 1741 5076 1775
rect 4949 1656 4983 1690
rect 210 1443 244 1477
rect 210 1371 244 1405
rect 421 1450 455 1484
rect 421 1378 455 1412
rect 1196 1450 1230 1484
rect 1196 1378 1230 1412
rect 2993 1450 3027 1484
rect 2993 1378 3027 1412
rect 3730 1428 3764 1462
rect 4864 1493 4898 1527
rect 4864 1421 4898 1455
rect 441 1123 459 1157
rect 459 1123 475 1157
rect 513 1123 527 1157
rect 527 1123 547 1157
rect 585 1123 595 1157
rect 595 1123 619 1157
rect 657 1123 663 1157
rect 663 1123 691 1157
rect 729 1123 731 1157
rect 731 1123 763 1157
rect 801 1123 833 1157
rect 833 1123 835 1157
rect 873 1123 901 1157
rect 901 1123 907 1157
rect 945 1123 969 1157
rect 969 1123 979 1157
rect 1017 1123 1037 1157
rect 1037 1123 1051 1157
rect 1089 1123 1105 1157
rect 1105 1123 1123 1157
rect 1161 1123 1173 1157
rect 1173 1123 1195 1157
rect 1233 1123 1241 1157
rect 1241 1123 1267 1157
rect 1305 1123 1309 1157
rect 1309 1123 1339 1157
rect 1377 1123 1411 1157
rect 1503 1123 1515 1157
rect 1515 1123 1537 1157
rect 1575 1123 1583 1157
rect 1583 1123 1609 1157
rect 1647 1123 1651 1157
rect 1651 1123 1681 1157
rect 1719 1123 1753 1157
rect 1791 1123 1821 1157
rect 1821 1123 1825 1157
rect 1863 1123 1889 1157
rect 1889 1123 1897 1157
rect 1935 1123 1957 1157
rect 1957 1123 1969 1157
rect 2007 1123 2025 1157
rect 2025 1123 2041 1157
rect 2079 1123 2093 1157
rect 2093 1123 2113 1157
rect 2151 1123 2161 1157
rect 2161 1123 2185 1157
rect 2223 1123 2229 1157
rect 2229 1123 2257 1157
rect 2295 1123 2297 1157
rect 2297 1123 2329 1157
rect 2367 1123 2399 1157
rect 2399 1123 2401 1157
rect 2439 1123 2467 1157
rect 2467 1123 2473 1157
rect 2889 1123 2899 1157
rect 2899 1123 2923 1157
rect 2961 1123 2967 1157
rect 2967 1123 2995 1157
rect 3033 1123 3035 1157
rect 3035 1123 3067 1157
rect 3105 1123 3137 1157
rect 3137 1123 3139 1157
rect 3177 1123 3205 1157
rect 3205 1123 3211 1157
rect 3249 1123 3273 1157
rect 3273 1123 3283 1157
rect 3321 1123 3341 1157
rect 3341 1123 3355 1157
rect 3393 1123 3409 1157
rect 3409 1123 3427 1157
rect 3465 1123 3477 1157
rect 3477 1123 3499 1157
rect 3537 1123 3545 1157
rect 3545 1123 3571 1157
rect 3609 1123 3613 1157
rect 3613 1123 3643 1157
rect 3681 1123 3715 1157
rect 3753 1123 3783 1157
rect 3783 1123 3787 1157
rect 3825 1123 3851 1157
rect 3851 1123 3859 1157
rect 3897 1123 3919 1157
rect 3919 1123 3931 1157
rect 3969 1123 3987 1157
rect 3987 1123 4003 1157
rect 4041 1123 4055 1157
rect 4055 1123 4075 1157
rect 4113 1123 4123 1157
rect 4123 1123 4147 1157
rect 4185 1123 4191 1157
rect 4191 1123 4219 1157
rect 4257 1123 4259 1157
rect 4259 1123 4291 1157
rect 4329 1123 4361 1157
rect 4361 1123 4363 1157
rect 4401 1123 4429 1157
rect 4429 1123 4435 1157
rect 4473 1123 4497 1157
rect 4497 1123 4507 1157
rect 4545 1123 4565 1157
rect 4565 1123 4579 1157
rect 4617 1123 4633 1157
rect 4633 1123 4651 1157
rect 4689 1123 4701 1157
rect 4701 1123 4723 1157
rect 4761 1123 4769 1157
rect 4769 1123 4795 1157
rect 4833 1123 4837 1157
rect 4837 1123 4867 1157
rect 4905 1123 4939 1157
rect 4977 1123 5007 1157
rect 5007 1123 5011 1157
rect 5049 1123 5075 1157
rect 5075 1123 5083 1157
rect 5121 1123 5143 1157
rect 5143 1123 5155 1157
rect 685 862 719 896
rect 4860 891 4894 925
rect 685 790 719 824
rect 2993 796 3027 830
rect 1993 757 2027 791
rect 2065 757 2099 791
rect 30 719 64 753
rect 2993 724 3027 758
rect 3261 796 3295 830
rect 3261 724 3295 758
rect 3645 803 3679 837
rect 3645 731 3679 765
rect 3737 805 3771 839
rect 3737 733 3771 767
rect 4121 805 4155 839
rect 4121 733 4155 767
rect 4860 819 4894 853
rect 30 647 64 681
rect 332 655 366 689
rect 332 583 366 617
rect 589 655 623 689
rect 589 583 623 617
rect -56 499 -22 533
rect -56 427 -22 461
rect 119 499 153 533
rect 783 655 817 689
rect 1728 688 1762 722
rect 783 583 817 617
rect 1075 651 1109 685
rect 1728 616 1762 650
rect 2893 663 2927 697
rect 1075 579 1109 613
rect 986 540 1020 574
rect 119 427 153 461
rect 421 492 455 526
rect 2893 591 2927 625
rect 3087 663 3121 697
rect 3087 591 3121 625
rect 3345 663 3379 697
rect 3345 591 3379 625
rect 986 468 1020 502
rect 3559 521 3593 555
rect 4474 673 4508 707
rect 4474 601 4508 635
rect 421 420 455 454
rect 3559 449 3593 483
rect 4036 521 4070 555
rect 4036 449 4070 483
rect 4209 521 4243 555
rect 4209 449 4243 483
rect 4392 525 4426 559
rect 4392 453 4426 487
rect 4561 525 4595 559
rect 4949 776 4983 810
rect 4949 704 4983 738
rect 4561 453 4595 487
rect 5033 528 5067 562
rect 5033 456 5067 490
rect 2223 276 2257 310
rect 2295 276 2329 310
rect 337 117 371 151
rect 409 117 441 151
rect 441 117 443 151
rect 481 117 509 151
rect 509 117 515 151
rect 553 117 577 151
rect 577 117 587 151
rect 625 117 645 151
rect 645 117 659 151
rect 697 117 713 151
rect 713 117 731 151
rect 769 117 781 151
rect 781 117 803 151
rect 841 117 849 151
rect 849 117 875 151
rect 913 117 917 151
rect 917 117 947 151
rect 985 117 1019 151
rect 1057 117 1087 151
rect 1087 117 1091 151
rect 1129 117 1155 151
rect 1155 117 1163 151
rect 1201 117 1223 151
rect 1223 117 1235 151
rect 2817 142 2851 176
rect 2889 142 2899 176
rect 2899 142 2923 176
rect 2961 142 2967 176
rect 2967 142 2995 176
rect 3033 142 3035 176
rect 3035 142 3067 176
rect 3105 142 3137 176
rect 3137 142 3139 176
rect 3177 142 3205 176
rect 3205 142 3211 176
rect 3249 142 3273 176
rect 3273 142 3283 176
rect 3321 142 3341 176
rect 3341 142 3355 176
rect 3393 142 3409 176
rect 3409 142 3427 176
rect 3465 142 3477 176
rect 3477 142 3499 176
rect 3537 142 3545 176
rect 3545 142 3571 176
rect 3609 142 3613 176
rect 3613 142 3643 176
rect 3681 142 3715 176
rect 3753 142 3783 176
rect 3783 142 3787 176
rect 3825 142 3851 176
rect 3851 142 3859 176
rect 3897 142 3919 176
rect 3919 142 3931 176
rect 3969 142 3987 176
rect 3987 142 4003 176
rect 4041 142 4055 176
rect 4055 142 4075 176
rect 4113 142 4123 176
rect 4123 142 4147 176
rect 4185 142 4191 176
rect 4191 142 4219 176
rect 4257 142 4259 176
rect 4259 142 4291 176
rect 4329 142 4361 176
rect 4361 142 4363 176
rect 4401 142 4429 176
rect 4429 142 4435 176
rect 4473 142 4497 176
rect 4497 142 4507 176
rect 4545 142 4565 176
rect 4565 142 4579 176
rect 4617 142 4633 176
rect 4633 142 4651 176
rect 4689 142 4701 176
rect 4701 142 4723 176
rect 4761 142 4769 176
rect 4769 142 4795 176
rect 4833 142 4837 176
rect 4837 142 4867 176
rect 4905 142 4939 176
rect 4977 142 5007 176
rect 5007 142 5011 176
rect 5049 142 5075 176
rect 5075 142 5083 176
rect 5121 142 5143 176
rect 5143 142 5155 176
<< metal1 >>
rect 2192 3308 2231 3357
rect 2700 2797 2706 2849
rect 2758 2797 2777 2849
rect 2829 2797 3932 2849
rect 3984 2797 3996 2849
rect 4048 2797 4054 2849
rect 25 2705 31 2757
rect 83 2705 95 2757
rect 147 2705 2486 2757
rect 2538 2705 2550 2757
rect 2602 2705 2608 2757
rect 123 2613 129 2665
rect 181 2613 193 2665
rect 245 2613 2064 2665
rect 2116 2613 2128 2665
rect 2180 2613 3443 2665
rect 3495 2613 3507 2665
rect 3559 2613 4482 2665
rect 4534 2613 4546 2665
rect 4598 2613 4604 2665
rect -139 2521 -133 2573
rect -81 2521 -69 2573
rect -17 2521 1681 2573
rect 1733 2521 1745 2573
rect 1797 2521 4313 2573
rect 4365 2521 4377 2573
rect 4429 2521 4435 2573
rect 1080 2429 1413 2481
rect 1465 2429 1477 2481
rect 1529 2429 4867 2481
rect 4919 2429 4931 2481
rect 4983 2429 4989 2481
rect 1867 2337 1873 2389
rect 1925 2337 1937 2389
rect 1989 2337 4221 2389
rect 4273 2337 4285 2389
rect 4337 2337 4343 2389
rect 2784 2285 3714 2297
rect 2784 2251 2804 2285
rect 2838 2251 2876 2285
rect 2910 2251 2948 2285
rect 2982 2251 3020 2285
rect 3054 2251 3092 2285
rect 3126 2251 3164 2285
rect 3198 2251 3236 2285
rect 3270 2251 3308 2285
rect 3342 2251 3380 2285
rect 3414 2251 3452 2285
rect 3486 2251 3524 2285
rect 3558 2251 3596 2285
rect 3630 2251 3668 2285
rect 3702 2251 3714 2285
tri 2750 2211 2784 2245 se
rect 2784 2211 3714 2251
tri 2742 2203 2750 2211 se
rect 2750 2203 2804 2211
rect -175 2177 2804 2203
rect 2838 2177 2876 2211
rect 2910 2177 2948 2211
rect 2982 2177 3020 2211
rect 3054 2177 3092 2211
rect 3126 2177 3164 2211
rect 3198 2177 3236 2211
rect 3270 2177 3308 2211
rect 3342 2177 3380 2211
rect 3414 2177 3452 2211
rect 3486 2177 3524 2211
rect 3558 2177 3596 2211
rect 3630 2177 3668 2211
rect 3702 2177 3714 2211
rect -175 2150 3714 2177
tri 3714 2150 3861 2297 sw
rect -175 2146 5170 2150
rect -175 2112 331 2146
rect 365 2112 403 2146
rect 437 2112 475 2146
rect 509 2112 547 2146
rect 581 2112 619 2146
rect 653 2112 691 2146
rect 725 2112 763 2146
rect 797 2112 835 2146
rect 869 2112 907 2146
rect 941 2112 979 2146
rect 1013 2112 1051 2146
rect 1085 2112 1123 2146
rect 1157 2112 1195 2146
rect 1229 2112 1267 2146
rect 1301 2138 5170 2146
rect 1301 2112 2820 2138
rect -175 2104 2820 2112
rect 2854 2104 2892 2138
rect 2926 2104 2964 2138
rect 2998 2104 3036 2138
rect 3070 2104 3108 2138
rect 3142 2104 3180 2138
rect 3214 2104 3252 2138
rect 3286 2104 3324 2138
rect 3358 2104 3396 2138
rect 3430 2104 3468 2138
rect 3502 2104 3540 2138
rect 3574 2104 3612 2138
rect 3646 2104 3684 2138
rect 3718 2104 3756 2138
rect 3790 2104 3828 2138
rect 3862 2104 3900 2138
rect 3934 2104 3972 2138
rect 4006 2104 4044 2138
rect 4078 2104 4116 2138
rect 4150 2104 4188 2138
rect 4222 2104 4260 2138
rect 4294 2104 4332 2138
rect 4366 2104 4404 2138
rect 4438 2104 4476 2138
rect 4510 2104 4548 2138
rect 4582 2104 4620 2138
rect 4654 2104 4692 2138
rect 4726 2104 4764 2138
rect 4798 2104 4836 2138
rect 4870 2104 4908 2138
rect 4942 2104 4980 2138
rect 5014 2104 5052 2138
rect 5086 2104 5124 2138
rect 5158 2104 5170 2138
rect -175 2092 5170 2104
tri 5341 2097 5375 2131 nw
rect -175 2071 2809 2092
rect -175 1943 279 2071
rect 358 2015 525 2071
rect 1260 2040 2809 2071
rect 1260 2015 1293 2040
tri 1293 2015 1318 2040 nw
tri 2742 2015 2767 2040 ne
rect 2767 2015 2784 2040
tri 1260 1982 1293 2015 nw
tri 2767 1998 2784 2015 ne
rect 4250 1935 4254 2092
rect 4733 1935 4740 2092
rect 3630 1898 3682 1904
rect 3466 1881 3598 1893
rect -63 1856 -11 1862
rect -63 1792 -11 1804
rect -63 1732 -11 1740
rect 123 1856 175 1862
rect 123 1792 175 1804
rect 123 1732 175 1740
rect 679 1845 756 1857
rect 679 1811 685 1845
rect 719 1811 756 1845
rect 679 1773 756 1811
rect 679 1739 685 1773
rect 719 1739 756 1773
rect 679 1727 756 1739
rect 943 1854 989 1866
rect 943 1820 949 1854
rect 983 1820 989 1854
rect 943 1782 989 1820
rect 943 1748 949 1782
rect 983 1748 989 1782
rect 943 1727 989 1748
rect 1122 1854 1168 1865
tri 1168 1854 1173 1859 sw
rect 1122 1853 1173 1854
rect 1122 1819 1128 1853
rect 1162 1843 1173 1853
tri 1173 1843 1184 1854 sw
rect 3257 1848 3309 1854
rect 1162 1842 1184 1843
tri 1184 1842 1185 1843 sw
rect 1162 1839 1185 1842
tri 1185 1839 1188 1842 sw
rect 1162 1830 1188 1839
tri 1188 1830 1197 1839 sw
rect 1585 1833 1637 1839
rect 1162 1819 1197 1830
tri 1197 1819 1208 1830 sw
rect 1122 1796 1208 1819
tri 1208 1796 1231 1819 sw
tri 1562 1796 1585 1819 se
rect 1122 1794 1231 1796
tri 1231 1794 1233 1796 sw
tri 1560 1794 1562 1796 se
rect 1562 1794 1585 1796
rect 1122 1781 1585 1794
rect 1122 1747 1128 1781
rect 1162 1769 1637 1781
rect 1162 1756 1585 1769
rect 1162 1747 1168 1756
tri 1168 1753 1171 1756 nw
tri 1541 1753 1544 1756 ne
rect 1544 1753 1585 1756
rect 1122 1735 1168 1747
tri 1544 1735 1562 1753 ne
rect 1562 1735 1585 1753
tri 1562 1729 1568 1735 ne
rect 1568 1729 1585 1735
tri 989 1727 991 1729 sw
tri 1568 1727 1570 1729 ne
rect 1570 1727 1585 1729
rect 943 1724 991 1727
tri 991 1724 994 1727 sw
tri 1570 1724 1573 1727 ne
rect 1573 1724 1585 1727
rect 943 1711 994 1724
tri 994 1711 1007 1724 sw
tri 1573 1712 1585 1724 ne
rect 1585 1711 1637 1717
rect 1752 1830 1798 1842
rect 1752 1796 1758 1830
rect 1792 1796 1798 1830
rect 1752 1771 1798 1796
tri 1798 1771 1825 1798 sw
rect 3257 1777 3309 1796
rect 1752 1770 1825 1771
tri 1825 1770 1826 1771 sw
rect 1752 1764 1826 1770
tri 1826 1764 1832 1770 sw
rect 1752 1758 2048 1764
rect 1752 1724 1758 1758
rect 1792 1724 2048 1758
rect 1752 1712 2048 1724
rect 2100 1712 2112 1764
rect 2164 1712 2170 1764
rect 2289 1753 2335 1755
tri 2335 1753 2337 1755 sw
rect 2289 1743 2337 1753
rect 327 1699 373 1711
tri 581 1709 583 1711 se
rect 583 1709 629 1711
tri 629 1709 631 1711 sw
rect 943 1709 1007 1711
tri 1007 1709 1009 1711 sw
rect 2289 1709 2295 1743
rect 2329 1736 2337 1743
tri 2337 1736 2354 1753 sw
tri 2507 1736 2524 1753 se
rect 2524 1747 2576 1753
rect 2329 1732 2354 1736
tri 2354 1732 2358 1736 sw
tri 2503 1732 2507 1736 se
rect 2507 1732 2524 1736
rect 2329 1709 2524 1732
tri 577 1705 581 1709 se
rect 581 1708 631 1709
tri 631 1708 632 1709 sw
rect 943 1708 1009 1709
tri 1009 1708 1010 1709 sw
rect 581 1706 632 1708
tri 632 1706 634 1708 sw
rect 581 1705 634 1706
tri 373 1699 379 1705 sw
tri 571 1699 577 1705 se
rect 577 1699 634 1705
rect 327 1665 333 1699
rect 367 1672 379 1699
tri 379 1672 406 1699 sw
tri 544 1672 571 1699 se
rect 571 1672 589 1699
rect 367 1665 589 1672
rect 623 1696 634 1699
tri 634 1696 644 1706 sw
tri 767 1696 777 1706 se
rect 777 1696 823 1708
rect 623 1672 644 1696
tri 644 1672 668 1696 sw
tri 743 1672 767 1696 se
rect 767 1672 783 1696
rect 623 1665 783 1672
rect 327 1662 783 1665
rect 817 1662 823 1696
rect 327 1627 823 1662
rect 327 1593 333 1627
rect 367 1608 589 1627
rect 367 1593 385 1608
tri 385 1593 400 1608 nw
tri 556 1593 571 1608 ne
rect 571 1593 589 1608
rect 623 1624 823 1627
rect 943 1689 1010 1708
tri 1010 1689 1029 1708 sw
rect 2289 1695 2524 1709
rect 3518 1877 3598 1881
rect 3518 1843 3558 1877
rect 3592 1843 3598 1877
rect 3518 1829 3598 1843
rect 3466 1817 3598 1829
rect 3518 1805 3598 1817
rect 3518 1771 3558 1805
rect 3592 1771 3598 1805
tri 3682 1891 3695 1904 sw
rect 3682 1882 3695 1891
tri 3695 1882 3704 1891 sw
tri 4374 1882 4383 1891 se
rect 4383 1885 4519 1891
rect 4383 1882 4467 1885
rect 3682 1879 4467 1882
rect 3682 1846 4389 1879
rect 3630 1845 4389 1846
rect 4423 1845 4467 1879
rect 3630 1836 4467 1845
rect 3630 1834 3699 1836
rect 3682 1813 3699 1834
tri 3699 1813 3722 1836 nw
tri 4355 1813 4378 1836 ne
rect 4378 1833 4467 1836
rect 4378 1819 4519 1833
rect 4378 1813 4467 1819
rect 3682 1807 3693 1813
tri 3693 1807 3699 1813 nw
tri 4378 1808 4383 1813 ne
rect 3682 1802 3688 1807
tri 3688 1802 3693 1807 nw
rect 4055 1802 4343 1808
tri 3682 1796 3688 1802 nw
rect 3630 1776 3682 1782
rect 3518 1765 3598 1771
rect 3466 1759 3598 1765
rect 4055 1768 4067 1802
rect 4101 1768 4139 1802
rect 4173 1768 4225 1802
rect 4259 1768 4297 1802
rect 4331 1768 4343 1802
rect 4055 1762 4343 1768
rect 4383 1807 4467 1813
rect 4383 1773 4389 1807
rect 4423 1773 4467 1807
rect 4383 1767 4467 1773
rect 4383 1761 4519 1767
rect 4803 1847 5082 1859
rect 4803 1813 5042 1847
rect 5076 1813 5082 1847
tri 4802 1761 4803 1762 se
rect 4803 1761 4862 1813
tri 4862 1779 4896 1813 nw
tri 5002 1779 5036 1813 ne
rect 5036 1775 5082 1813
rect 5540 1805 5851 2006
tri 4800 1759 4802 1761 se
rect 4802 1759 4862 1761
tri 4775 1734 4800 1759 se
rect 4800 1734 4862 1759
rect 3257 1719 3309 1725
rect 3639 1721 3685 1733
tri 3685 1721 3689 1725 sw
tri 3901 1721 3905 1725 se
rect 3905 1721 3951 1733
rect 943 1671 1029 1689
tri 1029 1671 1047 1689 sw
rect 2289 1683 2576 1695
rect 2289 1680 2524 1683
rect 2289 1671 2365 1680
rect 943 1664 1047 1671
tri 1047 1664 1054 1671 sw
rect 943 1658 2145 1664
rect 943 1654 2027 1658
tri 943 1624 973 1654 ne
rect 973 1624 2027 1654
rect 2061 1624 2099 1658
rect 2133 1624 2145 1658
rect 2289 1637 2295 1671
rect 2329 1655 2365 1671
tri 2365 1655 2390 1680 nw
tri 2490 1655 2515 1680 ne
rect 2515 1655 2524 1680
rect 2329 1649 2359 1655
tri 2359 1649 2365 1655 nw
tri 2515 1649 2521 1655 ne
rect 2521 1649 2524 1655
rect 2329 1637 2335 1649
rect 2289 1625 2335 1637
tri 2335 1625 2359 1649 nw
tri 2521 1646 2524 1649 ne
rect 2524 1625 2576 1631
rect 2887 1689 2933 1701
tri 2933 1689 2940 1696 sw
tri 3074 1689 3081 1696 se
rect 3081 1689 3127 1701
tri 3127 1689 3134 1696 sw
tri 3332 1689 3339 1696 se
rect 3339 1689 3385 1701
rect 2887 1655 2893 1689
rect 2927 1662 2940 1689
tri 2940 1662 2967 1689 sw
tri 3047 1662 3074 1689 se
rect 3074 1662 3087 1689
rect 2927 1655 3087 1662
rect 3121 1662 3134 1689
tri 3134 1662 3161 1689 sw
tri 3305 1662 3332 1689 se
rect 3332 1662 3345 1689
rect 3121 1655 3345 1662
rect 3379 1655 3385 1689
rect 623 1608 783 1624
rect 623 1593 638 1608
rect 327 1590 382 1593
tri 382 1590 385 1593 nw
tri 571 1590 574 1593 ne
rect 574 1590 638 1593
tri 638 1590 656 1608 nw
tri 751 1590 769 1608 ne
rect 769 1590 783 1608
rect 817 1590 823 1624
tri 973 1618 979 1624 ne
rect 979 1618 2145 1624
rect 327 1583 375 1590
tri 375 1583 382 1590 nw
tri 574 1583 581 1590 ne
rect 581 1583 631 1590
tri 631 1583 638 1590 nw
tri 769 1583 776 1590 ne
rect 776 1583 823 1590
rect 327 1581 373 1583
tri 373 1581 375 1583 nw
tri 581 1581 583 1583 ne
rect 583 1581 629 1583
tri 629 1581 631 1583 nw
tri 776 1582 777 1583 ne
rect 777 1578 823 1583
rect 2887 1617 3385 1655
rect 2887 1583 2893 1617
rect 2927 1598 3087 1617
rect 2927 1583 2945 1598
tri 2945 1583 2960 1598 nw
tri 3054 1583 3069 1598 ne
rect 3069 1583 3087 1598
rect 3121 1598 3345 1617
rect 3121 1583 3139 1598
tri 3139 1583 3154 1598 nw
tri 3312 1583 3327 1598 ne
rect 3327 1583 3345 1598
rect 3379 1583 3385 1617
rect 3639 1687 3645 1721
rect 3679 1691 3689 1721
tri 3689 1691 3719 1721 sw
tri 3871 1691 3901 1721 se
rect 3901 1691 3911 1721
rect 3679 1687 3911 1691
rect 3945 1687 3951 1721
rect 3639 1649 3951 1687
rect 4095 1682 4101 1734
rect 4153 1682 4165 1734
rect 4217 1728 4241 1734
tri 4241 1728 4247 1734 sw
tri 4769 1728 4775 1734 se
rect 4775 1728 4862 1734
rect 4217 1682 4862 1728
rect 4943 1762 4989 1774
rect 4943 1728 4949 1762
rect 4983 1728 4989 1762
rect 5036 1741 5042 1775
rect 5076 1741 5082 1775
rect 5036 1729 5082 1741
rect 4943 1690 4989 1728
tri 4935 1656 4943 1664 se
rect 4943 1656 4949 1690
rect 4983 1656 4989 1690
rect 7159 1677 7237 1745
tri 4934 1655 4935 1656 se
rect 4935 1655 4989 1656
rect 3639 1615 3645 1649
rect 3679 1645 3911 1649
rect 3679 1640 3714 1645
tri 3714 1640 3719 1645 nw
tri 3871 1640 3876 1645 ne
rect 3876 1640 3911 1645
rect 3679 1625 3699 1640
tri 3699 1625 3714 1640 nw
tri 3876 1625 3891 1640 ne
rect 3891 1625 3911 1640
rect 3679 1618 3692 1625
tri 3692 1618 3699 1625 nw
tri 3891 1618 3898 1625 ne
rect 3898 1618 3911 1625
rect 3679 1615 3689 1618
tri 3689 1615 3692 1618 nw
tri 3898 1615 3901 1618 ne
rect 3901 1615 3911 1618
rect 3945 1615 3951 1649
rect 3639 1603 3685 1615
tri 3685 1611 3689 1615 nw
tri 3901 1611 3905 1615 ne
rect 3905 1603 3951 1615
rect 3984 1649 4037 1655
rect 2887 1571 2933 1583
tri 2933 1571 2945 1583 nw
tri 3069 1571 3081 1583 ne
rect 3081 1571 3127 1583
tri 3127 1571 3139 1583 nw
tri 3327 1571 3339 1583 ne
rect 3339 1571 3385 1583
rect 4036 1597 4037 1649
tri 4925 1646 4934 1655 se
rect 4934 1646 4989 1655
tri 4919 1640 4925 1646 se
rect 4925 1640 4989 1646
rect 3984 1583 4037 1597
rect 3724 1534 3770 1546
rect 3724 1500 3730 1534
rect 3764 1500 3770 1534
rect 4036 1531 4037 1583
rect 3984 1525 4037 1531
rect 4200 1634 4252 1640
tri 4252 1630 4262 1640 sw
tri 4909 1630 4919 1640 se
rect 4919 1630 4989 1640
rect 4252 1625 4262 1630
tri 4262 1625 4267 1630 sw
rect 4252 1624 4267 1625
tri 4267 1624 4268 1625 sw
rect 4252 1582 4520 1624
rect 4200 1578 4520 1582
rect 4200 1570 4252 1578
tri 4252 1552 4278 1578 nw
tri 4440 1552 4466 1578 ne
rect 4466 1552 4520 1578
tri 4466 1550 4468 1552 ne
rect 4468 1550 4520 1552
rect 4200 1512 4252 1518
rect 4291 1544 4343 1550
tri 4468 1546 4472 1550 ne
rect 4472 1546 4520 1550
tri 4472 1544 4474 1546 ne
rect 3724 1499 3770 1500
tri 3770 1499 3779 1508 sw
tri 4282 1499 4291 1508 se
rect 410 1493 462 1499
rect 3724 1496 3779 1499
tri 3779 1496 3782 1499 sw
tri 4279 1496 4282 1499 se
rect 4282 1496 4291 1499
rect 201 1483 253 1489
rect 201 1417 253 1431
tri 462 1484 466 1488 sw
tri 1186 1484 1190 1488 se
rect 1190 1484 1236 1496
rect 462 1454 466 1484
tri 466 1454 496 1484 sw
tri 1156 1454 1186 1484 se
rect 1186 1454 1196 1484
rect 462 1450 1196 1454
rect 1230 1450 1236 1484
rect 462 1441 1236 1450
rect 410 1424 1236 1441
rect 2987 1484 3033 1496
rect 2987 1450 2993 1484
rect 3027 1450 3033 1484
tri 1656 1428 1667 1439 se
rect 462 1412 1236 1424
tri 1649 1421 1656 1428 se
rect 1656 1421 1667 1428
tri 1640 1412 1649 1421 se
rect 1649 1412 1667 1421
rect 462 1408 1196 1412
rect 462 1378 466 1408
tri 466 1378 496 1408 nw
tri 1156 1378 1186 1408 ne
rect 1186 1378 1196 1408
rect 1230 1378 1236 1412
tri 1606 1378 1640 1412 se
rect 1640 1378 1667 1412
tri 462 1374 466 1378 nw
tri 1186 1374 1190 1378 ne
rect 410 1366 462 1372
rect 1190 1366 1236 1378
tri 1594 1366 1606 1378 se
rect 1606 1366 1667 1378
rect 201 1359 253 1365
tri 1587 1359 1594 1366 se
rect 1594 1359 1667 1366
tri 1551 1323 1587 1359 se
rect 1587 1323 1667 1359
tri -185 1160 -154 1191 se
rect 107 1121 279 1323
rect 1173 1309 1667 1323
rect 2384 1428 2417 1439
tri 2417 1428 2428 1439 sw
rect 2384 1421 2428 1428
tri 2428 1421 2435 1428 sw
rect 2384 1418 2435 1421
tri 2435 1418 2438 1421 sw
rect 2384 1412 2438 1418
tri 2438 1412 2444 1418 sw
rect 2987 1412 3033 1450
rect 3724 1493 3782 1496
tri 3782 1493 3785 1496 sw
tri 4276 1493 4279 1496 se
rect 4279 1493 4291 1496
rect 3724 1474 3785 1493
tri 3785 1474 3804 1493 sw
tri 4257 1474 4276 1493 se
rect 4276 1492 4291 1493
rect 4276 1480 4343 1492
rect 4276 1474 4291 1480
rect 3724 1462 4291 1474
rect 3724 1428 3730 1462
rect 3764 1428 4291 1462
rect 3724 1422 4343 1428
rect 4474 1496 4520 1546
rect 4559 1618 4989 1630
tri 7077 1625 7098 1646 ne
rect 7098 1625 7332 1646
tri 7098 1618 7105 1625 ne
rect 7105 1618 7332 1625
rect 4559 1584 4565 1618
rect 4599 1584 4989 1618
tri 7105 1616 7107 1618 ne
rect 7107 1616 7332 1618
tri 7332 1616 7362 1646 nw
rect 4559 1578 4633 1584
tri 4633 1578 4639 1584 nw
rect 4559 1546 4605 1578
tri 4605 1550 4633 1578 nw
rect 4559 1512 4565 1546
rect 4599 1512 4605 1546
rect 7159 1541 7237 1609
rect 4559 1500 4605 1512
rect 4858 1527 4904 1539
tri 4520 1496 4522 1498 sw
tri 4856 1496 4858 1498 se
rect 4858 1496 4864 1527
rect 4474 1493 4522 1496
tri 4522 1493 4525 1496 sw
tri 4853 1493 4856 1496 se
rect 4856 1493 4864 1496
rect 4898 1493 4904 1527
rect 4474 1490 4525 1493
tri 4525 1490 4528 1493 sw
tri 4850 1490 4853 1493 se
rect 4853 1490 4904 1493
tri 5341 1490 5375 1524 sw
rect 4474 1464 4528 1490
tri 4528 1464 4554 1490 sw
tri 4824 1464 4850 1490 se
rect 4850 1464 4904 1490
rect 4474 1455 4904 1464
rect 3724 1421 3775 1422
tri 3775 1421 3776 1422 nw
rect 4474 1421 4864 1455
rect 4898 1421 4904 1455
rect 5798 1449 5833 1488
rect 6826 1452 6865 1496
rect 3724 1418 3772 1421
tri 3772 1418 3775 1421 nw
rect 4474 1418 4904 1421
rect 3724 1416 3770 1418
tri 3770 1416 3772 1418 nw
tri 4673 1416 4675 1418 ne
rect 4675 1416 4808 1418
tri 4675 1412 4679 1416 ne
rect 4679 1412 4808 1416
tri 4808 1412 4814 1418 nw
tri 4849 1412 4855 1418 ne
rect 4855 1412 4904 1418
rect 2384 1409 2444 1412
tri 2444 1409 2447 1412 sw
rect 2384 1378 2447 1409
tri 2447 1378 2478 1409 sw
rect 2987 1378 2993 1412
rect 3027 1378 3033 1412
tri 4855 1409 4858 1412 ne
rect 4858 1409 4904 1412
rect 7371 1409 7459 1454
rect 2384 1366 2478 1378
tri 2478 1366 2490 1378 sw
rect 2987 1366 3033 1378
rect 2384 1359 2490 1366
tri 2490 1359 2497 1366 sw
rect 2384 1323 2497 1359
tri 2497 1323 2533 1359 sw
rect 2384 1315 2533 1323
tri 2533 1315 2541 1323 sw
rect 2384 1309 4761 1315
rect 384 1169 695 1237
rect 1173 1177 4761 1309
rect 1148 1169 4761 1177
tri 5171 1169 5201 1199 sw
rect 353 1157 5167 1169
rect 5171 1168 5201 1169
tri 5201 1168 5202 1169 sw
rect 353 1123 441 1157
rect 475 1123 513 1157
rect 547 1123 585 1157
rect 619 1123 657 1157
rect 691 1123 729 1157
rect 763 1123 801 1157
rect 835 1123 873 1157
rect 907 1123 945 1157
rect 979 1123 1017 1157
rect 1051 1123 1089 1157
rect 1123 1123 1161 1157
rect 1195 1123 1233 1157
rect 1267 1123 1305 1157
rect 1339 1123 1377 1157
rect 1411 1123 1503 1157
rect 1537 1123 1575 1157
rect 1609 1123 1647 1157
rect 1681 1123 1719 1157
rect 1753 1123 1791 1157
rect 1825 1123 1863 1157
rect 1897 1123 1935 1157
rect 1969 1123 2007 1157
rect 2041 1123 2079 1157
rect 2113 1123 2151 1157
rect 2185 1123 2223 1157
rect 2257 1123 2295 1157
rect 2329 1123 2367 1157
rect 2401 1123 2439 1157
rect 2473 1123 2889 1157
rect 2923 1123 2961 1157
rect 2995 1123 3033 1157
rect 3067 1123 3105 1157
rect 3139 1123 3177 1157
rect 3211 1123 3249 1157
rect 3283 1123 3321 1157
rect 3355 1123 3393 1157
rect 3427 1123 3465 1157
rect 3499 1123 3537 1157
rect 3571 1123 3609 1157
rect 3643 1123 3681 1157
rect 3715 1123 3753 1157
rect 3787 1123 3825 1157
rect 3859 1123 3897 1157
rect 3931 1123 3969 1157
rect 4003 1123 4041 1157
rect 4075 1123 4113 1157
rect 4147 1123 4185 1157
rect 4219 1123 4257 1157
rect 4291 1123 4329 1157
rect 4363 1123 4401 1157
rect 4435 1123 4473 1157
rect 4507 1123 4545 1157
rect 4579 1123 4617 1157
rect 4651 1123 4689 1157
rect 4723 1123 4761 1157
rect 4795 1123 4833 1157
rect 4867 1123 4905 1157
rect 4939 1123 4977 1157
rect 5011 1123 5049 1157
rect 5083 1123 5121 1157
rect 5155 1123 5167 1157
rect 5483 1123 5522 1168
rect 279 957 306 1120
rect 353 1111 5167 1123
rect 384 1005 4761 1111
rect 441 965 4761 1005
rect 441 957 2497 965
tri 2497 957 2505 965 nw
tri 1521 937 1541 957 ne
rect 1541 944 2477 957
rect 1541 937 1634 944
tri 1541 925 1553 937 ne
rect 1553 925 1634 937
tri 1553 922 1556 925 ne
rect 1556 922 1634 925
tri 1556 908 1570 922 ne
rect 1570 908 1634 922
rect 679 896 810 908
rect 679 862 685 896
rect 719 862 810 896
tri 1570 891 1587 908 ne
rect 1587 891 1634 908
tri 1587 864 1614 891 ne
rect 1614 864 1634 891
rect 679 824 810 862
tri 1614 853 1625 864 ne
rect 1625 853 1634 864
tri 1625 844 1634 853 ne
rect 2384 937 2477 944
tri 2477 937 2497 957 nw
rect 2384 925 2465 937
tri 2465 925 2477 937 nw
tri 4842 925 4854 937 se
rect 4854 925 4900 937
rect 2384 922 2462 925
tri 2462 922 2465 925 nw
tri 4839 922 4842 925 se
rect 4842 922 4860 925
rect 2384 908 2448 922
tri 2448 908 2462 922 nw
tri 2599 908 2613 922 se
rect 2613 916 4860 922
rect 2613 908 3984 916
rect 2384 891 2431 908
tri 2431 891 2448 908 nw
tri 2582 891 2599 908 se
rect 2599 891 3984 908
rect 2384 864 2404 891
tri 2404 864 2431 891 nw
tri 2555 864 2582 891 se
rect 2582 879 3984 891
rect 2582 864 2613 879
tri 2613 864 2628 879 nw
tri 3950 864 3965 879 ne
rect 3965 864 3984 879
rect 4036 891 4860 916
rect 4894 891 4900 925
rect 4036 879 4900 891
rect 4036 864 4055 879
tri 4055 864 4070 879 nw
tri 4820 864 4835 879 ne
rect 4835 864 4900 879
rect 2384 853 2393 864
tri 2393 853 2404 864 nw
tri 2544 853 2555 864 se
rect 2555 853 2602 864
tri 2602 853 2613 864 nw
tri 3965 853 3976 864 ne
rect 3976 853 4044 864
tri 4044 853 4055 864 nw
tri 4835 853 4846 864 ne
rect 4846 853 4900 864
tri 2384 844 2393 853 nw
tri 2535 844 2544 853 se
rect 2544 844 2588 853
tri 2530 839 2535 844 se
rect 2535 839 2588 844
tri 2588 839 2602 853 nw
tri 3976 851 3978 853 ne
rect 3978 852 4036 853
rect 3978 851 3984 852
tri 2528 837 2530 839 se
rect 2530 837 2586 839
tri 2586 837 2588 839 nw
tri 2521 830 2528 837 se
rect 2528 830 2579 837
tri 2579 830 2586 837 nw
rect 2987 830 3033 842
rect 679 790 685 824
rect 719 790 810 824
tri 2500 809 2521 830 se
rect 2521 809 2558 830
tri 2558 809 2579 830 nw
tri 2497 806 2500 809 se
rect 2500 806 2555 809
tri 2555 806 2558 809 nw
tri 2488 797 2497 806 se
rect 2497 797 2545 806
rect 679 778 810 790
rect 24 763 70 765
rect 21 757 73 763
rect 21 693 73 705
rect 1719 742 1771 748
rect 1841 745 1847 797
rect 1899 745 1911 797
rect 1963 791 2111 797
tri 2487 796 2488 797 se
rect 2488 796 2545 797
tri 2545 796 2555 806 nw
rect 2987 796 2993 830
rect 3027 796 3033 830
rect 1963 757 1993 791
rect 2027 757 2065 791
rect 2099 757 2111 791
tri 2474 783 2487 796 se
rect 2487 783 2532 796
tri 2532 783 2545 796 nw
rect 1963 751 2111 757
rect 2344 776 2525 783
tri 2525 776 2532 783 nw
rect 2344 767 2516 776
tri 2516 767 2525 776 nw
rect 2344 765 2514 767
tri 2514 765 2516 767 nw
rect 2344 758 2507 765
tri 2507 758 2514 765 nw
rect 2987 758 3033 796
rect 2344 751 2500 758
tri 2500 751 2507 758 nw
rect 1963 745 1975 751
tri 1975 745 1981 751 nw
rect 2344 748 2497 751
tri 2497 748 2500 751 nw
rect 2344 741 2490 748
tri 2490 741 2497 748 nw
rect 21 635 73 641
rect 326 689 372 701
tri 372 689 384 701 sw
tri 571 689 583 701 se
rect 583 689 629 701
tri 629 689 641 701 sw
tri 765 689 777 701 se
rect 777 689 823 701
rect 326 655 332 689
rect 366 674 384 689
tri 384 674 399 689 sw
tri 556 674 571 689 se
rect 571 674 589 689
rect 366 655 589 674
rect 623 674 641 689
tri 641 674 656 689 sw
tri 750 674 765 689 se
rect 765 674 783 689
rect 623 655 783 674
rect 817 655 823 689
rect 326 617 823 655
rect 326 583 332 617
rect 366 610 589 617
rect 366 583 379 610
tri 379 583 406 610 nw
tri 549 583 576 610 ne
rect 576 583 589 610
rect 623 610 783 617
rect 623 583 636 610
tri 636 583 663 610 nw
tri 744 583 771 610 ne
rect 771 583 783 610
rect 817 583 823 617
rect 1069 688 1347 697
tri 1347 688 1356 697 sw
rect 2987 724 2993 758
rect 3027 724 3033 758
rect 2987 712 3033 724
rect 3255 839 3301 842
tri 3301 839 3304 842 sw
rect 3255 837 3304 839
tri 3304 837 3306 839 sw
rect 3639 837 3685 849
rect 3255 834 3306 837
tri 3306 834 3309 837 sw
rect 3255 830 3309 834
rect 3255 796 3261 830
rect 3295 822 3309 830
tri 3309 822 3321 834 sw
tri 3627 822 3639 834 se
rect 3639 822 3645 837
rect 3295 809 3321 822
tri 3321 809 3334 822 sw
tri 3614 809 3627 822 se
rect 3627 809 3645 822
rect 3295 806 3334 809
tri 3334 806 3337 809 sw
tri 3611 806 3614 809 se
rect 3614 806 3645 809
rect 3295 803 3337 806
tri 3337 803 3340 806 sw
tri 3608 803 3611 806 se
rect 3611 803 3645 806
rect 3679 803 3685 837
rect 3295 802 3340 803
tri 3340 802 3341 803 sw
tri 3607 802 3608 803 se
rect 3608 802 3685 803
rect 3295 801 3341 802
tri 3341 801 3342 802 sw
tri 3606 801 3607 802 se
rect 3607 801 3685 802
rect 3295 800 3342 801
tri 3342 800 3343 801 sw
tri 3605 800 3606 801 se
rect 3606 800 3685 801
rect 3295 796 3685 800
rect 3255 765 3685 796
rect 3255 758 3645 765
rect 3255 724 3261 758
rect 3295 754 3645 758
rect 3295 751 3332 754
tri 3332 751 3335 754 nw
tri 3605 751 3608 754 ne
rect 3608 751 3645 754
rect 3295 748 3329 751
tri 3329 748 3332 751 nw
tri 3608 748 3611 751 ne
rect 3611 748 3645 751
rect 3295 741 3322 748
tri 3322 741 3329 748 nw
tri 3611 741 3618 748 ne
rect 3618 741 3645 748
rect 3295 731 3312 741
tri 3312 731 3322 741 nw
tri 3618 731 3628 741 ne
rect 3628 731 3645 741
rect 3679 731 3685 765
rect 3295 724 3302 731
rect 3255 721 3302 724
tri 3302 721 3312 731 nw
tri 3628 721 3638 731 ne
rect 3638 721 3685 731
rect 3731 839 3777 851
tri 3978 845 3984 851 ne
rect 3731 805 3737 839
rect 3771 805 3777 839
rect 3731 783 3777 805
tri 3777 783 3795 801 sw
tri 4036 845 4044 853 nw
tri 4846 851 4848 853 ne
rect 4848 851 4860 853
rect 4115 839 4161 851
tri 4848 845 4854 851 ne
rect 4115 805 4121 839
rect 4155 805 4161 839
rect 4854 819 4860 851
rect 4894 819 4900 853
rect 5751 829 5918 985
rect 4854 807 4900 819
rect 4937 812 4989 822
rect 3984 794 4036 800
tri 4108 794 4115 801 se
rect 4115 794 4161 805
tri 4097 783 4108 794 se
rect 4108 783 4161 794
tri 4918 783 4937 802 se
rect 3731 781 3795 783
tri 3795 781 3797 783 sw
tri 4095 781 4097 783 se
rect 4097 781 4161 783
tri 4916 781 4918 783 se
rect 4918 781 4937 783
rect 3731 776 3797 781
tri 3797 776 3802 781 sw
tri 4090 776 4095 781 se
rect 4095 776 4161 781
rect 3731 767 3802 776
tri 3802 767 3811 776 sw
tri 4081 767 4090 776 se
rect 4090 767 4161 776
rect 3731 733 3737 767
rect 3771 766 3811 767
tri 3811 766 3812 767 sw
tri 4080 766 4081 767 se
rect 4081 766 4121 767
rect 3771 733 4121 766
rect 4155 733 4161 767
rect 3731 721 4161 733
rect 4210 776 4675 781
tri 4675 776 4680 781 sw
tri 4911 776 4916 781 se
rect 4916 776 4937 781
rect 4210 760 4937 776
tri 7318 767 7360 809 ne
rect 4210 748 4989 760
rect 4210 747 4937 748
rect 4210 741 4272 747
tri 4272 741 4278 747 nw
tri 4619 742 4624 747 ne
rect 4624 742 4937 747
tri 4909 741 4910 742 ne
rect 4910 741 4937 742
rect 4210 738 4269 741
tri 4269 738 4272 741 nw
tri 4910 738 4913 741 ne
rect 4913 738 4937 741
rect 4210 725 4256 738
tri 4256 725 4269 738 nw
tri 4913 725 4926 738 ne
rect 4926 725 4937 738
tri 4206 721 4210 725 se
rect 4210 721 4245 725
rect 3255 712 3301 721
tri 3301 720 3302 721 nw
tri 3638 720 3639 721 ne
rect 3639 719 3685 721
tri 4204 719 4206 721 se
rect 4206 719 4245 721
tri 4200 715 4204 719 se
rect 4204 715 4245 719
rect 1719 688 1728 690
rect 1762 688 1771 690
rect 1069 685 1356 688
rect 1069 651 1075 685
rect 1109 663 1356 685
tri 1356 663 1381 688 sw
rect 1719 678 1771 688
rect 1109 651 1381 663
rect 1069 650 1381 651
tri 1381 650 1394 663 sw
rect 1069 616 1394 650
tri 1394 616 1428 650 sw
rect 1719 616 1728 626
rect 1762 616 1771 626
rect 1069 613 1428 616
rect 326 579 375 583
tri 375 579 379 583 nw
tri 576 579 580 583 ne
rect 580 579 632 583
tri 632 579 636 583 nw
tri 771 579 775 583 ne
rect 775 579 823 583
rect 326 571 372 579
tri 372 576 375 579 nw
tri 580 576 583 579 ne
rect 583 571 629 579
tri 629 576 632 579 nw
tri 775 577 777 579 ne
rect 777 571 823 579
rect 980 574 1026 586
rect -65 539 -13 545
rect -65 473 -13 487
rect -65 415 -13 421
rect 110 539 162 545
rect 980 540 986 574
rect 1020 540 1026 574
rect 1069 579 1075 613
rect 1109 607 1428 613
tri 1428 607 1437 616 sw
rect 1109 604 1437 607
tri 1437 604 1440 607 sw
rect 1719 604 1771 616
rect 2887 707 2933 709
tri 2933 707 2935 709 sw
tri 3079 707 3081 709 se
rect 3081 707 3127 709
tri 3127 707 3129 709 sw
tri 3337 707 3339 709 se
rect 3339 707 3385 709
rect 2887 697 2935 707
tri 2935 697 2945 707 sw
tri 3069 697 3079 707 se
rect 3079 697 3129 707
tri 3129 697 3139 707 sw
tri 3327 697 3337 707 se
rect 3337 697 3385 707
rect 2887 663 2893 697
rect 2927 682 2945 697
tri 2945 682 2960 697 sw
tri 3054 682 3069 697 se
rect 3069 682 3087 697
rect 2927 663 3087 682
rect 3121 682 3139 697
tri 3139 682 3154 697 sw
tri 3312 682 3327 697 se
rect 3327 682 3345 697
rect 3121 663 3345 682
rect 3379 663 3385 697
rect 3474 663 3480 715
rect 3532 663 3544 715
rect 3596 714 3602 715
tri 3602 714 3603 715 sw
tri 4199 714 4200 715 se
rect 4200 714 4245 715
tri 4245 714 4256 725 nw
tri 4926 719 4932 725 ne
rect 4932 719 4937 725
rect 3596 707 3603 714
tri 3603 707 3610 714 sw
tri 4192 707 4199 714 se
rect 4199 707 4244 714
tri 4244 713 4245 714 nw
rect 3596 691 3610 707
tri 3610 691 3626 707 sw
tri 4176 691 4192 707 se
rect 4192 691 4244 707
rect 3596 663 4244 691
rect 4468 707 4514 719
tri 4932 714 4937 719 ne
rect 4468 673 4474 707
rect 4508 673 4514 707
rect 7360 714 7412 809
tri 7412 767 7454 809 nw
rect 4937 690 4989 696
tri 4462 663 4468 669 se
rect 4468 663 4514 673
rect 2887 625 3385 663
tri 4434 635 4462 663 se
rect 4462 635 4514 663
rect 1109 591 1440 604
tri 1440 591 1453 604 sw
rect 2887 591 2893 625
rect 2927 618 3087 625
rect 2927 604 2953 618
tri 2953 604 2967 618 nw
tri 3047 604 3061 618 ne
rect 3061 604 3087 618
rect 2927 591 2940 604
tri 2940 591 2953 604 nw
tri 3061 591 3074 604 ne
rect 3074 591 3087 604
rect 3121 618 3345 625
rect 3121 591 3134 618
tri 3134 591 3161 618 nw
tri 3305 591 3332 618 ne
rect 3332 591 3345 618
rect 3379 591 3385 625
rect 1109 579 1453 591
rect 1069 567 1453 579
tri 1453 567 1477 591 sw
rect 2887 579 2933 591
tri 2933 584 2940 591 nw
tri 3074 584 3081 591 ne
rect 3081 579 3127 591
tri 3127 584 3134 591 nw
tri 3332 584 3339 591 ne
rect 3339 579 3385 591
rect 3425 601 4474 635
rect 4508 601 4514 635
rect 3425 574 3466 601
tri 3466 574 3493 601 nw
tri 4456 589 4468 601 ne
rect 4468 589 4514 601
tri 1293 562 1298 567 ne
rect 1298 562 1477 567
tri 1477 562 1482 567 sw
tri 1298 559 1301 562 ne
rect 1301 559 1482 562
tri 1482 559 1485 562 sw
tri 1301 555 1305 559 ne
rect 1305 555 1485 559
tri 1485 555 1489 559 sw
tri 1305 553 1307 555 ne
rect 1307 553 1489 555
tri 1489 553 1491 555 sw
rect 110 473 162 487
rect 110 415 162 421
rect 415 526 461 538
rect 415 492 421 526
rect 455 521 461 526
tri 461 521 478 538 sw
tri 963 521 980 538 se
rect 980 521 1026 540
tri 1307 521 1339 553 ne
rect 1339 547 1520 553
rect 1339 521 1468 547
rect 455 504 478 521
tri 478 504 495 521 sw
tri 946 504 963 521 se
rect 963 504 1026 521
rect 455 502 1026 504
rect 455 492 986 502
rect 415 470 986 492
rect 415 468 489 470
tri 489 468 491 470 nw
tri 966 468 968 470 ne
rect 968 468 986 470
rect 1020 468 1026 502
tri 1339 490 1370 521 ne
rect 1370 495 1468 521
tri 3400 521 3425 546 se
rect 3425 521 3459 574
tri 3459 567 3466 574 nw
tri 3391 512 3400 521 se
rect 3400 512 3459 521
rect 1370 490 1520 495
tri 1370 487 1373 490 ne
rect 1373 487 1520 490
tri 1373 483 1377 487 ne
rect 1377 483 1520 487
rect 415 456 477 468
tri 477 456 489 468 nw
tri 968 456 980 468 ne
rect 980 456 1026 468
tri 1377 456 1404 483 ne
rect 1404 481 1520 483
rect 1404 456 1468 481
rect 415 454 470 456
rect 415 420 421 454
rect 455 449 470 454
tri 470 449 477 456 nw
tri 1404 449 1411 456 ne
rect 1411 449 1468 456
rect 455 420 461 449
tri 461 440 470 449 nw
tri 1411 440 1420 449 ne
rect 1420 440 1468 449
tri 1420 423 1437 440 ne
rect 1437 429 1468 440
rect 3257 460 3263 512
rect 3315 460 3327 512
rect 3379 460 3459 512
rect 3550 561 3602 567
rect 3550 494 3602 509
rect 3550 436 3602 442
rect 4027 561 4079 567
rect 4027 494 4079 509
rect 4027 436 4079 442
rect 4200 561 4252 567
rect 4200 494 4252 509
rect 4200 436 4252 442
rect 4383 565 4435 571
rect 4383 498 4435 513
rect 4383 440 4435 446
rect 4552 565 4604 571
rect 4552 498 4604 513
rect 5024 568 5076 574
rect 5024 504 5076 516
rect 5024 446 5076 452
rect 4552 440 4604 446
rect 5027 444 5073 446
rect 1437 423 1520 429
rect 415 408 461 420
tri 2776 337 2785 346 se
rect 2785 345 5202 346
rect 2785 337 3730 345
rect 929 163 931 337
tri 1250 310 1277 337 sw
tri 2761 322 2776 337 se
rect 2776 322 3730 337
tri 2488 316 2494 322 se
rect 2494 316 2518 322
rect 2211 310 2518 316
rect 1250 306 1277 310
tri 1277 306 1281 310 sw
rect 1235 163 1634 306
rect 2211 276 2223 310
rect 2257 276 2295 310
rect 2329 276 2518 310
tri 1634 242 1663 271 sw
rect 2211 270 2518 276
rect 2570 270 2582 322
rect 2634 270 2640 322
tri 2709 270 2761 322 se
rect 2761 293 3730 322
rect 3782 293 3808 345
rect 3860 293 3887 345
rect 3939 293 5202 345
rect 2761 270 5202 293
tri 2681 242 2709 270 se
rect 2709 266 5202 270
rect 2709 242 3730 266
rect 317 151 1634 163
rect 317 122 337 151
tri 300 117 305 122 ne
rect 305 117 337 122
rect 371 117 409 151
rect 443 117 481 151
rect 515 117 553 151
rect 587 117 625 151
rect 659 117 697 151
rect 731 117 769 151
rect 803 117 841 151
rect 875 117 913 151
rect 947 117 985 151
rect 1019 117 1057 151
rect 1091 117 1129 151
rect 1163 117 1201 151
rect 1235 117 1634 151
tri 305 105 317 117 ne
rect 317 112 1634 117
rect 2384 214 3730 242
rect 3782 214 3808 266
rect 3860 214 3887 266
rect 3939 214 5202 266
rect 2384 187 5202 214
rect 2384 176 3730 187
rect 3782 176 3808 187
rect 2384 142 2817 176
rect 2851 142 2889 176
rect 2923 142 2961 176
rect 2995 142 3033 176
rect 3067 142 3105 176
rect 3139 142 3177 176
rect 3211 142 3249 176
rect 3283 142 3321 176
rect 3355 142 3393 176
rect 3427 142 3465 176
rect 3499 142 3537 176
rect 3571 142 3609 176
rect 3643 142 3681 176
rect 3715 142 3730 176
rect 3787 142 3808 176
rect 2384 135 3730 142
rect 3782 135 3808 142
rect 3860 135 3887 187
rect 3939 176 5202 187
rect 3939 142 3969 176
rect 4003 142 4041 176
rect 4075 142 4113 176
rect 4147 142 4185 176
rect 4219 142 4257 176
rect 4291 142 4329 176
rect 4363 142 4401 176
rect 4435 142 4473 176
rect 4507 142 4545 176
rect 4579 142 4617 176
rect 4651 142 4689 176
rect 4723 142 4761 176
rect 4795 142 4833 176
rect 4867 142 4905 176
rect 4939 142 4977 176
rect 5011 142 5049 176
rect 5083 142 5121 176
rect 5155 142 5202 176
rect 3939 135 5202 142
rect 2384 130 5202 135
rect 2384 112 2805 130
tri 2805 112 2823 130 nw
rect 317 105 1247 112
tri 1247 105 1254 112 nw
<< via1 >>
rect 2706 2797 2758 2849
rect 2777 2797 2829 2849
rect 3932 2797 3984 2849
rect 3996 2797 4048 2849
rect 31 2705 83 2757
rect 95 2705 147 2757
rect 2486 2705 2538 2757
rect 2550 2705 2602 2757
rect 129 2613 181 2665
rect 193 2613 245 2665
rect 2064 2613 2116 2665
rect 2128 2613 2180 2665
rect 3443 2613 3495 2665
rect 3507 2613 3559 2665
rect 4482 2613 4534 2665
rect 4546 2613 4598 2665
rect -133 2521 -81 2573
rect -69 2521 -17 2573
rect 1681 2521 1733 2573
rect 1745 2521 1797 2573
rect 4313 2521 4365 2573
rect 4377 2521 4429 2573
rect 1413 2429 1465 2481
rect 1477 2429 1529 2481
rect 4867 2429 4919 2481
rect 4931 2429 4983 2481
rect 1873 2337 1925 2389
rect 1937 2337 1989 2389
rect 4221 2337 4273 2389
rect 4285 2337 4337 2389
rect -63 1850 -11 1856
rect -63 1816 -54 1850
rect -54 1816 -20 1850
rect -20 1816 -11 1850
rect -63 1804 -11 1816
rect -63 1778 -11 1792
rect -63 1744 -54 1778
rect -54 1744 -20 1778
rect -20 1744 -11 1778
rect -63 1740 -11 1744
rect 123 1850 175 1856
rect 123 1816 132 1850
rect 132 1816 166 1850
rect 166 1816 175 1850
rect 123 1804 175 1816
rect 123 1778 175 1792
rect 123 1744 132 1778
rect 132 1744 166 1778
rect 166 1744 175 1778
rect 123 1740 175 1744
rect 3257 1842 3309 1848
rect 1585 1781 1637 1833
rect 1585 1717 1637 1769
rect 3257 1808 3267 1842
rect 3267 1808 3301 1842
rect 3301 1808 3309 1842
rect 3257 1796 3309 1808
rect 3257 1770 3309 1777
rect 2048 1712 2100 1764
rect 2112 1712 2164 1764
rect 2524 1695 2576 1747
rect 3257 1736 3267 1770
rect 3267 1736 3301 1770
rect 3301 1736 3309 1770
rect 3466 1829 3518 1881
rect 3466 1765 3518 1817
rect 3630 1846 3682 1898
rect 3630 1782 3682 1834
rect 4467 1833 4519 1885
rect 4467 1767 4519 1819
rect 3257 1725 3309 1736
rect 2524 1631 2576 1683
rect 4101 1682 4153 1734
rect 4165 1682 4217 1734
rect 3984 1643 4036 1649
rect 3984 1609 3997 1643
rect 3997 1609 4031 1643
rect 4031 1609 4036 1643
rect 3984 1597 4036 1609
rect 3984 1571 4036 1583
rect 3984 1537 3997 1571
rect 3997 1537 4031 1571
rect 4031 1537 4036 1571
rect 3984 1531 4036 1537
rect 4200 1582 4252 1634
rect 4200 1518 4252 1570
rect 201 1477 253 1483
rect 201 1443 210 1477
rect 210 1443 244 1477
rect 244 1443 253 1477
rect 201 1431 253 1443
rect 201 1405 253 1417
rect 201 1371 210 1405
rect 210 1371 244 1405
rect 244 1371 253 1405
rect 201 1365 253 1371
rect 410 1484 462 1493
rect 410 1450 421 1484
rect 421 1450 455 1484
rect 455 1450 462 1484
rect 410 1441 462 1450
rect 410 1412 462 1424
rect 410 1378 421 1412
rect 421 1378 455 1412
rect 455 1378 462 1412
rect 410 1372 462 1378
rect 4291 1492 4343 1544
rect 4291 1428 4343 1480
rect 3984 864 4036 916
rect 21 753 73 757
rect 21 719 30 753
rect 30 719 64 753
rect 64 719 73 753
rect 21 705 73 719
rect 1847 745 1899 797
rect 1911 745 1963 797
rect 1719 722 1771 742
rect 21 681 73 693
rect 21 647 30 681
rect 30 647 64 681
rect 64 647 73 681
rect 21 641 73 647
rect 1719 690 1728 722
rect 1728 690 1762 722
rect 1762 690 1771 722
rect 3984 800 4036 852
rect 4937 810 4989 812
rect 4937 776 4949 810
rect 4949 776 4983 810
rect 4983 776 4989 810
rect 4937 760 4989 776
rect 4937 738 4989 748
rect 1719 650 1771 678
rect 1719 626 1728 650
rect 1728 626 1762 650
rect 1762 626 1771 650
rect -65 533 -13 539
rect -65 499 -56 533
rect -56 499 -22 533
rect -22 499 -13 533
rect -65 487 -13 499
rect -65 461 -13 473
rect -65 427 -56 461
rect -56 427 -22 461
rect -22 427 -13 461
rect -65 421 -13 427
rect 110 533 162 539
rect 3480 663 3532 715
rect 3544 663 3596 715
rect 4937 704 4949 738
rect 4949 704 4983 738
rect 4983 704 4989 738
rect 4937 696 4989 704
rect 110 499 119 533
rect 119 499 153 533
rect 153 499 162 533
rect 110 487 162 499
rect 110 461 162 473
rect 110 427 119 461
rect 119 427 153 461
rect 153 427 162 461
rect 110 421 162 427
rect 1468 495 1520 547
rect 1468 429 1520 481
rect 3263 460 3315 512
rect 3327 460 3379 512
rect 3550 555 3602 561
rect 3550 521 3559 555
rect 3559 521 3593 555
rect 3593 521 3602 555
rect 3550 509 3602 521
rect 3550 483 3602 494
rect 3550 449 3559 483
rect 3559 449 3593 483
rect 3593 449 3602 483
rect 3550 442 3602 449
rect 4027 555 4079 561
rect 4027 521 4036 555
rect 4036 521 4070 555
rect 4070 521 4079 555
rect 4027 509 4079 521
rect 4027 483 4079 494
rect 4027 449 4036 483
rect 4036 449 4070 483
rect 4070 449 4079 483
rect 4027 442 4079 449
rect 4200 555 4252 561
rect 4200 521 4209 555
rect 4209 521 4243 555
rect 4243 521 4252 555
rect 4200 509 4252 521
rect 4200 483 4252 494
rect 4200 449 4209 483
rect 4209 449 4243 483
rect 4243 449 4252 483
rect 4200 442 4252 449
rect 4383 559 4435 565
rect 4383 525 4392 559
rect 4392 525 4426 559
rect 4426 525 4435 559
rect 4383 513 4435 525
rect 4383 487 4435 498
rect 4383 453 4392 487
rect 4392 453 4426 487
rect 4426 453 4435 487
rect 4383 446 4435 453
rect 4552 559 4604 565
rect 4552 525 4561 559
rect 4561 525 4595 559
rect 4595 525 4604 559
rect 4552 513 4604 525
rect 4552 487 4604 498
rect 4552 453 4561 487
rect 4561 453 4595 487
rect 4595 453 4604 487
rect 4552 446 4604 453
rect 5024 562 5076 568
rect 5024 528 5033 562
rect 5033 528 5067 562
rect 5067 528 5076 562
rect 5024 516 5076 528
rect 5024 490 5076 504
rect 5024 456 5033 490
rect 5033 456 5067 490
rect 5067 456 5076 490
rect 5024 452 5076 456
rect 2518 270 2570 322
rect 2582 270 2634 322
rect 3730 293 3782 345
rect 3808 293 3860 345
rect 3887 293 3939 345
rect 3730 214 3782 266
rect 3808 214 3860 266
rect 3887 214 3939 266
rect 3730 176 3782 187
rect 3808 176 3860 187
rect 3730 142 3753 176
rect 3753 142 3782 176
rect 3808 142 3825 176
rect 3825 142 3859 176
rect 3859 142 3860 176
rect 3730 135 3782 142
rect 3808 135 3860 142
rect 3887 176 3939 187
rect 3887 142 3897 176
rect 3897 142 3931 176
rect 3931 142 3939 176
rect 3887 135 3939 142
<< metal2 >>
tri 1744 2797 1796 2849 se
rect 1796 2797 2706 2849
rect 2758 2797 2777 2849
rect 2829 2797 2835 2849
rect 3926 2797 3932 2849
rect 3984 2797 3996 2849
rect 4048 2797 4054 2849
tri 1722 2775 1744 2797 se
rect 1744 2775 1796 2797
tri 1796 2775 1818 2797 nw
tri 3946 2775 3968 2797 ne
rect 3968 2775 4032 2797
tri 4032 2775 4054 2797 nw
tri 1710 2763 1722 2775 se
rect 1722 2763 1784 2775
tri 1784 2763 1796 2775 nw
tri 3968 2763 3980 2775 ne
tri 1704 2757 1710 2763 se
rect 1710 2757 1778 2763
tri 1778 2757 1784 2763 nw
rect 25 2705 31 2757
rect 83 2705 95 2757
rect 147 2705 153 2757
tri 1652 2705 1704 2757 se
rect 1704 2705 1726 2757
tri 1726 2705 1778 2757 nw
rect 2480 2705 2486 2757
rect 2538 2705 2550 2757
rect 2602 2705 2608 2757
rect 25 2701 107 2705
tri 107 2701 111 2705 nw
tri 1648 2701 1652 2705 se
rect 1652 2701 1722 2705
tri 1722 2701 1726 2705 nw
tri 2490 2701 2494 2705 ne
rect 2494 2701 2576 2705
rect -139 2521 -133 2573
rect -81 2521 -69 2573
rect -17 2521 -11 2573
tri -97 2487 -63 2521 ne
rect -63 1856 -11 2521
rect -63 1792 -11 1804
rect -63 1734 -11 1740
tri 9 1631 25 1647 se
rect 25 1631 77 2701
tri 77 2671 107 2701 nw
tri 1618 2671 1648 2701 se
rect 1648 2671 1686 2701
tri 1612 2665 1618 2671 se
rect 1618 2665 1686 2671
tri 1686 2665 1722 2701 nw
tri 2494 2671 2524 2701 ne
rect 123 2613 129 2665
rect 181 2613 193 2665
rect 245 2613 251 2665
tri 1585 2638 1612 2665 se
rect 1612 2638 1659 2665
tri 1659 2638 1686 2665 nw
rect 123 1856 175 2613
tri 175 2579 209 2613 nw
rect 1407 2429 1413 2481
rect 1465 2429 1477 2481
rect 1529 2429 1535 2481
tri 1434 2395 1468 2429 ne
rect 123 1792 175 1804
rect 123 1734 175 1740
tri 3 1625 9 1631 se
rect 9 1625 77 1631
tri -13 1609 3 1625 se
rect 3 1609 61 1625
tri 61 1609 77 1625 nw
tri -25 1597 -13 1609 se
rect -13 1597 49 1609
tri 49 1597 61 1609 nw
tri -39 1583 -25 1597 se
rect -25 1583 35 1597
tri 35 1583 49 1597 nw
tri -65 1557 -39 1583 se
rect -39 1557 -13 1583
rect -65 539 -13 1557
tri -13 1535 35 1583 nw
rect 410 1493 462 1499
rect 201 1483 253 1489
rect 201 1417 253 1431
rect 410 1424 462 1441
rect 410 1366 462 1372
tri 179 1154 201 1176 se
rect 201 1154 253 1365
tri 162 1137 179 1154 se
rect 179 1137 236 1154
tri 236 1137 253 1154 nw
tri 110 1085 162 1137 se
rect 21 757 73 763
rect 21 693 73 705
rect 21 635 73 641
rect -65 473 -13 487
rect -65 415 -13 421
rect 110 539 162 1085
tri 162 1063 236 1137 nw
rect 110 473 162 487
rect 1468 547 1520 2429
tri 1520 2414 1535 2429 nw
rect 1585 1833 1637 2638
tri 1637 2616 1659 2638 nw
rect 2058 2613 2064 2665
rect 2116 2613 2128 2665
rect 2180 2613 2186 2665
tri 2068 2579 2102 2613 ne
rect 1675 2521 1681 2573
rect 1733 2521 1745 2573
rect 1797 2521 1803 2573
tri 1685 2489 1717 2521 ne
rect 1717 2489 1771 2521
tri 1771 2489 1803 2521 nw
tri 1717 2487 1719 2489 ne
rect 1585 1769 1637 1781
rect 1585 1711 1637 1717
rect 1719 742 1771 2489
rect 1867 2337 1873 2389
rect 1925 2337 1937 2389
rect 1989 2337 1995 2389
tri 1867 2333 1871 2337 ne
tri 1844 800 1871 827 se
rect 1871 800 1917 2337
tri 1917 2303 1951 2337 nw
tri 2100 1796 2102 1798 se
rect 2102 1796 2148 2613
tri 2148 2581 2180 2613 nw
tri 2514 2429 2524 2439 se
rect 2524 2429 2576 2701
tri 2576 2673 2608 2705 nw
rect 3437 2613 3443 2665
rect 3495 2613 3507 2665
rect 3559 2613 3565 2665
tri 3437 2584 3466 2613 ne
tri 2490 2405 2514 2429 se
rect 2514 2405 2576 2429
rect 2434 2353 2576 2405
rect 2434 2337 2504 2353
tri 2504 2337 2520 2353 nw
rect 2434 2179 2486 2337
tri 2486 2319 2504 2337 nw
tri 2486 2179 2520 2213 sw
rect 2434 2127 2576 2179
tri 2490 2093 2524 2127 ne
tri 2081 1777 2100 1796 se
rect 2100 1777 2148 1796
tri 2148 1777 2157 1786 sw
tri 2068 1764 2081 1777 se
rect 2081 1764 2157 1777
tri 2157 1764 2170 1777 sw
rect 2042 1712 2048 1764
rect 2100 1712 2112 1764
rect 2164 1712 2170 1764
rect 2524 1747 2576 2127
rect 3466 1881 3518 2613
tri 3518 2579 3552 2613 nw
rect 3980 2521 4032 2775
rect 4476 2613 4482 2665
rect 4534 2613 4546 2665
rect 4598 2613 4604 2665
tri 4518 2579 4552 2613 ne
tri 4032 2521 4036 2525 sw
rect 4307 2521 4313 2573
rect 4365 2521 4377 2573
rect 4429 2521 4435 2573
rect 3980 2491 4036 2521
tri 4036 2491 4066 2521 sw
tri 4349 2491 4379 2521 ne
rect 4379 2491 4435 2521
rect 3980 2439 4143 2491
tri 4379 2487 4383 2491 ne
tri 4057 2429 4067 2439 ne
rect 4067 2429 4143 2439
tri 4067 2405 4091 2429 ne
rect 2524 1683 2576 1695
tri 1917 800 1948 831 sw
tri 1841 797 1844 800 se
rect 1844 797 1948 800
tri 1948 797 1951 800 sw
rect 1841 745 1847 797
rect 1899 745 1911 797
rect 1963 745 1969 797
rect 1719 678 1771 690
rect 1719 620 1771 626
rect 1468 481 1520 495
rect 1468 423 1520 429
rect 110 415 162 421
rect 2524 345 2576 1631
rect 3257 1848 3309 1854
rect 3257 1777 3309 1796
rect 3466 1817 3518 1829
rect 3466 1759 3518 1765
rect 3630 1898 3682 1904
rect 3630 1834 3682 1846
rect 3257 512 3309 1725
rect 3474 663 3480 715
rect 3532 663 3544 715
rect 3596 663 3602 715
tri 3562 568 3630 636 se
rect 3630 568 3682 1782
rect 4091 1767 4143 2429
rect 4215 2337 4221 2389
rect 4273 2337 4285 2389
rect 4337 2337 4343 2389
tri 4257 2303 4291 2337 ne
tri 4143 1767 4144 1768 sw
rect 4091 1734 4144 1767
tri 4144 1734 4177 1767 sw
rect 4091 1682 4101 1734
rect 4153 1682 4165 1734
rect 4217 1682 4223 1734
rect 3984 1649 4036 1655
rect 3984 1583 4036 1597
rect 3984 916 4036 1531
rect 3984 852 4036 864
rect 3984 794 4036 800
tri 3561 567 3562 568 se
rect 3562 567 3682 568
rect 3550 561 3682 567
tri 3309 512 3343 546 sw
rect 3257 460 3263 512
rect 3315 460 3327 512
rect 3379 460 3385 512
rect 3602 528 3682 561
tri 4027 614 4091 678 se
rect 4091 656 4143 1682
tri 4143 1648 4177 1682 nw
rect 4091 614 4101 656
tri 4101 614 4143 656 nw
rect 4200 1634 4252 1640
rect 4200 1570 4252 1582
rect 4027 561 4079 614
tri 4079 592 4101 614 nw
rect 3602 509 3639 528
tri 3639 509 3658 528 nw
rect 3550 504 3634 509
tri 3634 504 3639 509 nw
rect 3550 498 3628 504
tri 3628 498 3634 504 nw
rect 3550 494 3624 498
tri 3624 494 3628 498 nw
rect 4027 494 4079 509
tri 3602 472 3624 494 nw
tri 2576 345 2587 356 sw
tri 2512 322 2524 334 se
rect 2524 322 2587 345
tri 2587 322 2610 345 sw
rect 2512 270 2518 322
rect 2570 270 2582 322
rect 2634 270 2640 322
rect 3550 285 3602 442
rect 3724 345 3945 346
rect 3724 293 3730 345
rect 3782 293 3808 345
rect 3860 293 3887 345
rect 3939 293 3945 345
rect 3724 266 3945 293
rect 4027 269 4079 442
rect 4200 561 4252 1518
rect 4291 1544 4343 2337
rect 4291 1480 4343 1492
rect 4291 1422 4343 1428
rect 4200 494 4252 509
rect 4200 285 4252 442
rect 4383 565 4435 2491
rect 4383 498 4435 513
rect 4383 440 4435 446
rect 4467 1885 4519 1891
rect 4467 1819 4519 1833
rect 4467 305 4519 1767
rect 4552 565 4604 2613
rect 4861 2429 4867 2481
rect 4919 2429 4931 2481
rect 4983 2429 4989 2481
tri 4903 2395 4937 2429 ne
rect 4937 812 4989 2429
rect 4937 748 4989 760
rect 4937 690 4989 696
rect 4552 498 4604 513
rect 4552 440 4604 446
rect 5024 568 5076 587
rect 5024 504 5076 516
rect 5024 412 5076 452
rect 3724 214 3730 266
rect 3782 214 3808 266
rect 3860 214 3887 266
rect 3939 214 3945 266
rect 3724 187 3945 214
rect 3724 135 3730 187
rect 3782 135 3808 187
rect 3860 135 3887 187
rect 3939 135 3945 187
rect 3724 134 3945 135
use sky130_fd_io__com_ctl_ls_octl  sky130_fd_io__com_ctl_ls_octl_0
timestamp 1619729480
transform 1 0 5445 0 -1 2130
box -71 10 2077 2019
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1619729480
transform 1 0 3095 0 -1 2174
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1619729480
transform 1 0 3095 0 1 106
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_2
timestamp 1619729480
transform -1 0 618 0 1 98
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_3
timestamp 1619729480
transform -1 0 1270 0 1 98
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_4
timestamp 1619729480
transform -1 0 618 0 -1 2182
box -46 24 399 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1619729480
transform 1 0 3747 0 -1 2174
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_1
timestamp 1619729480
transform -1 0 3929 0 -1 2174
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_2
timestamp 1619729480
transform -1 0 4757 0 -1 2174
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_3
timestamp 1619729480
transform 1 0 4699 0 1 106
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_4
timestamp 1619729480
transform -1 0 4405 0 1 106
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_5
timestamp 1619729480
transform 1 0 3395 0 1 106
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_6
timestamp 1619729480
transform 1 0 4223 0 1 106
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_7
timestamp 1619729480
transform -1 0 318 0 1 98
box -42 24 569 1116
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_0
timestamp 1619729480
transform 1 0 2743 0 -1 2174
box 0 24 534 1116
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_1
timestamp 1619729480
transform -1 0 3277 0 1 106
box 0 24 534 1116
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_2
timestamp 1619729480
transform -1 0 970 0 -1 2182
box 0 24 534 1116
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_3
timestamp 1619729480
transform -1 0 970 0 1 98
box 0 24 534 1116
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1619729480
transform 1 0 4699 0 -1 2174
box 0 24 534 1116
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_1
timestamp 1619729480
transform 1 0 788 0 -1 2182
box 0 24 534 1116
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_2
timestamp 1619729480
transform 1 0 -216 0 -1 2182
box 0 24 534 1116
use sky130_fd_io__hvsbt_xor  sky130_fd_io__hvsbt_xor_0
timestamp 1619729480
transform -1 0 2723 0 1 -63
box 95 75 1333 1135
use sky130_fd_io__hvsbt_xor  sky130_fd_io__hvsbt_xor_1
timestamp 1619729480
transform -1 0 2756 0 -1 2346
box 95 75 1333 1135
use sky130_fd_io__hvsbt_inv_x1_i2c_fix  sky130_fd_io__hvsbt_inv_x1_i2c_fix_0
timestamp 1619729480
transform 1 0 2032 0 -1 3724
box -1 41 358 1116
<< labels >>
flabel metal2 s 27 664 64 728 3 FreeSans 520 0 0 0 PDEN_H_N[2]
flabel metal2 s 5032 478 5063 543 3 FreeSans 520 0 0 0 VREG_EN_H_N
flabel metal2 s 416 1379 454 1471 3 FreeSans 520 0 0 0 PUEN_0_H
flabel metal2 s 3554 290 3598 339 3 FreeSans 520 90 0 0 DM_H_N[0]
flabel metal2 s 4209 296 4244 341 3 FreeSans 520 90 0 0 DM_H_N[2]
flabel metal2 s 3989 891 4020 985 3 FreeSans 520 180 0 0 PUEN_2OR1_H
flabel metal2 s 4385 471 4434 524 3 FreeSans 520 90 0 0 DM_H[1]
flabel metal2 s 4553 463 4602 526 3 FreeSans 520 90 0 0 DM_H[0]
flabel metal2 s 2538 336 2564 385 3 FreeSans 520 90 0 0 DM_H[2]
flabel metal2 s 4036 297 4070 346 3 FreeSans 520 90 0 0 DM_H_N[1]
flabel metal2 s 3576 314 3576 314 3 FreeSans 520 90 0 0 DM_H_N[0]
flabel metal2 s 4004 938 4004 938 3 FreeSans 520 180 0 0 PUEN_2OR1_H
flabel metal2 s 4227 318 4227 318 3 FreeSans 520 90 0 0 DM_H_N[2]
flabel comment s 4058 183 4058 183 0 FreeSans 440 90 0 0 DM_H_N[1]
flabel comment s 4586 866 4586 866 0 FreeSans 440 270 0 0 DM_H[0]
flabel comment s 4408 849 4408 849 0 FreeSans 440 270 0 0 DM_H[1]
flabel comment s 5067 1248 5067 1248 0 FreeSans 440 90 0 0 DM_H[2]
flabel comment s 4234 179 4234 179 0 FreeSans 440 90 0 0 DM_H_N[2]
flabel comment s 3582 245 3582 245 0 FreeSans 440 270 0 0 DM_H_N[0]
flabel metal1 s 682 1761 722 1838 3 FreeSans 520 0 0 0 PUEN_H[0]
flabel metal1 s 5751 829 5918 985 3 FreeSans 520 180 0 0 VGND
flabel metal1 s 5540 1805 5851 2006 3 FreeSans 520 180 0 0 VCC_IO
flabel metal1 s 682 793 722 870 3 FreeSans 520 0 0 0 PUEN_H[1]
flabel metal1 s 7159 1677 7237 1745 3 FreeSans 520 0 0 0 VPWR
flabel metal1 s 5798 1449 5833 1488 3 FreeSans 520 0 0 0 SLOW_H
flabel metal1 s 6826 1452 6865 1496 3 FreeSans 520 0 0 0 HLD_I_H_N
flabel metal1 s 7159 1541 7237 1609 3 FreeSans 520 0 0 0 VPWR
flabel metal1 s 7371 1409 7459 1454 3 FreeSans 520 0 0 0 SLOW
flabel metal1 s 2192 3308 2231 3357 3 FreeSans 520 0 0 0 OD_H
flabel metal1 s 5483 1123 5522 1168 3 FreeSans 520 0 0 0 SLOW_H_N
flabel metal1 s 384 1005 695 1237 3 FreeSans 520 180 0 0 VCC_IO
flabel metal1 s 358 2015 525 2171 3 FreeSans 520 180 0 0 VGND
flabel metal1 s 2994 770 3024 830 3 FreeSans 520 180 0 0 PDEN_H_N[1]
flabel metal1 s 2992 1405 3026 1469 3 FreeSans 520 180 0 0 PDEN_H_N[0]
flabel metal1 s 2852 152 3019 322 3 FreeSans 520 180 0 0 VGND
flabel metal1 s 2851 1028 3162 1260 3 FreeSans 520 180 0 0 VCC_IO
flabel metal1 s 2852 2117 3019 2273 3 FreeSans 520 180 0 0 VGND
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 36668874
string GDS_START 36596094
<< end >>
