magic
tech sky130A
magscale 1 2
timestamp 1619729485
<< metal4 >>
rect 0 35957 287 40800
rect 0 14807 529 19800
rect 0 13617 296 14507
rect 0 12447 325 13337
rect 0 12081 4635 12147
rect 0 11425 4582 12021
rect 0 11129 4310 11365
rect 0 10473 4187 11069
rect 0 10347 3915 10413
rect 0 9117 295 10047
rect 0 8147 267 8837
rect 0 7177 277 7867
rect 0 5967 320 6897
rect 0 4757 305 5687
rect 0 3787 294 4477
rect 0 2577 757 3507
rect 0 1207 470 2297
rect 407 0 1497 254
rect 1777 0 2707 254
rect 2987 0 3677 251
rect 3957 0 4887 254
rect 5167 0 6097 254
rect 6377 0 7067 254
rect 7347 0 8037 254
rect 8317 0 9247 254
rect 9547 0 9613 4715
rect 9673 0 10269 4175
rect 10329 0 10565 4311
rect 10625 0 11221 5382
rect 11281 0 11347 5435
rect 11647 0 12537 254
rect 12817 0 13707 254
rect 14007 0 19000 371
rect 35157 0 40000 254
<< obsm4 >>
rect 367 35877 40000 40800
rect 0 19880 40000 35877
rect 609 14727 40000 19880
rect 0 14587 40000 14727
rect 376 13537 40000 14587
rect 0 13417 40000 13537
rect 405 12367 40000 13417
rect 0 12227 40000 12367
rect 4715 12001 40000 12227
rect 4662 11345 40000 12001
rect 4390 11049 40000 11345
rect 4267 10393 40000 11049
rect 3995 10267 40000 10393
rect 0 10127 40000 10267
rect 375 9037 40000 10127
rect 0 8917 40000 9037
rect 347 8067 40000 8917
rect 0 7947 40000 8067
rect 357 7097 40000 7947
rect 0 6977 40000 7097
rect 400 5887 40000 6977
rect 0 5767 40000 5887
rect 385 5515 40000 5767
rect 385 5462 11201 5515
rect 385 4795 10545 5462
rect 385 4677 9467 4795
rect 0 4557 9467 4677
rect 374 3707 9467 4557
rect 0 3587 9467 3707
rect 837 2497 9467 3587
rect 0 2377 9467 2497
tri 0 1127 80 1207 ne
rect 80 1127 407 1207
rect 550 1127 9467 2377
rect 0 334 9467 1127
rect 0 251 327 334
rect 1577 251 1697 334
rect 2787 331 3877 334
rect 2787 251 2907 331
rect 3757 251 3877 331
rect 4967 251 5087 334
rect 6177 251 6297 334
rect 7147 251 7267 334
rect 8117 251 8237 334
rect 9327 251 9467 334
rect 9693 4391 10545 4795
rect 9693 4255 10249 4391
rect 11427 451 40000 5515
rect 11427 334 13927 451
rect 11427 251 11567 334
rect 12617 251 12737 334
rect 13787 251 13927 334
rect 19080 334 40000 451
rect 19080 251 35077 334
<< metal5 >>
rect 0 14807 529 19797
rect 0 13637 296 14487
rect 0 12467 325 13317
rect 0 10347 4631 12147
rect 0 9137 295 10027
rect 0 8167 267 8817
rect 0 7197 277 7847
rect 0 5987 320 6877
rect 0 4777 305 5667
rect 0 3807 294 4457
rect 0 2597 757 3487
rect 0 1227 470 2277
rect 427 0 1477 254
rect 1797 0 2687 254
rect 3007 0 3657 251
rect 3977 0 4867 254
rect 5187 0 6077 254
rect 6397 0 7047 254
rect 7368 0 8017 254
rect 8337 0 9227 254
rect 9547 0 11347 5431
rect 11667 0 12517 254
rect 12837 0 13687 254
rect 14007 0 18997 371
<< obsm5 >>
rect 0 20117 40000 40800
rect 849 14487 40000 20117
rect 616 13637 40000 14487
rect 645 12467 40000 13637
rect 4951 10027 40000 12467
rect 615 8817 40000 10027
rect 587 8167 40000 8817
rect 597 7197 40000 8167
rect 640 5751 40000 7197
rect 640 5667 9227 5751
rect 625 4457 9227 5667
rect 614 3807 9227 4457
rect 1077 2277 9227 3807
tri 0 907 320 1227 ne
rect 320 907 427 1227
rect 790 907 9227 2277
rect 0 574 9227 907
rect 0 0 107 574
rect 3007 571 3657 574
rect 11667 691 40000 5751
rect 11667 574 13687 691
rect 19317 0 40000 691
<< labels >>
rlabel metal4 s 0 11425 4582 12021 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 10625 0 11221 5382 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 10473 4187 11069 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal4 s 9673 0 10269 4175 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal5 s 0 10347 4631 12147 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 126 11204 128 11206 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 8167 267 8817 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10347 3915 10413 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 8147 267 8837 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 11129 4310 11365 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 12081 4635 12147 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 7368 0 8017 254 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 9547 0 11347 5431 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 10257 126 10259 128 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 11281 0 11347 5435 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 10329 0 10565 4311 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 7347 0 8037 254 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 9547 0 9613 4715 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 3807 294 4457 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 0 3787 294 4477 6 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 3007 0 3657 251 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2987 0 3677 251 6 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 0 7197 277 7847 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal4 s 0 7177 277 7867 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal5 s 6397 0 7047 254 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal4 s 6377 0 7067 254 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal5 s 0 13637 296 14487 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal4 s 0 13617 296 14507 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal5 s 12837 0 13687 254 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal4 s 12817 0 13707 254 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal5 s 0 1227 470 2277 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal4 s 0 1207 470 2297 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal5 s 427 0 1477 254 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal4 s 407 0 1497 254 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal5 s 0 14807 529 19797 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 4777 305 5667 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 4757 305 5687 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 14807 529 19800 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 3977 0 4867 254 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 14007 0 18997 371 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 14007 0 19000 371 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 3957 0 4887 254 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 2597 757 3487 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 0 2577 757 3507 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 1797 0 2687 254 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 1777 0 2707 254 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 0 5987 320 6877 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 5967 320 6897 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 35957 287 40800 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 126 38973 128 38975 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 5187 0 6077 254 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 5167 0 6097 254 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 35157 0 40000 254 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 38173 126 38175 128 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 0 9137 295 10027 6 VSSD
port 11 nsew ground bidirectional
rlabel metal4 s 0 9117 295 10047 6 VSSD
port 11 nsew ground bidirectional
rlabel metal5 s 8337 0 9227 254 6 VSSD
port 11 nsew ground bidirectional
rlabel metal4 s 8317 0 9247 254 6 VSSD
port 11 nsew ground bidirectional
rlabel metal5 s 0 12467 325 13317 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel metal4 s 0 12447 325 13337 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel metal5 s 11667 0 12517 254 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel metal4 s 11647 0 12537 254 6 VSSIO_Q
port 12 nsew ground bidirectional
<< properties >>
string LEFclass ENDCAP TOPRIGHT
string FIXED_BBOX 0 0 40000 40800
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_END 1673972
string GDS_START 1661258
<< end >>
