magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1260 -1236 1404 1288
<< labels >>
flabel comment s 62 25 62 25 2 FreeSans 50 0 0 0 EM1S
flabel comment s 94 27 94 27 0 FreeSans 50 0 0 0 B
flabel comment s 50 27 50 27 0 FreeSans 50 0 0 0 A
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 17385662
string GDS_START 17384958
<< end >>
