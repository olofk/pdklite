magic
tech sky130A
magscale 1 2
timestamp 1640697677
<< pwell >>
rect 894 2323 918 2374
rect 2544 2323 2568 2374
rect 1179 1269 1189 1279
rect 894 821 918 872
rect 2544 821 2568 872
<< obsli1 >>
rect 0 0 3366 3070
<< obsm1 >>
rect 0 3004 3366 3070
rect 0 1568 66 3004
rect 99 2318 127 2976
rect 155 2346 183 3004
rect 211 2318 239 2976
rect 267 2346 295 3004
rect 323 2318 351 2976
rect 379 2346 407 3004
rect 435 2318 463 2976
rect 491 2346 519 3004
rect 547 2318 575 2976
rect 603 2346 631 3004
rect 659 2318 687 2976
rect 715 2346 743 3004
rect 771 2318 799 2976
rect 831 2318 885 2976
rect 917 2318 945 2976
rect 973 2346 1001 3004
rect 1029 2318 1057 2976
rect 1085 2346 1113 3004
rect 1141 2318 1169 2976
rect 1197 2346 1225 3004
rect 1253 2318 1281 2976
rect 1309 2346 1337 3004
rect 1365 2318 1393 2976
rect 1421 2346 1449 3004
rect 1477 2318 1505 2976
rect 1533 2346 1561 3004
rect 1589 2318 1617 2976
rect 99 2254 1617 2318
rect 99 1596 127 2254
rect 155 1568 183 2226
rect 211 1596 239 2254
rect 267 1568 295 2226
rect 323 1596 351 2254
rect 379 1568 407 2226
rect 435 1596 463 2254
rect 491 1568 519 2226
rect 547 1596 575 2254
rect 603 1568 631 2226
rect 659 1596 687 2254
rect 715 1568 743 2226
rect 771 1596 799 2254
rect 831 1596 885 2254
rect 917 1596 945 2254
rect 973 1568 1001 2226
rect 1029 1596 1057 2254
rect 1085 1568 1113 2226
rect 1141 1596 1169 2254
rect 1197 1568 1225 2226
rect 1253 1596 1281 2254
rect 1309 1568 1337 2226
rect 1365 1596 1393 2254
rect 1421 1568 1449 2226
rect 1477 1596 1505 2254
rect 1533 1568 1561 2226
rect 1589 1596 1617 2254
rect 1650 1568 1716 3004
rect 1749 2318 1777 2976
rect 1805 2346 1833 3004
rect 1861 2318 1889 2976
rect 1917 2346 1945 3004
rect 1973 2318 2001 2976
rect 2029 2346 2057 3004
rect 2085 2318 2113 2976
rect 2141 2346 2169 3004
rect 2197 2318 2225 2976
rect 2253 2346 2281 3004
rect 2309 2318 2337 2976
rect 2365 2346 2393 3004
rect 2421 2318 2449 2976
rect 2481 2318 2535 2976
rect 2567 2318 2595 2976
rect 2623 2346 2651 3004
rect 2679 2318 2707 2976
rect 2735 2346 2763 3004
rect 2791 2318 2819 2976
rect 2847 2346 2875 3004
rect 2903 2318 2931 2976
rect 2959 2346 2987 3004
rect 3015 2318 3043 2976
rect 3071 2346 3099 3004
rect 3127 2318 3155 2976
rect 3183 2346 3211 3004
rect 3239 2318 3267 2976
rect 1749 2254 3267 2318
rect 1749 1596 1777 2254
rect 1805 1568 1833 2226
rect 1861 1596 1889 2254
rect 1917 1568 1945 2226
rect 1973 1596 2001 2254
rect 2029 1568 2057 2226
rect 2085 1596 2113 2254
rect 2141 1568 2169 2226
rect 2197 1596 2225 2254
rect 2253 1568 2281 2226
rect 2309 1596 2337 2254
rect 2365 1568 2393 2226
rect 2421 1596 2449 2254
rect 2481 1596 2535 2254
rect 2567 1596 2595 2254
rect 2623 1568 2651 2226
rect 2679 1596 2707 2254
rect 2735 1568 2763 2226
rect 2791 1596 2819 2254
rect 2847 1568 2875 2226
rect 2903 1596 2931 2254
rect 2959 1568 2987 2226
rect 3015 1596 3043 2254
rect 3071 1568 3099 2226
rect 3127 1596 3155 2254
rect 3183 1568 3211 2226
rect 3239 1596 3267 2254
rect 3300 1568 3366 3004
rect 0 1502 3366 1568
rect 0 66 66 1502
rect 99 816 127 1474
rect 155 844 183 1502
rect 211 816 239 1474
rect 267 844 295 1502
rect 323 816 351 1474
rect 379 844 407 1502
rect 435 816 463 1474
rect 491 844 519 1502
rect 547 816 575 1474
rect 603 844 631 1502
rect 659 816 687 1474
rect 715 844 743 1502
rect 771 816 799 1474
rect 831 816 885 1474
rect 917 816 945 1474
rect 973 844 1001 1502
rect 1029 816 1057 1474
rect 1085 844 1113 1502
rect 1141 816 1169 1474
rect 1197 844 1225 1502
rect 1253 816 1281 1474
rect 1309 844 1337 1502
rect 1365 816 1393 1474
rect 1421 844 1449 1502
rect 1477 816 1505 1474
rect 1533 844 1561 1502
rect 1589 816 1617 1474
rect 99 752 1617 816
rect 99 94 127 752
rect 155 66 183 724
rect 211 94 239 752
rect 267 66 295 724
rect 323 94 351 752
rect 379 66 407 724
rect 435 94 463 752
rect 491 66 519 724
rect 547 94 575 752
rect 603 66 631 724
rect 659 94 687 752
rect 715 66 743 724
rect 771 94 799 752
rect 831 94 885 752
rect 917 94 945 752
rect 973 66 1001 724
rect 1029 94 1057 752
rect 1085 66 1113 724
rect 1141 94 1169 752
rect 1197 66 1225 724
rect 1253 94 1281 752
rect 1309 66 1337 724
rect 1365 94 1393 752
rect 1421 66 1449 724
rect 1477 94 1505 752
rect 1533 66 1561 724
rect 1589 94 1617 752
rect 1650 66 1716 1502
rect 1749 816 1777 1474
rect 1805 844 1833 1502
rect 1861 816 1889 1474
rect 1917 844 1945 1502
rect 1973 816 2001 1474
rect 2029 844 2057 1502
rect 2085 816 2113 1474
rect 2141 844 2169 1502
rect 2197 816 2225 1474
rect 2253 844 2281 1502
rect 2309 816 2337 1474
rect 2365 844 2393 1502
rect 2421 816 2449 1474
rect 2481 816 2535 1474
rect 2567 816 2595 1474
rect 2623 844 2651 1502
rect 2679 816 2707 1474
rect 2735 844 2763 1502
rect 2791 816 2819 1474
rect 2847 844 2875 1502
rect 2903 816 2931 1474
rect 2959 844 2987 1502
rect 3015 816 3043 1474
rect 3071 844 3099 1502
rect 3127 816 3155 1474
rect 3183 844 3211 1502
rect 3239 816 3267 1474
rect 1749 752 3267 816
rect 1749 94 1777 752
rect 1805 66 1833 724
rect 1861 94 1889 752
rect 1917 66 1945 724
rect 1973 94 2001 752
rect 2029 66 2057 724
rect 2085 94 2113 752
rect 2141 66 2169 724
rect 2197 94 2225 752
rect 2253 66 2281 724
rect 2309 94 2337 752
rect 2365 66 2393 724
rect 2421 94 2449 752
rect 2481 94 2535 752
rect 2567 94 2595 752
rect 2623 66 2651 724
rect 2679 94 2707 752
rect 2735 66 2763 724
rect 2791 94 2819 752
rect 2847 66 2875 724
rect 2903 94 2931 752
rect 2959 66 2987 724
rect 3015 94 3043 752
rect 3071 66 3099 724
rect 3127 94 3155 752
rect 3183 66 3211 724
rect 3239 94 3267 752
rect 3300 66 3366 1502
rect 0 0 3366 66
<< obsm2 >>
rect 0 3004 803 3070
rect 0 2920 66 3004
rect 831 2976 885 3070
rect 913 3004 2453 3070
rect 94 2948 1622 2976
rect 0 2892 802 2920
rect 0 2808 66 2892
rect 830 2864 886 2948
rect 1650 2920 1716 3004
rect 2481 2976 2535 3070
rect 2563 3004 3366 3070
rect 1744 2948 3272 2976
rect 914 2892 2452 2920
rect 94 2836 1622 2864
rect 0 2780 802 2808
rect 0 2696 66 2780
rect 830 2752 886 2836
rect 1650 2808 1716 2892
rect 2480 2864 2536 2948
rect 3300 2920 3366 3004
rect 2564 2892 3366 2920
rect 1744 2836 3272 2864
rect 914 2780 2452 2808
rect 94 2724 1622 2752
rect 0 2668 802 2696
rect 0 2584 66 2668
rect 830 2640 886 2724
rect 1650 2696 1716 2780
rect 2480 2752 2536 2836
rect 3300 2808 3366 2892
rect 2564 2780 3366 2808
rect 1744 2724 3272 2752
rect 914 2668 2452 2696
rect 94 2612 1622 2640
rect 0 2556 802 2584
rect 0 2472 66 2556
rect 830 2528 886 2612
rect 1650 2584 1716 2668
rect 2480 2640 2536 2724
rect 3300 2696 3366 2780
rect 2564 2668 3366 2696
rect 1744 2612 3272 2640
rect 914 2556 2452 2584
rect 94 2500 1622 2528
rect 0 2444 802 2472
rect 0 2341 66 2444
rect 830 2416 886 2500
rect 1650 2472 1716 2556
rect 2480 2528 2536 2612
rect 3300 2584 3366 2668
rect 2564 2556 3366 2584
rect 1744 2500 3272 2528
rect 914 2444 2452 2472
rect 94 2342 1622 2416
rect 830 2314 886 2342
rect 1650 2341 1716 2444
rect 2480 2416 2536 2500
rect 3300 2472 3366 2556
rect 2564 2444 3366 2472
rect 1744 2342 3272 2416
rect 2480 2314 2536 2342
rect 3300 2341 3366 2444
rect 74 2313 1642 2314
rect 1724 2313 3292 2314
rect 0 2259 3366 2313
rect 74 2258 1642 2259
rect 1724 2258 3292 2259
rect 0 2128 66 2231
rect 830 2230 886 2258
rect 94 2156 1622 2230
rect 0 2100 802 2128
rect 0 2016 66 2100
rect 830 2072 886 2156
rect 1650 2128 1716 2231
rect 2480 2230 2536 2258
rect 1744 2156 3272 2230
rect 914 2100 2452 2128
rect 94 2044 1622 2072
rect 0 1988 802 2016
rect 0 1904 66 1988
rect 830 1960 886 2044
rect 1650 2016 1716 2100
rect 2480 2072 2536 2156
rect 3300 2128 3366 2231
rect 2564 2100 3366 2128
rect 1744 2044 3272 2072
rect 914 1988 2452 2016
rect 94 1932 1622 1960
rect 0 1876 802 1904
rect 0 1792 66 1876
rect 830 1848 886 1932
rect 1650 1904 1716 1988
rect 2480 1960 2536 2044
rect 3300 2016 3366 2100
rect 2564 1988 3366 2016
rect 1744 1932 3272 1960
rect 914 1876 2452 1904
rect 94 1820 1622 1848
rect 0 1764 802 1792
rect 0 1680 66 1764
rect 830 1736 886 1820
rect 1650 1792 1716 1876
rect 2480 1848 2536 1932
rect 3300 1904 3366 1988
rect 2564 1876 3366 1904
rect 1744 1820 3272 1848
rect 914 1764 2452 1792
rect 94 1708 1622 1736
rect 0 1652 802 1680
rect 0 1568 66 1652
rect 830 1624 886 1708
rect 1650 1680 1716 1764
rect 2480 1736 2536 1820
rect 3300 1792 3366 1876
rect 2564 1764 3366 1792
rect 1744 1708 3272 1736
rect 914 1652 2452 1680
rect 94 1596 1622 1624
rect 0 1502 803 1568
rect 0 1418 66 1502
rect 831 1474 885 1596
rect 1650 1568 1716 1652
rect 2480 1624 2536 1708
rect 3300 1680 3366 1764
rect 2564 1652 3366 1680
rect 1744 1596 3272 1624
rect 913 1502 2453 1568
rect 94 1446 1622 1474
rect 0 1390 802 1418
rect 0 1306 66 1390
rect 830 1362 886 1446
rect 1650 1418 1716 1502
rect 2481 1474 2535 1596
rect 3300 1568 3366 1652
rect 2563 1502 3366 1568
rect 1744 1446 3272 1474
rect 914 1390 2452 1418
rect 94 1334 1622 1362
rect 0 1278 802 1306
rect 0 1194 66 1278
rect 830 1250 886 1334
rect 1650 1306 1716 1390
rect 2480 1362 2536 1446
rect 3300 1418 3366 1502
rect 2564 1390 3366 1418
rect 1744 1334 3272 1362
rect 914 1278 2452 1306
rect 94 1222 1622 1250
rect 0 1166 802 1194
rect 0 1082 66 1166
rect 830 1138 886 1222
rect 1650 1194 1716 1278
rect 2480 1250 2536 1334
rect 3300 1306 3366 1390
rect 2564 1278 3366 1306
rect 1744 1222 3272 1250
rect 914 1166 2452 1194
rect 94 1110 1622 1138
rect 0 1054 802 1082
rect 0 970 66 1054
rect 830 1026 886 1110
rect 1650 1082 1716 1166
rect 2480 1138 2536 1222
rect 3300 1194 3366 1278
rect 2564 1166 3366 1194
rect 1744 1110 3272 1138
rect 914 1054 2452 1082
rect 94 998 1622 1026
rect 0 942 802 970
rect 0 839 66 942
rect 830 914 886 998
rect 1650 970 1716 1054
rect 2480 1026 2536 1110
rect 3300 1082 3366 1166
rect 2564 1054 3366 1082
rect 1744 998 3272 1026
rect 914 942 2452 970
rect 94 840 1622 914
rect 830 812 886 840
rect 1650 839 1716 942
rect 2480 914 2536 998
rect 3300 970 3366 1054
rect 2564 942 3366 970
rect 1744 840 3272 914
rect 2480 812 2536 840
rect 3300 839 3366 942
rect 74 811 1642 812
rect 1724 811 3292 812
rect 0 757 3366 811
rect 74 756 1642 757
rect 1724 756 3292 757
rect 0 626 66 729
rect 830 728 886 756
rect 94 654 1622 728
rect 0 598 802 626
rect 0 514 66 598
rect 830 570 886 654
rect 1650 626 1716 729
rect 2480 728 2536 756
rect 1744 654 3272 728
rect 914 598 2452 626
rect 94 542 1622 570
rect 0 486 802 514
rect 0 402 66 486
rect 830 458 886 542
rect 1650 514 1716 598
rect 2480 570 2536 654
rect 3300 626 3366 729
rect 2564 598 3366 626
rect 1744 542 3272 570
rect 914 486 2452 514
rect 94 430 1622 458
rect 0 374 802 402
rect 0 290 66 374
rect 830 346 886 430
rect 1650 402 1716 486
rect 2480 458 2536 542
rect 3300 514 3366 598
rect 2564 486 3366 514
rect 1744 430 3272 458
rect 914 374 2452 402
rect 94 318 1622 346
rect 0 262 802 290
rect 0 178 66 262
rect 830 234 886 318
rect 1650 290 1716 374
rect 2480 346 2536 430
rect 3300 402 3366 486
rect 2564 374 3366 402
rect 1744 318 3272 346
rect 914 262 2452 290
rect 94 206 1622 234
rect 0 150 802 178
rect 0 66 66 150
rect 830 122 886 206
rect 1650 178 1716 262
rect 2480 234 2536 318
rect 3300 290 3366 374
rect 2564 262 3366 290
rect 1744 206 3272 234
rect 914 150 2452 178
rect 94 94 1622 122
rect 0 0 803 66
rect 831 0 885 94
rect 1650 66 1716 150
rect 2480 122 2536 206
rect 3300 178 3366 262
rect 2564 150 3366 178
rect 1744 94 3272 122
rect 913 0 2453 66
rect 2481 0 2535 94
rect 3300 66 3366 150
rect 2563 0 3366 66
<< metal3 >>
rect 0 3004 3366 3070
rect 0 1568 66 3004
rect 126 2319 204 2944
rect 264 2379 342 3004
rect 402 2319 480 2944
rect 540 2379 618 3004
rect 678 2319 756 2944
rect 819 2379 897 3004
rect 960 2319 1038 2944
rect 1098 2379 1176 3004
rect 1236 2319 1314 2944
rect 1374 2379 1452 3004
rect 1512 2319 1590 2944
rect 126 2253 1590 2319
rect 126 1628 204 2253
rect 264 1568 342 2193
rect 402 1628 480 2253
rect 540 1568 618 2193
rect 678 1628 756 2253
rect 819 1568 897 2193
rect 960 1628 1038 2253
rect 1098 1568 1176 2193
rect 1236 1628 1314 2253
rect 1374 1568 1452 2193
rect 1512 1628 1590 2253
rect 1650 1568 1716 3004
rect 1776 2319 1854 2944
rect 1914 2379 1992 3004
rect 2052 2319 2130 2944
rect 2190 2379 2268 3004
rect 2328 2319 2406 2944
rect 2469 2379 2547 3004
rect 2610 2319 2688 2944
rect 2748 2379 2826 3004
rect 2886 2319 2964 2944
rect 3024 2379 3102 3004
rect 3162 2319 3240 2944
rect 1776 2253 3240 2319
rect 1776 1628 1854 2253
rect 1914 1568 1992 2193
rect 2052 1628 2130 2253
rect 2190 1568 2268 2193
rect 2328 1628 2406 2253
rect 2469 1568 2547 2193
rect 2610 1628 2688 2253
rect 2748 1568 2826 2193
rect 2886 1628 2964 2253
rect 3024 1568 3102 2193
rect 3162 1628 3240 2253
rect 3300 1568 3366 3004
rect 0 1502 3366 1568
rect 0 66 66 1502
rect 126 817 204 1442
rect 264 877 342 1502
rect 402 817 480 1442
rect 540 877 618 1502
rect 678 817 756 1442
rect 819 877 897 1502
rect 960 817 1038 1442
rect 1098 877 1176 1502
rect 1236 817 1314 1442
rect 1374 877 1452 1502
rect 1512 817 1590 1442
rect 126 751 1590 817
rect 126 126 204 751
rect 264 66 342 691
rect 402 126 480 751
rect 540 66 618 691
rect 678 126 756 751
rect 819 66 897 691
rect 960 126 1038 751
rect 1098 66 1176 691
rect 1236 126 1314 751
rect 1374 66 1452 691
rect 1512 126 1590 751
rect 1650 66 1716 1502
rect 1776 817 1854 1442
rect 1914 877 1992 1502
rect 2052 817 2130 1442
rect 2190 877 2268 1502
rect 2328 817 2406 1442
rect 2469 877 2547 1502
rect 2610 817 2688 1442
rect 2748 877 2826 1502
rect 2886 817 2964 1442
rect 3024 877 3102 1502
rect 3162 817 3240 1442
rect 1776 751 3240 817
rect 1776 126 1854 751
rect 1914 66 1992 691
rect 2052 126 2130 751
rect 2190 66 2268 691
rect 2328 126 2406 751
rect 2469 66 2547 691
rect 2610 126 2688 751
rect 2748 66 2826 691
rect 2886 126 2964 751
rect 3024 66 3102 691
rect 3162 126 3240 751
rect 3300 66 3366 1502
rect 0 0 3366 66
<< obsm4 >>
rect 63 2605 465 3007
rect 658 2605 1060 3007
rect 1251 2605 1653 3007
rect 1713 2605 2115 3007
rect 2308 2605 2710 3007
rect 2901 2605 3303 3007
rect 63 2086 465 2488
rect 658 2086 1060 2488
rect 1251 2086 1653 2488
rect 1713 2086 2115 2488
rect 2308 2086 2710 2488
rect 2901 2086 3303 2488
rect 63 1565 465 1967
rect 658 1565 1060 1967
rect 1251 1565 1653 1967
rect 1713 1565 2115 1967
rect 2308 1565 2710 1967
rect 2901 1565 3303 1967
rect 63 1103 465 1505
rect 658 1103 1060 1505
rect 1251 1103 1653 1505
rect 1713 1103 2115 1505
rect 2308 1103 2710 1505
rect 2901 1103 3303 1505
rect 63 584 465 986
rect 658 584 1060 986
rect 1251 584 1653 986
rect 1713 584 2115 986
rect 2308 584 2710 986
rect 2901 584 3303 986
rect 63 63 465 465
rect 658 63 1060 465
rect 1251 63 1653 465
rect 1713 63 2115 465
rect 2308 63 2710 465
rect 2901 63 3303 465
<< metal5 >>
rect 0 0 3366 3070
<< labels >>
rlabel metal3 s 3300 1568 3366 3004 6 C0
port 1 nsew
rlabel metal3 s 3300 66 3366 1502 6 C0
port 1 nsew
rlabel metal3 s 3024 2379 3102 3004 6 C0
port 1 nsew
rlabel metal3 s 3024 1568 3102 2193 6 C0
port 1 nsew
rlabel metal3 s 3024 877 3102 1502 6 C0
port 1 nsew
rlabel metal3 s 3024 66 3102 691 6 C0
port 1 nsew
rlabel metal3 s 2748 2379 2826 3004 6 C0
port 1 nsew
rlabel metal3 s 2748 1568 2826 2193 6 C0
port 1 nsew
rlabel metal3 s 2748 877 2826 1502 6 C0
port 1 nsew
rlabel metal3 s 2748 66 2826 691 6 C0
port 1 nsew
rlabel metal3 s 2469 2379 2547 3004 6 C0
port 1 nsew
rlabel metal3 s 2469 1568 2547 2193 6 C0
port 1 nsew
rlabel metal3 s 2469 877 2547 1502 6 C0
port 1 nsew
rlabel metal3 s 2469 66 2547 691 6 C0
port 1 nsew
rlabel metal3 s 2190 2379 2268 3004 6 C0
port 1 nsew
rlabel metal3 s 2190 1568 2268 2193 6 C0
port 1 nsew
rlabel metal3 s 2190 877 2268 1502 6 C0
port 1 nsew
rlabel metal3 s 2190 66 2268 691 6 C0
port 1 nsew
rlabel metal3 s 1914 2379 1992 3004 6 C0
port 1 nsew
rlabel metal3 s 1914 1568 1992 2193 6 C0
port 1 nsew
rlabel metal3 s 1914 877 1992 1502 6 C0
port 1 nsew
rlabel metal3 s 1914 66 1992 691 6 C0
port 1 nsew
rlabel metal3 s 1650 1568 1716 3004 6 C0
port 1 nsew
rlabel metal3 s 1650 66 1716 1502 6 C0
port 1 nsew
rlabel metal3 s 1374 2379 1452 3004 6 C0
port 1 nsew
rlabel metal3 s 1374 1568 1452 2193 6 C0
port 1 nsew
rlabel metal3 s 1374 877 1452 1502 6 C0
port 1 nsew
rlabel metal3 s 1374 66 1452 691 6 C0
port 1 nsew
rlabel metal3 s 1098 2379 1176 3004 6 C0
port 1 nsew
rlabel metal3 s 1098 1568 1176 2193 6 C0
port 1 nsew
rlabel metal3 s 1098 877 1176 1502 6 C0
port 1 nsew
rlabel metal3 s 1098 66 1176 691 6 C0
port 1 nsew
rlabel metal3 s 819 2379 897 3004 6 C0
port 1 nsew
rlabel metal3 s 819 1568 897 2193 6 C0
port 1 nsew
rlabel metal3 s 819 877 897 1502 6 C0
port 1 nsew
rlabel metal3 s 819 66 897 691 6 C0
port 1 nsew
rlabel metal3 s 540 2379 618 3004 6 C0
port 1 nsew
rlabel metal3 s 540 1568 618 2193 6 C0
port 1 nsew
rlabel metal3 s 540 877 618 1502 6 C0
port 1 nsew
rlabel metal3 s 540 66 618 691 6 C0
port 1 nsew
rlabel metal3 s 264 2379 342 3004 6 C0
port 1 nsew
rlabel metal3 s 264 1568 342 2193 6 C0
port 1 nsew
rlabel metal3 s 264 877 342 1502 6 C0
port 1 nsew
rlabel metal3 s 264 66 342 691 6 C0
port 1 nsew
rlabel metal3 s 0 3004 3366 3070 6 C0
port 1 nsew
rlabel metal3 s 0 1568 66 3004 6 C0
port 1 nsew
rlabel metal3 s 0 1502 3366 1568 6 C0
port 1 nsew
rlabel metal3 s 0 66 66 1502 6 C0
port 1 nsew
rlabel metal3 s 0 0 3366 66 6 C0
port 1 nsew
rlabel metal3 s 3162 2319 3240 2944 6 C1
port 2 nsew
rlabel metal3 s 3162 1628 3240 2253 6 C1
port 2 nsew
rlabel metal3 s 3162 817 3240 1442 6 C1
port 2 nsew
rlabel metal3 s 3162 126 3240 751 6 C1
port 2 nsew
rlabel metal3 s 2886 2319 2964 2944 6 C1
port 2 nsew
rlabel metal3 s 2886 1628 2964 2253 6 C1
port 2 nsew
rlabel metal3 s 2886 817 2964 1442 6 C1
port 2 nsew
rlabel metal3 s 2886 126 2964 751 6 C1
port 2 nsew
rlabel metal3 s 2610 2319 2688 2944 6 C1
port 2 nsew
rlabel metal3 s 2610 1628 2688 2253 6 C1
port 2 nsew
rlabel metal3 s 2610 817 2688 1442 6 C1
port 2 nsew
rlabel metal3 s 2610 126 2688 751 6 C1
port 2 nsew
rlabel metal3 s 2328 2319 2406 2944 6 C1
port 2 nsew
rlabel metal3 s 2328 1628 2406 2253 6 C1
port 2 nsew
rlabel metal3 s 2328 817 2406 1442 6 C1
port 2 nsew
rlabel metal3 s 2328 126 2406 751 6 C1
port 2 nsew
rlabel metal3 s 2052 2319 2130 2944 6 C1
port 2 nsew
rlabel metal3 s 2052 1628 2130 2253 6 C1
port 2 nsew
rlabel metal3 s 2052 817 2130 1442 6 C1
port 2 nsew
rlabel metal3 s 2052 126 2130 751 6 C1
port 2 nsew
rlabel metal3 s 1776 2319 1854 2944 6 C1
port 2 nsew
rlabel metal3 s 1776 2253 3240 2319 6 C1
port 2 nsew
rlabel metal3 s 1776 1628 1854 2253 6 C1
port 2 nsew
rlabel metal3 s 1776 817 1854 1442 6 C1
port 2 nsew
rlabel metal3 s 1776 751 3240 817 6 C1
port 2 nsew
rlabel metal3 s 1776 126 1854 751 6 C1
port 2 nsew
rlabel metal3 s 1512 2319 1590 2944 6 C1
port 2 nsew
rlabel metal3 s 1512 1628 1590 2253 6 C1
port 2 nsew
rlabel metal3 s 1512 817 1590 1442 6 C1
port 2 nsew
rlabel metal3 s 1512 126 1590 751 6 C1
port 2 nsew
rlabel metal3 s 1236 2319 1314 2944 6 C1
port 2 nsew
rlabel metal3 s 1236 1628 1314 2253 6 C1
port 2 nsew
rlabel metal3 s 1236 817 1314 1442 6 C1
port 2 nsew
rlabel metal3 s 1236 126 1314 751 6 C1
port 2 nsew
rlabel metal3 s 960 2319 1038 2944 6 C1
port 2 nsew
rlabel metal3 s 960 1628 1038 2253 6 C1
port 2 nsew
rlabel metal3 s 960 817 1038 1442 6 C1
port 2 nsew
rlabel metal3 s 960 126 1038 751 6 C1
port 2 nsew
rlabel metal3 s 678 2319 756 2944 6 C1
port 2 nsew
rlabel metal3 s 678 1628 756 2253 6 C1
port 2 nsew
rlabel metal3 s 678 817 756 1442 6 C1
port 2 nsew
rlabel metal3 s 678 126 756 751 6 C1
port 2 nsew
rlabel metal3 s 402 2319 480 2944 6 C1
port 2 nsew
rlabel metal3 s 402 1628 480 2253 6 C1
port 2 nsew
rlabel metal3 s 402 817 480 1442 6 C1
port 2 nsew
rlabel metal3 s 402 126 480 751 6 C1
port 2 nsew
rlabel metal3 s 126 2319 204 2944 6 C1
port 2 nsew
rlabel metal3 s 126 2253 1590 2319 6 C1
port 2 nsew
rlabel metal3 s 126 1628 204 2253 6 C1
port 2 nsew
rlabel metal3 s 126 817 204 1442 6 C1
port 2 nsew
rlabel metal3 s 126 751 1590 817 6 C1
port 2 nsew
rlabel metal3 s 126 126 204 751 6 C1
port 2 nsew
rlabel metal5 s 0 0 3366 3070 6 M5
port 3 nsew
rlabel pwell s 1179 1269 1189 1279 6 SUB
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 3366 3070
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 380426
string GDS_START 379846
<< end >>
