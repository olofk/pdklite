magic
tech sky130A
magscale 1 2
timestamp 1619729571
<< checkpaint >>
rect -1512 -1494 2595 2038
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 751 47 781 177
rect 835 47 865 177
rect 919 47 949 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 751 297 781 497
rect 835 297 865 497
rect 919 297 949 497
<< ndiff >>
rect 27 129 79 177
rect 27 95 35 129
rect 69 95 79 129
rect 27 47 79 95
rect 109 97 163 177
rect 109 63 119 97
rect 153 63 163 97
rect 109 47 163 63
rect 193 129 247 177
rect 193 95 203 129
rect 237 95 247 129
rect 193 47 247 95
rect 277 97 331 177
rect 277 63 287 97
rect 321 63 331 97
rect 277 47 331 63
rect 361 129 415 177
rect 361 95 371 129
rect 405 95 415 129
rect 361 47 415 95
rect 445 97 499 177
rect 445 63 455 97
rect 489 63 499 97
rect 445 47 499 63
rect 529 129 583 177
rect 529 95 539 129
rect 573 95 583 129
rect 529 47 583 95
rect 613 97 667 177
rect 613 63 623 97
rect 657 63 667 97
rect 613 47 667 63
rect 697 129 751 177
rect 697 95 707 129
rect 741 95 751 129
rect 697 47 751 95
rect 781 97 835 177
rect 781 63 791 97
rect 825 63 835 97
rect 781 47 835 63
rect 865 129 919 177
rect 865 95 875 129
rect 909 95 919 129
rect 865 47 919 95
rect 949 161 1001 177
rect 949 127 959 161
rect 993 127 1001 161
rect 949 93 1001 127
rect 949 59 959 93
rect 993 59 1001 93
rect 949 47 1001 59
<< pdiff >>
rect 27 479 79 497
rect 27 445 35 479
rect 69 445 79 479
rect 27 411 79 445
rect 27 377 35 411
rect 69 377 79 411
rect 27 343 79 377
rect 27 309 35 343
rect 69 309 79 343
rect 27 297 79 309
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 297 163 383
rect 193 479 247 497
rect 193 445 203 479
rect 237 445 247 479
rect 193 411 247 445
rect 193 377 203 411
rect 237 377 247 411
rect 193 343 247 377
rect 193 309 203 343
rect 237 309 247 343
rect 193 297 247 309
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 417 331 451
rect 277 383 287 417
rect 321 383 331 417
rect 277 297 331 383
rect 361 463 415 497
rect 361 429 371 463
rect 405 429 415 463
rect 361 368 415 429
rect 361 334 371 368
rect 405 334 415 368
rect 361 297 415 334
rect 445 485 499 497
rect 445 451 455 485
rect 489 451 499 485
rect 445 417 499 451
rect 445 383 455 417
rect 489 383 499 417
rect 445 297 499 383
rect 529 463 583 497
rect 529 429 539 463
rect 573 429 583 463
rect 529 368 583 429
rect 529 334 539 368
rect 573 334 583 368
rect 529 297 583 334
rect 613 485 667 497
rect 613 451 623 485
rect 657 451 667 485
rect 613 417 667 451
rect 613 383 623 417
rect 657 383 667 417
rect 613 297 667 383
rect 697 463 751 497
rect 697 429 707 463
rect 741 429 751 463
rect 697 368 751 429
rect 697 334 707 368
rect 741 334 751 368
rect 697 297 751 334
rect 781 485 835 497
rect 781 451 791 485
rect 825 451 835 485
rect 781 417 835 451
rect 781 383 791 417
rect 825 383 835 417
rect 781 297 835 383
rect 865 463 919 497
rect 865 429 875 463
rect 909 429 919 463
rect 865 368 919 429
rect 865 334 875 368
rect 909 334 919 368
rect 865 297 919 334
rect 949 485 1001 497
rect 949 451 959 485
rect 993 451 1001 485
rect 949 417 1001 451
rect 949 383 959 417
rect 993 383 1001 417
rect 949 349 1001 383
rect 949 315 959 349
rect 993 315 1001 349
rect 949 297 1001 315
<< ndiffc >>
rect 35 95 69 129
rect 119 63 153 97
rect 203 95 237 129
rect 287 63 321 97
rect 371 95 405 129
rect 455 63 489 97
rect 539 95 573 129
rect 623 63 657 97
rect 707 95 741 129
rect 791 63 825 97
rect 875 95 909 129
rect 959 127 993 161
rect 959 59 993 93
<< pdiffc >>
rect 35 445 69 479
rect 35 377 69 411
rect 35 309 69 343
rect 119 451 153 485
rect 119 383 153 417
rect 203 445 237 479
rect 203 377 237 411
rect 203 309 237 343
rect 287 451 321 485
rect 287 383 321 417
rect 371 429 405 463
rect 371 334 405 368
rect 455 451 489 485
rect 455 383 489 417
rect 539 429 573 463
rect 539 334 573 368
rect 623 451 657 485
rect 623 383 657 417
rect 707 429 741 463
rect 707 334 741 368
rect 791 451 825 485
rect 791 383 825 417
rect 875 429 909 463
rect 875 334 909 368
rect 959 451 993 485
rect 959 383 993 417
rect 959 315 993 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 751 497 781 523
rect 835 497 865 523
rect 919 497 949 523
rect 79 261 109 297
rect 28 259 109 261
rect 163 259 193 297
rect 247 259 277 297
rect 28 249 277 259
rect 28 215 44 249
rect 78 215 112 249
rect 146 215 180 249
rect 214 215 277 249
rect 28 205 277 215
rect 28 203 109 205
rect 79 177 109 203
rect 163 177 193 205
rect 247 177 277 205
rect 331 259 361 297
rect 415 259 445 297
rect 499 259 529 297
rect 583 259 613 297
rect 667 259 697 297
rect 751 259 781 297
rect 835 259 865 297
rect 919 259 949 297
rect 331 249 949 259
rect 331 215 351 249
rect 385 215 419 249
rect 453 215 487 249
rect 521 215 555 249
rect 589 215 623 249
rect 657 215 691 249
rect 725 215 759 249
rect 793 215 949 249
rect 331 205 949 215
rect 331 177 361 205
rect 415 177 445 205
rect 499 177 529 205
rect 583 177 613 205
rect 667 177 697 205
rect 751 177 781 205
rect 835 177 865 205
rect 919 177 949 205
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 751 21 781 47
rect 835 21 865 47
rect 919 21 949 47
<< polycont >>
rect 44 215 78 249
rect 112 215 146 249
rect 180 215 214 249
rect 351 215 385 249
rect 419 215 453 249
rect 487 215 521 249
rect 555 215 589 249
rect 623 215 657 249
rect 691 215 725 249
rect 759 215 793 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 19 479 85 493
rect 19 445 35 479
rect 69 445 85 479
rect 19 411 85 445
rect 19 377 35 411
rect 69 377 85 411
rect 19 343 85 377
rect 119 485 153 527
rect 119 417 153 451
rect 119 367 153 383
rect 187 479 253 493
rect 187 445 203 479
rect 237 445 253 479
rect 187 411 253 445
rect 187 377 203 411
rect 237 377 253 411
rect 19 309 35 343
rect 69 323 85 343
rect 187 343 253 377
rect 287 485 321 527
rect 287 417 321 451
rect 287 367 321 383
rect 371 463 405 493
rect 371 368 405 429
rect 187 323 203 343
rect 69 309 203 323
rect 237 323 253 343
rect 439 485 505 527
rect 439 451 455 485
rect 489 451 505 485
rect 439 417 505 451
rect 439 383 455 417
rect 489 383 505 417
rect 439 367 505 383
rect 539 463 573 493
rect 539 368 573 429
rect 371 323 405 334
rect 607 485 673 527
rect 607 451 623 485
rect 657 451 673 485
rect 607 417 673 451
rect 607 383 623 417
rect 657 383 673 417
rect 607 367 673 383
rect 707 463 741 493
rect 707 368 741 429
rect 539 323 573 334
rect 775 485 841 527
rect 775 451 791 485
rect 825 451 841 485
rect 775 417 841 451
rect 775 383 791 417
rect 825 383 841 417
rect 775 367 841 383
rect 875 463 909 493
rect 875 368 909 429
rect 707 323 741 334
rect 875 323 909 334
rect 237 309 319 323
rect 19 289 319 309
rect 371 289 909 323
rect 943 485 1009 527
rect 943 451 959 485
rect 993 451 1009 485
rect 943 417 1009 451
rect 943 383 959 417
rect 993 383 1009 417
rect 943 349 1009 383
rect 943 315 959 349
rect 993 315 1009 349
rect 943 297 1009 315
rect 28 249 248 255
rect 28 215 44 249
rect 78 215 112 249
rect 146 215 180 249
rect 214 215 248 249
rect 284 249 319 289
rect 858 263 909 289
rect 858 255 974 263
rect 284 215 351 249
rect 385 215 419 249
rect 453 215 487 249
rect 521 215 555 249
rect 589 215 623 249
rect 657 215 691 249
rect 725 215 759 249
rect 793 215 809 249
rect 858 221 861 255
rect 895 221 933 255
rect 967 221 974 255
rect 284 181 319 215
rect 858 211 974 221
rect 858 181 909 211
rect 35 147 319 181
rect 371 147 909 181
rect 35 129 69 147
rect 203 129 237 147
rect 35 51 69 95
rect 103 97 169 113
rect 103 63 119 97
rect 153 63 169 97
rect 103 17 169 63
rect 371 129 405 147
rect 203 52 237 95
rect 271 97 337 113
rect 271 63 287 97
rect 321 63 337 97
rect 271 17 337 63
rect 539 129 573 147
rect 371 51 405 95
rect 439 97 505 113
rect 439 63 455 97
rect 489 63 505 97
rect 439 17 505 63
rect 707 129 741 147
rect 539 51 573 95
rect 607 97 673 113
rect 607 63 623 97
rect 657 63 673 97
rect 607 17 673 63
rect 875 129 909 147
rect 707 51 741 95
rect 775 97 841 113
rect 775 63 791 97
rect 825 63 841 97
rect 775 17 841 63
rect 875 51 909 95
rect 943 161 1009 177
rect 943 127 959 161
rect 993 127 1009 161
rect 943 93 1009 127
rect 943 59 959 93
rect 993 59 1009 93
rect 943 17 1009 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 861 221 895 255
rect 933 221 967 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 570 1104 592
rect 0 561 1046 570
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 0 518 1046 527
rect 1098 518 1110 570
rect 1162 518 1168 570
rect 0 496 1104 518
rect 404 212 410 264
rect 462 212 474 264
rect 526 252 532 264
rect 849 255 979 261
rect 849 252 861 255
rect 526 224 861 252
rect 526 212 532 224
rect 849 221 861 224
rect 895 221 933 255
rect 967 221 979 255
rect 849 215 979 221
rect 0 26 1104 48
rect 0 17 1046 26
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 0 -26 1046 -17
rect 1098 -26 1110 26
rect 1162 -26 1168 26
rect 0 -48 1104 -26
<< via1 >>
rect 1046 561 1098 570
rect 1046 527 1075 561
rect 1075 527 1098 561
rect 1046 518 1098 527
rect 1110 518 1162 570
rect 410 212 462 264
rect 474 212 526 264
rect 1046 17 1098 26
rect 1046 -17 1075 17
rect 1075 -17 1098 17
rect 1046 -26 1098 -17
rect 1110 -26 1162 26
<< metal2 >>
rect 1027 516 1036 572
rect 1092 570 1116 572
rect 1098 518 1110 570
rect 1092 516 1116 518
rect 1172 516 1181 572
rect 378 210 387 266
rect 443 264 467 266
rect 523 264 532 266
rect 462 212 467 264
rect 526 212 532 264
rect 443 210 467 212
rect 523 210 532 212
rect 1027 -28 1036 28
rect 1092 26 1116 28
rect 1098 -26 1110 26
rect 1092 -28 1116 -26
rect 1172 -28 1181 28
<< via2 >>
rect 1036 570 1092 572
rect 1116 570 1172 572
rect 1036 518 1046 570
rect 1046 518 1092 570
rect 1116 518 1162 570
rect 1162 518 1172 570
rect 1036 516 1092 518
rect 1116 516 1172 518
rect 387 264 443 266
rect 467 264 523 266
rect 387 212 410 264
rect 410 212 443 264
rect 467 212 474 264
rect 474 212 523 264
rect 387 210 443 212
rect 467 210 523 212
rect 1036 26 1092 28
rect 1116 26 1172 28
rect 1036 -26 1046 26
rect 1046 -26 1092 26
rect 1116 -26 1162 26
rect 1162 -26 1172 26
rect 1036 -28 1092 -26
rect 1116 -28 1172 -26
<< metal3 >>
rect 1026 576 1182 577
rect 1026 512 1032 576
rect 1096 512 1112 576
rect 1176 512 1182 576
rect 1026 511 1182 512
rect 377 270 533 271
rect -143 206 -137 270
rect -73 206 -57 270
rect 7 206 13 270
rect 377 206 383 270
rect 447 206 463 270
rect 527 206 533 270
rect 377 205 533 206
rect 1026 32 1182 33
rect 1026 -32 1032 32
rect 1096 -32 1112 32
rect 1176 -32 1182 32
rect 1026 -33 1182 -32
<< via3 >>
rect 1032 572 1096 576
rect 1032 516 1036 572
rect 1036 516 1092 572
rect 1092 516 1096 572
rect 1032 512 1096 516
rect 1112 572 1176 576
rect 1112 516 1116 572
rect 1116 516 1172 572
rect 1172 516 1176 572
rect 1112 512 1176 516
rect -137 206 -73 270
rect -57 206 7 270
rect 383 266 447 270
rect 383 210 387 266
rect 387 210 443 266
rect 443 210 447 266
rect 383 206 447 210
rect 463 266 527 270
rect 463 210 467 266
rect 467 210 523 266
rect 523 210 527 266
rect 463 206 527 210
rect 1032 28 1096 32
rect 1032 -28 1036 28
rect 1036 -28 1092 28
rect 1092 -28 1096 28
rect 1032 -32 1096 -28
rect 1112 28 1176 32
rect 1112 -28 1116 28
rect 1116 -28 1172 28
rect 1172 -28 1176 28
rect 1112 -32 1176 -28
<< via4 >>
rect 986 576 1222 723
rect 986 512 1032 576
rect 1032 512 1096 576
rect 1096 512 1112 576
rect 1112 512 1176 576
rect 1176 512 1222 576
rect 986 487 1222 512
rect -228 270 8 390
rect -228 206 -137 270
rect -137 206 -73 270
rect -73 206 -57 270
rect -57 206 7 270
rect 7 206 8 270
rect -228 154 8 206
rect 292 270 528 390
rect 292 206 383 270
rect 383 206 447 270
rect 447 206 463 270
rect 463 206 527 270
rect 527 206 528 270
rect 292 154 528 206
rect 986 32 1222 57
rect 986 -32 1032 32
rect 1032 -32 1096 32
rect 1096 -32 1112 32
rect 1112 -32 1176 32
rect 1176 -32 1222 32
rect 986 -179 1222 -32
<< metal5 >>
rect 232 432 552 765
rect 872 723 1335 778
rect 872 635 986 723
rect 872 595 892 615
rect 912 575 986 635
rect 872 487 986 575
rect 1222 487 1335 723
rect 872 432 1335 487
rect -252 390 552 432
rect -252 154 -228 390
rect 8 154 292 390
rect 528 154 552 390
rect -252 112 552 154
rect 232 -221 552 112
rect 872 57 1335 112
rect 872 -31 986 57
rect 872 -71 892 -51
rect 912 -91 986 -31
rect 872 -179 986 -91
rect 1222 -179 1335 57
rect 872 -234 1335 -179
<< rm5 >>
rect 872 615 912 635
rect 892 595 912 615
rect 872 575 912 595
rect 872 -51 912 -31
rect 892 -71 912 -51
rect 872 -91 912 -71
<< labels >>
flabel metal3 s -98 206 -34 270 0 FreeSans 600 0 0 0 X
port 6 nsew signal output
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel locali s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 probec_p_8
rlabel metal5 s 232 432 552 765 1 X
port 6 nsew signal output
rlabel metal5 s 232 -221 552 112 1 X
port 6 nsew signal output
rlabel metal5 s -252 112 552 432 1 X
port 6 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 4108534
string GDS_START 4095726
<< end >>
