magic
tech sky130A
magscale 1 2
timestamp 1619729571
<< checkpaint >>
rect -1298 -1308 2678 1852
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 30 -17 64 17
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 435 47 465 131
rect 530 47 560 119
rect 621 47 651 119
rect 716 47 746 131
rect 904 47 934 177
rect 988 47 1018 177
rect 1176 47 1206 131
rect 1271 47 1301 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 356 369 386 497
rect 440 369 470 497
rect 536 413 566 497
rect 644 413 674 497
rect 716 413 746 497
rect 904 297 934 497
rect 988 297 1018 497
rect 1176 369 1206 497
rect 1271 297 1301 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 119 351 131
rect 299 85 307 119
rect 341 85 351 119
rect 299 47 351 85
rect 381 89 435 131
rect 381 55 391 89
rect 425 55 435 89
rect 381 47 435 55
rect 465 119 515 131
rect 852 133 904 177
rect 666 119 716 131
rect 465 47 530 119
rect 560 107 621 119
rect 560 73 574 107
rect 608 73 621 107
rect 560 47 621 73
rect 651 47 716 119
rect 746 106 798 131
rect 746 72 756 106
rect 790 72 798 106
rect 746 47 798 72
rect 852 99 860 133
rect 894 99 904 133
rect 852 47 904 99
rect 934 93 988 177
rect 934 59 944 93
rect 978 59 988 93
rect 934 47 988 59
rect 1018 133 1070 177
rect 1018 99 1028 133
rect 1062 99 1070 133
rect 1221 131 1271 177
rect 1018 47 1070 99
rect 1124 119 1176 131
rect 1124 85 1132 119
rect 1166 85 1176 119
rect 1124 47 1176 85
rect 1206 93 1271 131
rect 1206 59 1227 93
rect 1261 59 1271 93
rect 1206 47 1271 59
rect 1301 129 1353 177
rect 1301 95 1311 129
rect 1345 95 1353 129
rect 1301 47 1353 95
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 304 483 356 497
rect 304 449 312 483
rect 346 449 356 483
rect 304 415 356 449
rect 304 381 312 415
rect 346 381 356 415
rect 304 369 356 381
rect 386 485 440 497
rect 386 451 396 485
rect 430 451 440 485
rect 386 417 440 451
rect 386 383 396 417
rect 430 383 440 417
rect 386 369 440 383
rect 470 413 536 497
rect 566 455 644 497
rect 566 421 600 455
rect 634 421 644 455
rect 566 413 644 421
rect 674 413 716 497
rect 746 485 798 497
rect 746 451 756 485
rect 790 451 798 485
rect 746 413 798 451
rect 852 471 904 497
rect 852 437 860 471
rect 894 437 904 471
rect 470 369 520 413
rect 852 368 904 437
rect 852 334 860 368
rect 894 334 904 368
rect 852 297 904 334
rect 934 484 988 497
rect 934 450 944 484
rect 978 450 988 484
rect 934 416 988 450
rect 934 382 944 416
rect 978 382 988 416
rect 934 297 988 382
rect 1018 475 1070 497
rect 1018 441 1028 475
rect 1062 441 1070 475
rect 1018 384 1070 441
rect 1018 350 1028 384
rect 1062 350 1070 384
rect 1124 450 1176 497
rect 1124 416 1132 450
rect 1166 416 1176 450
rect 1124 369 1176 416
rect 1206 485 1271 497
rect 1206 451 1227 485
rect 1261 451 1271 485
rect 1206 417 1271 451
rect 1206 383 1227 417
rect 1261 383 1271 417
rect 1206 369 1271 383
rect 1018 297 1070 350
rect 1221 297 1271 369
rect 1301 449 1353 497
rect 1301 415 1311 449
rect 1345 415 1353 449
rect 1301 381 1353 415
rect 1301 347 1311 381
rect 1345 347 1353 381
rect 1301 297 1353 347
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 85 341 119
rect 391 55 425 89
rect 574 73 608 107
rect 756 72 790 106
rect 860 99 894 133
rect 944 59 978 93
rect 1028 99 1062 133
rect 1132 85 1166 119
rect 1227 59 1261 93
rect 1311 95 1345 129
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 312 449 346 483
rect 312 381 346 415
rect 396 451 430 485
rect 396 383 430 417
rect 600 421 634 455
rect 756 451 790 485
rect 860 437 894 471
rect 860 334 894 368
rect 944 450 978 484
rect 944 382 978 416
rect 1028 441 1062 475
rect 1028 350 1062 384
rect 1132 416 1166 450
rect 1227 451 1261 485
rect 1227 383 1261 417
rect 1311 415 1345 449
rect 1311 347 1345 381
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 356 497 386 523
rect 440 497 470 523
rect 536 497 566 523
rect 644 497 674 523
rect 716 497 746 523
rect 904 497 934 523
rect 988 497 1018 523
rect 1176 497 1206 523
rect 1271 497 1301 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 22 264 76 280
rect 163 274 193 363
rect 356 343 386 369
rect 22 230 32 264
rect 66 230 76 264
rect 22 214 76 230
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 343 313 386 343
rect 343 241 373 313
rect 440 247 470 369
rect 536 337 566 413
rect 644 376 674 413
rect 512 321 566 337
rect 608 366 674 376
rect 608 332 624 366
rect 658 332 674 366
rect 608 325 674 332
rect 609 323 674 325
rect 610 322 674 323
rect 716 373 746 413
rect 716 357 804 373
rect 716 323 760 357
rect 794 323 804 357
rect 512 287 522 321
rect 556 299 566 321
rect 716 307 804 323
rect 556 295 570 299
rect 556 288 575 295
rect 556 287 581 288
rect 512 284 581 287
rect 512 283 588 284
rect 512 282 590 283
rect 512 281 592 282
rect 512 280 599 281
rect 512 279 602 280
rect 512 271 658 279
rect 536 251 658 271
rect 591 250 658 251
rect 594 249 658 250
rect 597 248 658 249
rect 599 247 658 248
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 295 225 373 241
rect 295 191 305 225
rect 339 191 373 225
rect 295 175 373 191
rect 416 231 470 247
rect 601 246 658 247
rect 606 243 658 246
rect 611 239 658 243
rect 614 235 658 239
rect 416 197 426 231
rect 460 197 470 231
rect 416 183 470 197
rect 418 182 470 183
rect 420 181 470 182
rect 513 207 581 209
rect 513 205 582 207
rect 513 199 583 205
rect 343 167 373 175
rect 343 166 374 167
rect 343 164 375 166
rect 343 163 376 164
rect 343 161 377 163
rect 343 160 378 161
rect 343 157 379 160
rect 343 146 381 157
rect 351 131 381 146
rect 435 131 465 181
rect 513 165 533 199
rect 567 165 583 199
rect 513 164 583 165
rect 513 161 582 164
rect 513 158 581 161
rect 513 153 579 158
rect 628 157 658 235
rect 627 156 658 157
rect 625 153 658 156
rect 513 146 560 153
rect 624 151 658 153
rect 623 148 658 151
rect 530 119 560 146
rect 622 145 658 148
rect 621 144 658 145
rect 621 143 657 144
rect 621 142 655 143
rect 621 140 654 142
rect 621 139 653 140
rect 621 137 652 139
rect 621 119 651 137
rect 716 131 746 307
rect 1176 354 1206 369
rect 1175 324 1206 354
rect 904 265 934 297
rect 988 265 1018 297
rect 1175 265 1205 324
rect 1271 265 1301 297
rect 801 249 934 265
rect 801 215 811 249
rect 845 215 934 249
rect 801 199 934 215
rect 984 249 1205 265
rect 984 215 994 249
rect 1028 215 1205 249
rect 984 199 1205 215
rect 1247 249 1301 265
rect 1247 215 1257 249
rect 1291 215 1301 249
rect 1247 199 1301 215
rect 904 177 934 199
rect 988 177 1018 199
rect 1175 176 1205 199
rect 1271 177 1301 199
rect 1175 146 1206 176
rect 1176 131 1206 146
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 435 21 465 47
rect 530 21 560 47
rect 621 21 651 47
rect 716 21 746 47
rect 904 21 934 47
rect 988 21 1018 47
rect 1176 21 1206 47
rect 1271 21 1301 47
<< polycont >>
rect 32 230 66 264
rect 134 230 168 264
rect 624 332 658 366
rect 760 323 794 357
rect 522 287 556 321
rect 305 191 339 225
rect 426 197 460 231
rect 533 165 567 199
rect 811 215 845 249
rect 994 215 1028 249
rect 1257 215 1291 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 396 485 459 527
rect 237 443 248 477
rect 203 409 248 443
rect 69 375 156 393
rect 35 359 156 375
rect 18 264 66 325
rect 18 230 32 264
rect 18 197 66 230
rect 122 323 156 359
rect 122 280 156 289
rect 237 391 248 409
rect 203 357 214 375
rect 203 337 248 357
rect 296 449 312 483
rect 346 449 362 483
rect 296 415 362 449
rect 296 381 312 415
rect 346 381 362 415
rect 122 264 168 280
rect 122 230 134 264
rect 122 214 168 230
rect 122 161 156 214
rect 35 127 156 161
rect 35 119 69 127
rect 203 119 237 337
rect 296 333 362 381
rect 430 451 459 485
rect 756 485 790 527
rect 396 417 459 451
rect 584 421 600 455
rect 634 426 722 455
rect 756 435 790 451
rect 860 471 910 487
rect 894 437 910 471
rect 634 423 723 426
rect 634 421 724 423
rect 430 383 459 417
rect 672 418 725 421
rect 672 415 726 418
rect 675 412 726 415
rect 684 406 726 412
rect 686 403 726 406
rect 396 367 459 383
rect 499 391 556 401
rect 533 357 556 391
rect 296 299 433 333
rect 289 225 357 265
rect 289 191 305 225
rect 339 191 357 225
rect 399 247 433 299
rect 499 321 556 357
rect 499 287 522 321
rect 499 271 556 287
rect 590 366 658 382
rect 590 332 624 366
rect 590 323 658 332
rect 590 289 591 323
rect 625 289 658 323
rect 590 283 658 289
rect 399 231 473 247
rect 399 197 426 231
rect 460 197 473 231
rect 590 207 624 283
rect 692 265 726 403
rect 860 373 910 437
rect 760 368 910 373
rect 760 357 860 368
rect 794 334 860 357
rect 894 334 910 368
rect 944 484 994 527
rect 978 450 994 484
rect 944 416 994 450
rect 978 382 994 416
rect 944 366 994 382
rect 1028 475 1096 493
rect 1062 441 1096 475
rect 1028 384 1096 441
rect 1062 350 1096 384
rect 1028 334 1096 350
rect 794 324 910 334
rect 794 323 916 324
rect 760 307 916 323
rect 879 265 916 307
rect 692 249 845 265
rect 692 233 811 249
rect 399 181 473 197
rect 513 199 624 207
rect 399 157 433 181
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 307 123 433 157
rect 513 165 533 199
rect 567 165 624 199
rect 513 141 624 165
rect 671 215 811 233
rect 671 199 845 215
rect 879 249 1028 265
rect 879 215 994 249
rect 879 199 1028 215
rect 307 119 341 123
rect 671 107 705 199
rect 879 168 916 199
rect 860 133 916 168
rect 1062 149 1096 334
rect 307 69 341 85
rect 103 17 169 59
rect 375 55 391 89
rect 425 55 446 89
rect 558 73 574 107
rect 608 73 705 107
rect 753 106 819 122
rect 375 17 446 55
rect 753 72 756 106
rect 790 72 819 106
rect 894 132 916 133
rect 1028 133 1096 149
rect 1062 99 1096 133
rect 860 83 894 99
rect 928 93 994 99
rect 753 17 819 72
rect 928 59 944 93
rect 978 59 994 93
rect 1028 83 1096 99
rect 1132 450 1182 493
rect 1166 416 1182 450
rect 1132 265 1182 416
rect 1218 485 1277 527
rect 1218 451 1227 485
rect 1261 451 1277 485
rect 1218 417 1277 451
rect 1218 383 1227 417
rect 1261 383 1277 417
rect 1218 367 1277 383
rect 1311 449 1363 493
rect 1345 415 1363 449
rect 1311 381 1363 415
rect 1345 347 1363 381
rect 1311 301 1363 347
rect 1132 249 1291 265
rect 1132 215 1257 249
rect 1132 199 1291 215
rect 1132 119 1182 199
rect 1325 165 1363 301
rect 1166 85 1182 119
rect 1311 129 1363 165
rect 928 17 994 59
rect 1132 51 1182 85
rect 1218 93 1277 109
rect 1218 59 1227 93
rect 1261 59 1277 93
rect 1218 17 1277 59
rect 1345 95 1363 129
rect 1311 51 1363 95
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 122 289 156 323
rect 214 375 237 391
rect 237 375 248 391
rect 214 357 248 375
rect 499 357 533 391
rect 591 289 625 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 487 391 545 397
rect 487 388 499 391
rect 248 360 499 388
rect 248 357 260 360
rect 202 351 260 357
rect 487 357 499 360
rect 533 357 545 391
rect 487 351 545 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 579 323 637 329
rect 579 320 591 323
rect 156 292 591 320
rect 156 289 168 292
rect 110 283 168 289
rect 579 289 591 292
rect 625 289 637 323
rect 579 283 637 289
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
flabel locali s 1319 85 1353 119 0 FreeSans 200 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 315 221 349 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1039 357 1073 391 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1039 425 1073 459 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1039 85 1073 119 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1319 357 1353 391 0 FreeSans 200 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1319 425 1353 459 0 FreeSans 200 0 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 47 544 47 544 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 47 0 47 0 0 FreeSans 200 0 0 0 VGND
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
rlabel comment s 0 0 0 0 4 dlxbn_1
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1380 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 2956822
string GDS_START 2943820
<< end >>
