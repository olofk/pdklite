magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1288 -1260 1408 1357
use sky130_fd_pr__dfl1sd__example_559591418086  sky130_fd_pr__dfl1sd__example_559591418086_0
timestamp 1619729480
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_559591418086  sky130_fd_pr__dfl1sd__example_559591418086_1
timestamp 1619729480
transform 1 0 120 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 148 97 148 97 0 FreeSans 300 0 0 0 D
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 17292794
string GDS_START 17291748
<< end >>
