magic
tech sky130A
magscale 1 2
timestamp 1640697977
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 2 21 719 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
rect 527 47 557 177
rect 611 47 641 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 527 297 557 497
rect 611 297 641 497
<< ndiff >>
rect 28 163 83 177
rect 28 129 39 163
rect 73 129 83 163
rect 28 95 83 129
rect 28 61 39 95
rect 73 61 83 95
rect 28 47 83 61
rect 113 163 167 177
rect 113 129 123 163
rect 157 129 167 163
rect 113 95 167 129
rect 113 61 123 95
rect 157 61 167 95
rect 113 47 167 61
rect 197 95 251 177
rect 197 61 207 95
rect 241 61 251 95
rect 197 47 251 61
rect 281 163 335 177
rect 281 129 291 163
rect 325 129 335 163
rect 281 95 335 129
rect 281 61 291 95
rect 325 61 335 95
rect 281 47 335 61
rect 365 95 417 177
rect 365 61 375 95
rect 409 61 417 95
rect 365 47 417 61
rect 475 95 527 177
rect 475 61 483 95
rect 517 61 527 95
rect 475 47 527 61
rect 557 163 611 177
rect 557 129 567 163
rect 601 129 611 163
rect 557 95 611 129
rect 557 61 567 95
rect 601 61 611 95
rect 557 47 611 61
rect 641 95 693 177
rect 641 61 651 95
rect 685 61 693 95
rect 641 47 693 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 477 167 497
rect 113 443 123 477
rect 157 443 167 477
rect 113 409 167 443
rect 113 375 123 409
rect 157 375 167 409
rect 113 297 167 375
rect 197 477 251 497
rect 197 443 207 477
rect 241 443 251 477
rect 197 409 251 443
rect 197 375 207 409
rect 241 375 251 409
rect 197 341 251 375
rect 197 307 207 341
rect 241 307 251 341
rect 197 297 251 307
rect 281 477 335 497
rect 281 443 291 477
rect 325 443 335 477
rect 281 409 335 443
rect 281 375 291 409
rect 325 375 335 409
rect 281 297 335 375
rect 365 409 421 497
rect 365 375 375 409
rect 409 375 421 409
rect 365 341 421 375
rect 365 307 375 341
rect 409 307 421 341
rect 365 297 421 307
rect 475 477 527 497
rect 475 443 483 477
rect 517 443 527 477
rect 475 409 527 443
rect 475 375 483 409
rect 517 375 527 409
rect 475 297 527 375
rect 557 409 611 497
rect 557 375 567 409
rect 601 375 611 409
rect 557 341 611 375
rect 557 307 567 341
rect 601 307 611 341
rect 557 297 611 307
rect 641 477 693 497
rect 641 443 651 477
rect 685 443 693 477
rect 641 409 693 443
rect 641 375 651 409
rect 685 375 693 409
rect 641 297 693 375
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 123 129 157 163
rect 123 61 157 95
rect 207 61 241 95
rect 291 129 325 163
rect 291 61 325 95
rect 375 61 409 95
rect 483 61 517 95
rect 567 129 601 163
rect 567 61 601 95
rect 651 61 685 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 443 157 477
rect 123 375 157 409
rect 207 443 241 477
rect 207 375 241 409
rect 207 307 241 341
rect 291 443 325 477
rect 291 375 325 409
rect 375 375 409 409
rect 375 307 409 341
rect 483 443 517 477
rect 483 375 517 409
rect 567 375 601 409
rect 567 307 601 341
rect 651 443 685 477
rect 651 375 685 409
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 527 497 557 523
rect 611 497 641 523
rect 83 265 113 297
rect 167 265 197 297
rect 83 249 197 265
rect 83 215 112 249
rect 146 215 197 249
rect 83 199 197 215
rect 83 177 113 199
rect 167 177 197 199
rect 251 265 281 297
rect 335 265 365 297
rect 251 249 365 265
rect 251 215 288 249
rect 322 215 365 249
rect 251 199 365 215
rect 251 177 281 199
rect 335 177 365 199
rect 527 265 557 297
rect 611 265 641 297
rect 527 249 641 265
rect 527 215 543 249
rect 577 215 641 249
rect 527 199 641 215
rect 527 177 557 199
rect 611 177 641 199
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 335 21 365 47
rect 527 21 557 47
rect 611 21 641 47
<< polycont >>
rect 112 215 146 249
rect 288 215 322 249
rect 543 215 577 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 30 477 81 493
rect 30 443 39 477
rect 73 443 81 477
rect 30 409 81 443
rect 30 375 39 409
rect 73 375 81 409
rect 30 341 81 375
rect 115 477 165 527
rect 115 443 123 477
rect 157 443 165 477
rect 115 409 165 443
rect 115 375 123 409
rect 157 375 165 409
rect 115 359 165 375
rect 199 477 249 493
rect 199 443 207 477
rect 241 443 249 477
rect 199 409 249 443
rect 199 375 207 409
rect 241 375 249 409
rect 30 307 39 341
rect 73 325 81 341
rect 199 341 249 375
rect 283 477 693 493
rect 283 443 291 477
rect 325 459 483 477
rect 325 443 333 459
rect 283 409 333 443
rect 517 459 651 477
rect 517 443 525 459
rect 283 375 291 409
rect 325 375 333 409
rect 283 359 333 375
rect 367 409 417 425
rect 367 375 375 409
rect 409 375 417 409
rect 199 325 207 341
rect 73 307 207 325
rect 241 325 249 341
rect 367 341 417 375
rect 483 409 525 443
rect 643 443 651 459
rect 685 443 693 477
rect 517 375 525 409
rect 483 359 525 375
rect 567 409 609 425
rect 601 375 609 409
rect 367 325 375 341
rect 241 307 375 325
rect 409 307 417 341
rect 567 341 609 375
rect 643 409 693 443
rect 643 375 651 409
rect 685 375 693 409
rect 643 359 693 375
rect 30 291 417 307
rect 475 257 528 325
rect 601 325 609 341
rect 601 307 719 325
rect 567 291 719 307
rect 27 249 193 257
rect 27 215 112 249
rect 146 215 193 249
rect 227 249 437 257
rect 227 215 288 249
rect 322 215 437 249
rect 475 249 593 257
rect 475 215 543 249
rect 577 215 593 249
rect 627 181 719 291
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 107 163 719 181
rect 107 129 123 163
rect 157 145 291 163
rect 157 129 173 145
rect 107 95 173 129
rect 275 129 291 145
rect 325 145 567 163
rect 325 129 341 145
rect 107 61 123 95
rect 157 61 173 95
rect 107 51 173 61
rect 207 95 241 111
rect 207 17 241 61
rect 275 95 341 129
rect 551 129 567 145
rect 601 145 719 163
rect 601 129 617 145
rect 275 61 291 95
rect 325 61 341 95
rect 275 51 341 61
rect 375 95 517 111
rect 409 61 483 95
rect 375 17 517 61
rect 551 95 617 129
rect 551 61 567 95
rect 601 61 617 95
rect 551 51 617 61
rect 651 95 709 111
rect 685 61 709 95
rect 651 17 709 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 494 221 528 255 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 678 289 712 323 0 FreeSans 400 0 0 0 Y
port 8 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor3_2
rlabel metal1 s 0 -48 736 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 2020068
string GDS_START 2013520
string path 0.000 0.000 18.400 0.000 
<< end >>
