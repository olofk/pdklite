magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1260 -853 16260 41260
<< metal3 >>
rect 99 18950 4018 18953
rect 99 18886 162 18950
rect 226 18886 243 18950
rect 307 18886 324 18950
rect 388 18886 405 18950
rect 469 18886 486 18950
rect 550 18886 567 18950
rect 631 18886 648 18950
rect 712 18886 729 18950
rect 793 18886 810 18950
rect 874 18886 891 18950
rect 955 18886 972 18950
rect 1036 18886 1053 18950
rect 1117 18886 1134 18950
rect 1198 18886 1215 18950
rect 1279 18886 1296 18950
rect 1360 18886 1377 18950
rect 1441 18886 1458 18950
rect 1522 18886 1539 18950
rect 1603 18886 1620 18950
rect 1684 18886 1701 18950
rect 1765 18886 1782 18950
rect 1846 18886 1863 18950
rect 1927 18886 1944 18950
rect 2008 18886 2025 18950
rect 2089 18886 2106 18950
rect 2170 18886 2187 18950
rect 2251 18886 2268 18950
rect 2332 18886 2349 18950
rect 2413 18886 2430 18950
rect 2494 18886 2511 18950
rect 2575 18886 2592 18950
rect 2656 18886 2673 18950
rect 2737 18886 2754 18950
rect 2818 18886 2835 18950
rect 2899 18886 2916 18950
rect 2980 18886 2997 18950
rect 3061 18886 3078 18950
rect 3142 18886 3159 18950
rect 3223 18886 3240 18950
rect 3304 18886 3321 18950
rect 3385 18886 3402 18950
rect 3466 18886 3483 18950
rect 3547 18886 3563 18950
rect 3627 18886 3643 18950
rect 3707 18886 3723 18950
rect 3787 18886 3803 18950
rect 3867 18886 3883 18950
rect 3947 18886 4018 18950
rect 99 18866 4018 18886
rect 99 18802 162 18866
rect 226 18802 243 18866
rect 307 18802 324 18866
rect 388 18802 405 18866
rect 469 18802 486 18866
rect 550 18802 567 18866
rect 631 18802 648 18866
rect 712 18802 729 18866
rect 793 18802 810 18866
rect 874 18802 891 18866
rect 955 18802 972 18866
rect 1036 18802 1053 18866
rect 1117 18802 1134 18866
rect 1198 18802 1215 18866
rect 1279 18802 1296 18866
rect 1360 18802 1377 18866
rect 1441 18802 1458 18866
rect 1522 18802 1539 18866
rect 1603 18802 1620 18866
rect 1684 18802 1701 18866
rect 1765 18802 1782 18866
rect 1846 18802 1863 18866
rect 1927 18802 1944 18866
rect 2008 18802 2025 18866
rect 2089 18802 2106 18866
rect 2170 18802 2187 18866
rect 2251 18802 2268 18866
rect 2332 18802 2349 18866
rect 2413 18802 2430 18866
rect 2494 18802 2511 18866
rect 2575 18802 2592 18866
rect 2656 18802 2673 18866
rect 2737 18802 2754 18866
rect 2818 18802 2835 18866
rect 2899 18802 2916 18866
rect 2980 18802 2997 18866
rect 3061 18802 3078 18866
rect 3142 18802 3159 18866
rect 3223 18802 3240 18866
rect 3304 18802 3321 18866
rect 3385 18802 3402 18866
rect 3466 18802 3483 18866
rect 3547 18802 3563 18866
rect 3627 18802 3643 18866
rect 3707 18802 3723 18866
rect 3787 18802 3803 18866
rect 3867 18802 3883 18866
rect 3947 18802 4018 18866
rect 99 18782 4018 18802
rect 99 18718 162 18782
rect 226 18718 243 18782
rect 307 18718 324 18782
rect 388 18718 405 18782
rect 469 18718 486 18782
rect 550 18718 567 18782
rect 631 18718 648 18782
rect 712 18718 729 18782
rect 793 18718 810 18782
rect 874 18718 891 18782
rect 955 18718 972 18782
rect 1036 18718 1053 18782
rect 1117 18718 1134 18782
rect 1198 18718 1215 18782
rect 1279 18718 1296 18782
rect 1360 18718 1377 18782
rect 1441 18718 1458 18782
rect 1522 18718 1539 18782
rect 1603 18718 1620 18782
rect 1684 18718 1701 18782
rect 1765 18718 1782 18782
rect 1846 18718 1863 18782
rect 1927 18718 1944 18782
rect 2008 18718 2025 18782
rect 2089 18718 2106 18782
rect 2170 18718 2187 18782
rect 2251 18718 2268 18782
rect 2332 18718 2349 18782
rect 2413 18718 2430 18782
rect 2494 18718 2511 18782
rect 2575 18718 2592 18782
rect 2656 18718 2673 18782
rect 2737 18718 2754 18782
rect 2818 18718 2835 18782
rect 2899 18718 2916 18782
rect 2980 18718 2997 18782
rect 3061 18718 3078 18782
rect 3142 18718 3159 18782
rect 3223 18718 3240 18782
rect 3304 18718 3321 18782
rect 3385 18718 3402 18782
rect 3466 18718 3483 18782
rect 3547 18718 3563 18782
rect 3627 18718 3643 18782
rect 3707 18718 3723 18782
rect 3787 18718 3803 18782
rect 3867 18718 3883 18782
rect 3947 18771 4018 18782
tri 4018 18771 4200 18953 sw
tri 10812 18771 10994 18953 se
rect 10994 18950 14858 18953
rect 10994 18886 11065 18950
rect 11129 18886 11145 18950
rect 11209 18886 11225 18950
rect 11289 18886 11305 18950
rect 11369 18886 11385 18950
rect 11449 18886 11465 18950
rect 11529 18886 11546 18950
rect 11610 18886 11627 18950
rect 11691 18886 11708 18950
rect 11772 18886 11789 18950
rect 11853 18886 11870 18950
rect 11934 18886 11951 18950
rect 12015 18886 12032 18950
rect 12096 18886 12113 18950
rect 12177 18886 12194 18950
rect 12258 18886 12275 18950
rect 12339 18886 12356 18950
rect 12420 18886 12437 18950
rect 12501 18886 12518 18950
rect 12582 18886 12599 18950
rect 12663 18886 12680 18950
rect 12744 18886 12761 18950
rect 12825 18886 12842 18950
rect 12906 18886 12923 18950
rect 12987 18886 13004 18950
rect 13068 18886 13085 18950
rect 13149 18886 13166 18950
rect 13230 18886 13247 18950
rect 13311 18886 13328 18950
rect 13392 18886 13409 18950
rect 13473 18886 13490 18950
rect 13554 18886 13571 18950
rect 13635 18886 13652 18950
rect 13716 18886 13733 18950
rect 13797 18886 13814 18950
rect 13878 18886 13895 18950
rect 13959 18886 13976 18950
rect 14040 18886 14057 18950
rect 14121 18886 14138 18950
rect 14202 18886 14219 18950
rect 14283 18886 14300 18950
rect 14364 18886 14381 18950
rect 14445 18886 14462 18950
rect 14526 18886 14543 18950
rect 14607 18886 14624 18950
rect 14688 18886 14705 18950
rect 14769 18886 14786 18950
rect 14850 18886 14858 18950
rect 10994 18866 14858 18886
rect 10994 18802 11065 18866
rect 11129 18802 11145 18866
rect 11209 18802 11225 18866
rect 11289 18802 11305 18866
rect 11369 18802 11385 18866
rect 11449 18802 11465 18866
rect 11529 18802 11546 18866
rect 11610 18802 11627 18866
rect 11691 18802 11708 18866
rect 11772 18802 11789 18866
rect 11853 18802 11870 18866
rect 11934 18802 11951 18866
rect 12015 18802 12032 18866
rect 12096 18802 12113 18866
rect 12177 18802 12194 18866
rect 12258 18802 12275 18866
rect 12339 18802 12356 18866
rect 12420 18802 12437 18866
rect 12501 18802 12518 18866
rect 12582 18802 12599 18866
rect 12663 18802 12680 18866
rect 12744 18802 12761 18866
rect 12825 18802 12842 18866
rect 12906 18802 12923 18866
rect 12987 18802 13004 18866
rect 13068 18802 13085 18866
rect 13149 18802 13166 18866
rect 13230 18802 13247 18866
rect 13311 18802 13328 18866
rect 13392 18802 13409 18866
rect 13473 18802 13490 18866
rect 13554 18802 13571 18866
rect 13635 18802 13652 18866
rect 13716 18802 13733 18866
rect 13797 18802 13814 18866
rect 13878 18802 13895 18866
rect 13959 18802 13976 18866
rect 14040 18802 14057 18866
rect 14121 18802 14138 18866
rect 14202 18802 14219 18866
rect 14283 18802 14300 18866
rect 14364 18802 14381 18866
rect 14445 18802 14462 18866
rect 14526 18802 14543 18866
rect 14607 18802 14624 18866
rect 14688 18802 14705 18866
rect 14769 18802 14786 18866
rect 14850 18802 14858 18866
rect 10994 18782 14858 18802
rect 10994 18771 11065 18782
rect 3947 18765 4200 18771
rect 3947 18718 3994 18765
rect 99 18701 3994 18718
rect 4058 18701 4124 18765
rect 4188 18701 4200 18765
rect 99 18698 4200 18701
rect 99 18634 162 18698
rect 226 18634 243 18698
rect 307 18634 324 18698
rect 388 18634 405 18698
rect 469 18634 486 18698
rect 550 18634 567 18698
rect 631 18634 648 18698
rect 712 18634 729 18698
rect 793 18634 810 18698
rect 874 18634 891 18698
rect 955 18634 972 18698
rect 1036 18634 1053 18698
rect 1117 18634 1134 18698
rect 1198 18634 1215 18698
rect 1279 18634 1296 18698
rect 1360 18634 1377 18698
rect 1441 18634 1458 18698
rect 1522 18634 1539 18698
rect 1603 18634 1620 18698
rect 1684 18634 1701 18698
rect 1765 18634 1782 18698
rect 1846 18634 1863 18698
rect 1927 18634 1944 18698
rect 2008 18634 2025 18698
rect 2089 18634 2106 18698
rect 2170 18634 2187 18698
rect 2251 18634 2268 18698
rect 2332 18634 2349 18698
rect 2413 18634 2430 18698
rect 2494 18634 2511 18698
rect 2575 18634 2592 18698
rect 2656 18634 2673 18698
rect 2737 18634 2754 18698
rect 2818 18634 2835 18698
rect 2899 18634 2916 18698
rect 2980 18634 2997 18698
rect 3061 18634 3078 18698
rect 3142 18634 3159 18698
rect 3223 18634 3240 18698
rect 3304 18634 3321 18698
rect 3385 18634 3402 18698
rect 3466 18634 3483 18698
rect 3547 18634 3563 18698
rect 3627 18634 3643 18698
rect 3707 18634 3723 18698
rect 3787 18634 3803 18698
rect 3867 18634 3883 18698
rect 3947 18643 4200 18698
rect 3947 18634 3994 18643
rect 99 18614 3994 18634
rect 99 18550 162 18614
rect 226 18550 243 18614
rect 307 18550 324 18614
rect 388 18550 405 18614
rect 469 18550 486 18614
rect 550 18550 567 18614
rect 631 18550 648 18614
rect 712 18550 729 18614
rect 793 18550 810 18614
rect 874 18550 891 18614
rect 955 18550 972 18614
rect 1036 18550 1053 18614
rect 1117 18550 1134 18614
rect 1198 18550 1215 18614
rect 1279 18550 1296 18614
rect 1360 18550 1377 18614
rect 1441 18550 1458 18614
rect 1522 18550 1539 18614
rect 1603 18550 1620 18614
rect 1684 18550 1701 18614
rect 1765 18550 1782 18614
rect 1846 18550 1863 18614
rect 1927 18550 1944 18614
rect 2008 18550 2025 18614
rect 2089 18550 2106 18614
rect 2170 18550 2187 18614
rect 2251 18550 2268 18614
rect 2332 18550 2349 18614
rect 2413 18550 2430 18614
rect 2494 18550 2511 18614
rect 2575 18550 2592 18614
rect 2656 18550 2673 18614
rect 2737 18550 2754 18614
rect 2818 18550 2835 18614
rect 2899 18550 2916 18614
rect 2980 18550 2997 18614
rect 3061 18550 3078 18614
rect 3142 18550 3159 18614
rect 3223 18550 3240 18614
rect 3304 18550 3321 18614
rect 3385 18550 3402 18614
rect 3466 18550 3483 18614
rect 3547 18550 3563 18614
rect 3627 18550 3643 18614
rect 3707 18550 3723 18614
rect 3787 18550 3803 18614
rect 3867 18550 3883 18614
rect 3947 18579 3994 18614
rect 4058 18579 4124 18643
rect 4188 18579 4200 18643
rect 3947 18573 4200 18579
tri 4200 18573 4398 18771 sw
tri 10614 18573 10812 18771 se
rect 10812 18765 11065 18771
rect 10812 18701 10824 18765
rect 10888 18701 10954 18765
rect 11018 18718 11065 18765
rect 11129 18718 11145 18782
rect 11209 18718 11225 18782
rect 11289 18718 11305 18782
rect 11369 18718 11385 18782
rect 11449 18718 11465 18782
rect 11529 18718 11546 18782
rect 11610 18718 11627 18782
rect 11691 18718 11708 18782
rect 11772 18718 11789 18782
rect 11853 18718 11870 18782
rect 11934 18718 11951 18782
rect 12015 18718 12032 18782
rect 12096 18718 12113 18782
rect 12177 18718 12194 18782
rect 12258 18718 12275 18782
rect 12339 18718 12356 18782
rect 12420 18718 12437 18782
rect 12501 18718 12518 18782
rect 12582 18718 12599 18782
rect 12663 18718 12680 18782
rect 12744 18718 12761 18782
rect 12825 18718 12842 18782
rect 12906 18718 12923 18782
rect 12987 18718 13004 18782
rect 13068 18718 13085 18782
rect 13149 18718 13166 18782
rect 13230 18718 13247 18782
rect 13311 18718 13328 18782
rect 13392 18718 13409 18782
rect 13473 18718 13490 18782
rect 13554 18718 13571 18782
rect 13635 18718 13652 18782
rect 13716 18718 13733 18782
rect 13797 18718 13814 18782
rect 13878 18718 13895 18782
rect 13959 18718 13976 18782
rect 14040 18718 14057 18782
rect 14121 18718 14138 18782
rect 14202 18718 14219 18782
rect 14283 18718 14300 18782
rect 14364 18718 14381 18782
rect 14445 18718 14462 18782
rect 14526 18718 14543 18782
rect 14607 18718 14624 18782
rect 14688 18718 14705 18782
rect 14769 18718 14786 18782
rect 14850 18718 14858 18782
rect 11018 18701 14858 18718
rect 10812 18698 14858 18701
rect 10812 18643 11065 18698
rect 10812 18579 10824 18643
rect 10888 18579 10954 18643
rect 11018 18634 11065 18643
rect 11129 18634 11145 18698
rect 11209 18634 11225 18698
rect 11289 18634 11305 18698
rect 11369 18634 11385 18698
rect 11449 18634 11465 18698
rect 11529 18634 11546 18698
rect 11610 18634 11627 18698
rect 11691 18634 11708 18698
rect 11772 18634 11789 18698
rect 11853 18634 11870 18698
rect 11934 18634 11951 18698
rect 12015 18634 12032 18698
rect 12096 18634 12113 18698
rect 12177 18634 12194 18698
rect 12258 18634 12275 18698
rect 12339 18634 12356 18698
rect 12420 18634 12437 18698
rect 12501 18634 12518 18698
rect 12582 18634 12599 18698
rect 12663 18634 12680 18698
rect 12744 18634 12761 18698
rect 12825 18634 12842 18698
rect 12906 18634 12923 18698
rect 12987 18634 13004 18698
rect 13068 18634 13085 18698
rect 13149 18634 13166 18698
rect 13230 18634 13247 18698
rect 13311 18634 13328 18698
rect 13392 18634 13409 18698
rect 13473 18634 13490 18698
rect 13554 18634 13571 18698
rect 13635 18634 13652 18698
rect 13716 18634 13733 18698
rect 13797 18634 13814 18698
rect 13878 18634 13895 18698
rect 13959 18634 13976 18698
rect 14040 18634 14057 18698
rect 14121 18634 14138 18698
rect 14202 18634 14219 18698
rect 14283 18634 14300 18698
rect 14364 18634 14381 18698
rect 14445 18634 14462 18698
rect 14526 18634 14543 18698
rect 14607 18634 14624 18698
rect 14688 18634 14705 18698
rect 14769 18634 14786 18698
rect 14850 18634 14858 18698
rect 11018 18614 14858 18634
rect 11018 18579 11065 18614
rect 10812 18573 11065 18579
rect 3947 18550 4398 18573
rect 99 18530 4398 18550
rect 99 18466 162 18530
rect 226 18466 243 18530
rect 307 18466 324 18530
rect 388 18466 405 18530
rect 469 18466 486 18530
rect 550 18466 567 18530
rect 631 18466 648 18530
rect 712 18466 729 18530
rect 793 18466 810 18530
rect 874 18466 891 18530
rect 955 18466 972 18530
rect 1036 18466 1053 18530
rect 1117 18466 1134 18530
rect 1198 18466 1215 18530
rect 1279 18466 1296 18530
rect 1360 18466 1377 18530
rect 1441 18466 1458 18530
rect 1522 18466 1539 18530
rect 1603 18466 1620 18530
rect 1684 18466 1701 18530
rect 1765 18466 1782 18530
rect 1846 18466 1863 18530
rect 1927 18466 1944 18530
rect 2008 18466 2025 18530
rect 2089 18466 2106 18530
rect 2170 18466 2187 18530
rect 2251 18466 2268 18530
rect 2332 18466 2349 18530
rect 2413 18466 2430 18530
rect 2494 18466 2511 18530
rect 2575 18466 2592 18530
rect 2656 18466 2673 18530
rect 2737 18466 2754 18530
rect 2818 18466 2835 18530
rect 2899 18466 2916 18530
rect 2980 18466 2997 18530
rect 3061 18466 3078 18530
rect 3142 18466 3159 18530
rect 3223 18466 3240 18530
rect 3304 18466 3321 18530
rect 3385 18466 3402 18530
rect 3466 18466 3483 18530
rect 3547 18466 3563 18530
rect 3627 18466 3643 18530
rect 3707 18466 3723 18530
rect 3787 18466 3803 18530
rect 3867 18466 3883 18530
rect 3947 18514 4398 18530
tri 4398 18514 4457 18573 sw
tri 10555 18514 10614 18573 se
rect 10614 18550 11065 18573
rect 11129 18550 11145 18614
rect 11209 18550 11225 18614
rect 11289 18550 11305 18614
rect 11369 18550 11385 18614
rect 11449 18550 11465 18614
rect 11529 18550 11546 18614
rect 11610 18550 11627 18614
rect 11691 18550 11708 18614
rect 11772 18550 11789 18614
rect 11853 18550 11870 18614
rect 11934 18550 11951 18614
rect 12015 18550 12032 18614
rect 12096 18550 12113 18614
rect 12177 18550 12194 18614
rect 12258 18550 12275 18614
rect 12339 18550 12356 18614
rect 12420 18550 12437 18614
rect 12501 18550 12518 18614
rect 12582 18550 12599 18614
rect 12663 18550 12680 18614
rect 12744 18550 12761 18614
rect 12825 18550 12842 18614
rect 12906 18550 12923 18614
rect 12987 18550 13004 18614
rect 13068 18550 13085 18614
rect 13149 18550 13166 18614
rect 13230 18550 13247 18614
rect 13311 18550 13328 18614
rect 13392 18550 13409 18614
rect 13473 18550 13490 18614
rect 13554 18550 13571 18614
rect 13635 18550 13652 18614
rect 13716 18550 13733 18614
rect 13797 18550 13814 18614
rect 13878 18550 13895 18614
rect 13959 18550 13976 18614
rect 14040 18550 14057 18614
rect 14121 18550 14138 18614
rect 14202 18550 14219 18614
rect 14283 18550 14300 18614
rect 14364 18550 14381 18614
rect 14445 18550 14462 18614
rect 14526 18550 14543 18614
rect 14607 18550 14624 18614
rect 14688 18550 14705 18614
rect 14769 18550 14786 18614
rect 14850 18550 14858 18614
rect 10614 18530 14858 18550
rect 10614 18514 11065 18530
rect 3947 18512 4457 18514
rect 3947 18466 4016 18512
rect 99 18448 4016 18466
rect 4080 18448 4129 18512
rect 4193 18448 4242 18512
rect 4306 18448 4355 18512
rect 4419 18448 4457 18512
rect 99 18446 4457 18448
rect 99 18382 162 18446
rect 226 18382 243 18446
rect 307 18382 324 18446
rect 388 18382 405 18446
rect 469 18382 486 18446
rect 550 18382 567 18446
rect 631 18382 648 18446
rect 712 18382 729 18446
rect 793 18382 810 18446
rect 874 18382 891 18446
rect 955 18382 972 18446
rect 1036 18382 1053 18446
rect 1117 18382 1134 18446
rect 1198 18382 1215 18446
rect 1279 18382 1296 18446
rect 1360 18382 1377 18446
rect 1441 18382 1458 18446
rect 1522 18382 1539 18446
rect 1603 18382 1620 18446
rect 1684 18382 1701 18446
rect 1765 18382 1782 18446
rect 1846 18382 1863 18446
rect 1927 18382 1944 18446
rect 2008 18382 2025 18446
rect 2089 18382 2106 18446
rect 2170 18382 2187 18446
rect 2251 18382 2268 18446
rect 2332 18382 2349 18446
rect 2413 18382 2430 18446
rect 2494 18382 2511 18446
rect 2575 18382 2592 18446
rect 2656 18382 2673 18446
rect 2737 18382 2754 18446
rect 2818 18382 2835 18446
rect 2899 18382 2916 18446
rect 2980 18382 2997 18446
rect 3061 18382 3078 18446
rect 3142 18382 3159 18446
rect 3223 18382 3240 18446
rect 3304 18382 3321 18446
rect 3385 18382 3402 18446
rect 3466 18382 3483 18446
rect 3547 18382 3563 18446
rect 3627 18382 3643 18446
rect 3707 18382 3723 18446
rect 3787 18382 3803 18446
rect 3867 18382 3883 18446
rect 3947 18410 4457 18446
rect 3947 18382 4016 18410
rect 99 18362 4016 18382
rect 99 18298 162 18362
rect 226 18298 243 18362
rect 307 18298 324 18362
rect 388 18298 405 18362
rect 469 18298 486 18362
rect 550 18298 567 18362
rect 631 18298 648 18362
rect 712 18298 729 18362
rect 793 18298 810 18362
rect 874 18298 891 18362
rect 955 18298 972 18362
rect 1036 18298 1053 18362
rect 1117 18298 1134 18362
rect 1198 18298 1215 18362
rect 1279 18298 1296 18362
rect 1360 18298 1377 18362
rect 1441 18298 1458 18362
rect 1522 18298 1539 18362
rect 1603 18298 1620 18362
rect 1684 18298 1701 18362
rect 1765 18298 1782 18362
rect 1846 18298 1863 18362
rect 1927 18298 1944 18362
rect 2008 18298 2025 18362
rect 2089 18298 2106 18362
rect 2170 18298 2187 18362
rect 2251 18298 2268 18362
rect 2332 18298 2349 18362
rect 2413 18298 2430 18362
rect 2494 18298 2511 18362
rect 2575 18298 2592 18362
rect 2656 18298 2673 18362
rect 2737 18298 2754 18362
rect 2818 18298 2835 18362
rect 2899 18298 2916 18362
rect 2980 18298 2997 18362
rect 3061 18298 3078 18362
rect 3142 18298 3159 18362
rect 3223 18298 3240 18362
rect 3304 18298 3321 18362
rect 3385 18298 3402 18362
rect 3466 18298 3483 18362
rect 3547 18298 3563 18362
rect 3627 18298 3643 18362
rect 3707 18298 3723 18362
rect 3787 18298 3803 18362
rect 3867 18298 3883 18362
rect 3947 18346 4016 18362
rect 4080 18346 4129 18410
rect 4193 18346 4242 18410
rect 4306 18346 4355 18410
rect 4419 18346 4457 18410
rect 3947 18308 4457 18346
rect 3947 18298 4016 18308
rect 99 18278 4016 18298
rect 99 18214 162 18278
rect 226 18214 243 18278
rect 307 18214 324 18278
rect 388 18214 405 18278
rect 469 18214 486 18278
rect 550 18214 567 18278
rect 631 18214 648 18278
rect 712 18214 729 18278
rect 793 18214 810 18278
rect 874 18214 891 18278
rect 955 18214 972 18278
rect 1036 18214 1053 18278
rect 1117 18214 1134 18278
rect 1198 18214 1215 18278
rect 1279 18214 1296 18278
rect 1360 18214 1377 18278
rect 1441 18214 1458 18278
rect 1522 18214 1539 18278
rect 1603 18214 1620 18278
rect 1684 18214 1701 18278
rect 1765 18214 1782 18278
rect 1846 18214 1863 18278
rect 1927 18214 1944 18278
rect 2008 18214 2025 18278
rect 2089 18214 2106 18278
rect 2170 18214 2187 18278
rect 2251 18214 2268 18278
rect 2332 18214 2349 18278
rect 2413 18214 2430 18278
rect 2494 18214 2511 18278
rect 2575 18214 2592 18278
rect 2656 18214 2673 18278
rect 2737 18214 2754 18278
rect 2818 18214 2835 18278
rect 2899 18214 2916 18278
rect 2980 18214 2997 18278
rect 3061 18214 3078 18278
rect 3142 18214 3159 18278
rect 3223 18214 3240 18278
rect 3304 18214 3321 18278
rect 3385 18214 3402 18278
rect 3466 18214 3483 18278
rect 3547 18214 3563 18278
rect 3627 18214 3643 18278
rect 3707 18214 3723 18278
rect 3787 18214 3803 18278
rect 3867 18214 3883 18278
rect 3947 18244 4016 18278
rect 4080 18244 4129 18308
rect 4193 18244 4242 18308
rect 4306 18244 4355 18308
rect 4419 18297 4457 18308
tri 4457 18297 4674 18514 sw
tri 10338 18297 10555 18514 se
rect 10555 18512 11065 18514
rect 10555 18448 10593 18512
rect 10657 18448 10706 18512
rect 10770 18448 10819 18512
rect 10883 18448 10932 18512
rect 10996 18466 11065 18512
rect 11129 18466 11145 18530
rect 11209 18466 11225 18530
rect 11289 18466 11305 18530
rect 11369 18466 11385 18530
rect 11449 18466 11465 18530
rect 11529 18466 11546 18530
rect 11610 18466 11627 18530
rect 11691 18466 11708 18530
rect 11772 18466 11789 18530
rect 11853 18466 11870 18530
rect 11934 18466 11951 18530
rect 12015 18466 12032 18530
rect 12096 18466 12113 18530
rect 12177 18466 12194 18530
rect 12258 18466 12275 18530
rect 12339 18466 12356 18530
rect 12420 18466 12437 18530
rect 12501 18466 12518 18530
rect 12582 18466 12599 18530
rect 12663 18466 12680 18530
rect 12744 18466 12761 18530
rect 12825 18466 12842 18530
rect 12906 18466 12923 18530
rect 12987 18466 13004 18530
rect 13068 18466 13085 18530
rect 13149 18466 13166 18530
rect 13230 18466 13247 18530
rect 13311 18466 13328 18530
rect 13392 18466 13409 18530
rect 13473 18466 13490 18530
rect 13554 18466 13571 18530
rect 13635 18466 13652 18530
rect 13716 18466 13733 18530
rect 13797 18466 13814 18530
rect 13878 18466 13895 18530
rect 13959 18466 13976 18530
rect 14040 18466 14057 18530
rect 14121 18466 14138 18530
rect 14202 18466 14219 18530
rect 14283 18466 14300 18530
rect 14364 18466 14381 18530
rect 14445 18466 14462 18530
rect 14526 18466 14543 18530
rect 14607 18466 14624 18530
rect 14688 18466 14705 18530
rect 14769 18466 14786 18530
rect 14850 18466 14858 18530
rect 10996 18448 14858 18466
rect 10555 18446 14858 18448
rect 10555 18410 11065 18446
rect 10555 18346 10593 18410
rect 10657 18346 10706 18410
rect 10770 18346 10819 18410
rect 10883 18346 10932 18410
rect 10996 18382 11065 18410
rect 11129 18382 11145 18446
rect 11209 18382 11225 18446
rect 11289 18382 11305 18446
rect 11369 18382 11385 18446
rect 11449 18382 11465 18446
rect 11529 18382 11546 18446
rect 11610 18382 11627 18446
rect 11691 18382 11708 18446
rect 11772 18382 11789 18446
rect 11853 18382 11870 18446
rect 11934 18382 11951 18446
rect 12015 18382 12032 18446
rect 12096 18382 12113 18446
rect 12177 18382 12194 18446
rect 12258 18382 12275 18446
rect 12339 18382 12356 18446
rect 12420 18382 12437 18446
rect 12501 18382 12518 18446
rect 12582 18382 12599 18446
rect 12663 18382 12680 18446
rect 12744 18382 12761 18446
rect 12825 18382 12842 18446
rect 12906 18382 12923 18446
rect 12987 18382 13004 18446
rect 13068 18382 13085 18446
rect 13149 18382 13166 18446
rect 13230 18382 13247 18446
rect 13311 18382 13328 18446
rect 13392 18382 13409 18446
rect 13473 18382 13490 18446
rect 13554 18382 13571 18446
rect 13635 18382 13652 18446
rect 13716 18382 13733 18446
rect 13797 18382 13814 18446
rect 13878 18382 13895 18446
rect 13959 18382 13976 18446
rect 14040 18382 14057 18446
rect 14121 18382 14138 18446
rect 14202 18382 14219 18446
rect 14283 18382 14300 18446
rect 14364 18382 14381 18446
rect 14445 18382 14462 18446
rect 14526 18382 14543 18446
rect 14607 18382 14624 18446
rect 14688 18382 14705 18446
rect 14769 18382 14786 18446
rect 14850 18382 14858 18446
rect 10996 18362 14858 18382
rect 10996 18346 11065 18362
rect 10555 18308 11065 18346
rect 10555 18297 10593 18308
rect 4419 18244 4478 18297
rect 3947 18233 4478 18244
rect 4542 18233 4598 18297
rect 4662 18233 4674 18297
rect 3947 18214 4674 18233
rect 99 18206 4674 18214
rect 99 18194 4016 18206
rect 99 18130 162 18194
rect 226 18130 243 18194
rect 307 18130 324 18194
rect 388 18130 405 18194
rect 469 18130 486 18194
rect 550 18130 567 18194
rect 631 18130 648 18194
rect 712 18130 729 18194
rect 793 18130 810 18194
rect 874 18130 891 18194
rect 955 18130 972 18194
rect 1036 18130 1053 18194
rect 1117 18130 1134 18194
rect 1198 18130 1215 18194
rect 1279 18130 1296 18194
rect 1360 18130 1377 18194
rect 1441 18130 1458 18194
rect 1522 18130 1539 18194
rect 1603 18130 1620 18194
rect 1684 18130 1701 18194
rect 1765 18130 1782 18194
rect 1846 18130 1863 18194
rect 1927 18130 1944 18194
rect 2008 18130 2025 18194
rect 2089 18130 2106 18194
rect 2170 18130 2187 18194
rect 2251 18130 2268 18194
rect 2332 18130 2349 18194
rect 2413 18130 2430 18194
rect 2494 18130 2511 18194
rect 2575 18130 2592 18194
rect 2656 18130 2673 18194
rect 2737 18130 2754 18194
rect 2818 18130 2835 18194
rect 2899 18130 2916 18194
rect 2980 18130 2997 18194
rect 3061 18130 3078 18194
rect 3142 18130 3159 18194
rect 3223 18130 3240 18194
rect 3304 18130 3321 18194
rect 3385 18130 3402 18194
rect 3466 18130 3483 18194
rect 3547 18130 3563 18194
rect 3627 18130 3643 18194
rect 3707 18130 3723 18194
rect 3787 18130 3803 18194
rect 3867 18130 3883 18194
rect 3947 18142 4016 18194
rect 4080 18142 4129 18206
rect 4193 18142 4242 18206
rect 4306 18142 4355 18206
rect 4419 18183 4674 18206
rect 4419 18142 4478 18183
rect 3947 18130 4478 18142
rect 99 18119 4478 18130
rect 4542 18119 4598 18183
rect 4662 18119 4674 18183
tri 4674 18119 4852 18297 sw
tri 10160 18119 10338 18297 se
rect 10338 18233 10350 18297
rect 10414 18233 10470 18297
rect 10534 18244 10593 18297
rect 10657 18244 10706 18308
rect 10770 18244 10819 18308
rect 10883 18244 10932 18308
rect 10996 18298 11065 18308
rect 11129 18298 11145 18362
rect 11209 18298 11225 18362
rect 11289 18298 11305 18362
rect 11369 18298 11385 18362
rect 11449 18298 11465 18362
rect 11529 18298 11546 18362
rect 11610 18298 11627 18362
rect 11691 18298 11708 18362
rect 11772 18298 11789 18362
rect 11853 18298 11870 18362
rect 11934 18298 11951 18362
rect 12015 18298 12032 18362
rect 12096 18298 12113 18362
rect 12177 18298 12194 18362
rect 12258 18298 12275 18362
rect 12339 18298 12356 18362
rect 12420 18298 12437 18362
rect 12501 18298 12518 18362
rect 12582 18298 12599 18362
rect 12663 18298 12680 18362
rect 12744 18298 12761 18362
rect 12825 18298 12842 18362
rect 12906 18298 12923 18362
rect 12987 18298 13004 18362
rect 13068 18298 13085 18362
rect 13149 18298 13166 18362
rect 13230 18298 13247 18362
rect 13311 18298 13328 18362
rect 13392 18298 13409 18362
rect 13473 18298 13490 18362
rect 13554 18298 13571 18362
rect 13635 18298 13652 18362
rect 13716 18298 13733 18362
rect 13797 18298 13814 18362
rect 13878 18298 13895 18362
rect 13959 18298 13976 18362
rect 14040 18298 14057 18362
rect 14121 18298 14138 18362
rect 14202 18298 14219 18362
rect 14283 18298 14300 18362
rect 14364 18298 14381 18362
rect 14445 18298 14462 18362
rect 14526 18298 14543 18362
rect 14607 18298 14624 18362
rect 14688 18298 14705 18362
rect 14769 18298 14786 18362
rect 14850 18298 14858 18362
rect 10996 18278 14858 18298
rect 10996 18244 11065 18278
rect 10534 18233 11065 18244
rect 10338 18214 11065 18233
rect 11129 18214 11145 18278
rect 11209 18214 11225 18278
rect 11289 18214 11305 18278
rect 11369 18214 11385 18278
rect 11449 18214 11465 18278
rect 11529 18214 11546 18278
rect 11610 18214 11627 18278
rect 11691 18214 11708 18278
rect 11772 18214 11789 18278
rect 11853 18214 11870 18278
rect 11934 18214 11951 18278
rect 12015 18214 12032 18278
rect 12096 18214 12113 18278
rect 12177 18214 12194 18278
rect 12258 18214 12275 18278
rect 12339 18214 12356 18278
rect 12420 18214 12437 18278
rect 12501 18214 12518 18278
rect 12582 18214 12599 18278
rect 12663 18214 12680 18278
rect 12744 18214 12761 18278
rect 12825 18214 12842 18278
rect 12906 18214 12923 18278
rect 12987 18214 13004 18278
rect 13068 18214 13085 18278
rect 13149 18214 13166 18278
rect 13230 18214 13247 18278
rect 13311 18214 13328 18278
rect 13392 18214 13409 18278
rect 13473 18214 13490 18278
rect 13554 18214 13571 18278
rect 13635 18214 13652 18278
rect 13716 18214 13733 18278
rect 13797 18214 13814 18278
rect 13878 18214 13895 18278
rect 13959 18214 13976 18278
rect 14040 18214 14057 18278
rect 14121 18214 14138 18278
rect 14202 18214 14219 18278
rect 14283 18214 14300 18278
rect 14364 18214 14381 18278
rect 14445 18214 14462 18278
rect 14526 18214 14543 18278
rect 14607 18214 14624 18278
rect 14688 18214 14705 18278
rect 14769 18214 14786 18278
rect 14850 18214 14858 18278
rect 10338 18206 14858 18214
rect 10338 18183 10593 18206
rect 10338 18119 10350 18183
rect 10414 18119 10470 18183
rect 10534 18142 10593 18183
rect 10657 18142 10706 18206
rect 10770 18142 10819 18206
rect 10883 18142 10932 18206
rect 10996 18194 14858 18206
rect 10996 18142 11065 18194
rect 10534 18130 11065 18142
rect 11129 18130 11145 18194
rect 11209 18130 11225 18194
rect 11289 18130 11305 18194
rect 11369 18130 11385 18194
rect 11449 18130 11465 18194
rect 11529 18130 11546 18194
rect 11610 18130 11627 18194
rect 11691 18130 11708 18194
rect 11772 18130 11789 18194
rect 11853 18130 11870 18194
rect 11934 18130 11951 18194
rect 12015 18130 12032 18194
rect 12096 18130 12113 18194
rect 12177 18130 12194 18194
rect 12258 18130 12275 18194
rect 12339 18130 12356 18194
rect 12420 18130 12437 18194
rect 12501 18130 12518 18194
rect 12582 18130 12599 18194
rect 12663 18130 12680 18194
rect 12744 18130 12761 18194
rect 12825 18130 12842 18194
rect 12906 18130 12923 18194
rect 12987 18130 13004 18194
rect 13068 18130 13085 18194
rect 13149 18130 13166 18194
rect 13230 18130 13247 18194
rect 13311 18130 13328 18194
rect 13392 18130 13409 18194
rect 13473 18130 13490 18194
rect 13554 18130 13571 18194
rect 13635 18130 13652 18194
rect 13716 18130 13733 18194
rect 13797 18130 13814 18194
rect 13878 18130 13895 18194
rect 13959 18130 13976 18194
rect 14040 18130 14057 18194
rect 14121 18130 14138 18194
rect 14202 18130 14219 18194
rect 14283 18130 14300 18194
rect 14364 18130 14381 18194
rect 14445 18130 14462 18194
rect 14526 18130 14543 18194
rect 14607 18130 14624 18194
rect 14688 18130 14705 18194
rect 14769 18130 14786 18194
rect 14850 18130 14858 18194
rect 10534 18119 14858 18130
rect 99 18092 4852 18119
tri 4852 18092 4879 18119 sw
tri 10133 18092 10160 18119 se
rect 10160 18092 14858 18119
rect 99 18086 4879 18092
rect 99 14742 137 18086
rect 4841 14742 4879 18086
tri 10125 18084 10133 18092 se
rect 10133 18086 14858 18092
rect 10133 18084 10143 18086
rect 99 14725 4879 14742
rect 99 14661 137 14725
rect 201 14661 217 14725
rect 281 14661 297 14725
rect 361 14661 377 14725
rect 441 14661 457 14725
rect 521 14661 537 14725
rect 601 14661 617 14725
rect 681 14661 697 14725
rect 761 14661 777 14725
rect 841 14661 857 14725
rect 921 14661 937 14725
rect 1001 14661 1017 14725
rect 1081 14661 1097 14725
rect 1161 14661 1177 14725
rect 1241 14661 1257 14725
rect 1321 14661 1337 14725
rect 1401 14661 1417 14725
rect 1481 14661 1497 14725
rect 1561 14661 1577 14725
rect 1641 14661 1657 14725
rect 1721 14661 1737 14725
rect 1801 14661 1817 14725
rect 1881 14661 1897 14725
rect 1961 14661 1977 14725
rect 2041 14661 2057 14725
rect 2121 14661 2137 14725
rect 2201 14661 2217 14725
rect 2281 14661 2297 14725
rect 2361 14661 2377 14725
rect 2441 14661 2457 14725
rect 2521 14661 2537 14725
rect 2601 14661 2617 14725
rect 2681 14661 2697 14725
rect 2761 14661 2777 14725
rect 2841 14661 2857 14725
rect 2921 14661 2937 14725
rect 3001 14661 3017 14725
rect 3081 14661 3097 14725
rect 3161 14661 3177 14725
rect 3241 14661 3257 14725
rect 3321 14661 3337 14725
rect 3401 14661 3417 14725
rect 3481 14661 3497 14725
rect 3561 14661 3577 14725
rect 3641 14661 3657 14725
rect 3721 14661 3737 14725
rect 3801 14661 3817 14725
rect 3881 14661 3897 14725
rect 3961 14661 3977 14725
rect 4041 14661 4057 14725
rect 4121 14661 4137 14725
rect 4201 14661 4217 14725
rect 4281 14661 4297 14725
rect 4361 14661 4377 14725
rect 4441 14661 4457 14725
rect 4521 14661 4537 14725
rect 4601 14661 4617 14725
rect 4681 14661 4697 14725
rect 4761 14661 4777 14725
rect 4841 14661 4879 14725
rect 99 14644 4879 14661
rect 99 14580 137 14644
rect 201 14580 217 14644
rect 281 14580 297 14644
rect 361 14580 377 14644
rect 441 14580 457 14644
rect 521 14580 537 14644
rect 601 14580 617 14644
rect 681 14580 697 14644
rect 761 14580 777 14644
rect 841 14580 857 14644
rect 921 14580 937 14644
rect 1001 14580 1017 14644
rect 1081 14580 1097 14644
rect 1161 14580 1177 14644
rect 1241 14580 1257 14644
rect 1321 14580 1337 14644
rect 1401 14580 1417 14644
rect 1481 14580 1497 14644
rect 1561 14580 1577 14644
rect 1641 14580 1657 14644
rect 1721 14580 1737 14644
rect 1801 14580 1817 14644
rect 1881 14580 1897 14644
rect 1961 14580 1977 14644
rect 2041 14580 2057 14644
rect 2121 14580 2137 14644
rect 2201 14580 2217 14644
rect 2281 14580 2297 14644
rect 2361 14580 2377 14644
rect 2441 14580 2457 14644
rect 2521 14580 2537 14644
rect 2601 14580 2617 14644
rect 2681 14580 2697 14644
rect 2761 14580 2777 14644
rect 2841 14580 2857 14644
rect 2921 14580 2937 14644
rect 3001 14580 3017 14644
rect 3081 14580 3097 14644
rect 3161 14580 3177 14644
rect 3241 14580 3257 14644
rect 3321 14580 3337 14644
rect 3401 14580 3417 14644
rect 3481 14580 3497 14644
rect 3561 14580 3577 14644
rect 3641 14580 3657 14644
rect 3721 14580 3737 14644
rect 3801 14580 3817 14644
rect 3881 14580 3897 14644
rect 3961 14580 3977 14644
rect 4041 14580 4057 14644
rect 4121 14580 4137 14644
rect 4201 14580 4217 14644
rect 4281 14580 4297 14644
rect 4361 14580 4377 14644
rect 4441 14580 4457 14644
rect 4521 14580 4537 14644
rect 4601 14580 4617 14644
rect 4681 14580 4697 14644
rect 4761 14580 4777 14644
rect 4841 14580 4879 14644
rect 99 14563 4879 14580
rect 99 14499 137 14563
rect 201 14499 217 14563
rect 281 14499 297 14563
rect 361 14499 377 14563
rect 441 14499 457 14563
rect 521 14499 537 14563
rect 601 14499 617 14563
rect 681 14499 697 14563
rect 761 14499 777 14563
rect 841 14499 857 14563
rect 921 14499 937 14563
rect 1001 14499 1017 14563
rect 1081 14499 1097 14563
rect 1161 14499 1177 14563
rect 1241 14499 1257 14563
rect 1321 14499 1337 14563
rect 1401 14499 1417 14563
rect 1481 14499 1497 14563
rect 1561 14499 1577 14563
rect 1641 14499 1657 14563
rect 1721 14499 1737 14563
rect 1801 14499 1817 14563
rect 1881 14499 1897 14563
rect 1961 14499 1977 14563
rect 2041 14499 2057 14563
rect 2121 14499 2137 14563
rect 2201 14499 2217 14563
rect 2281 14499 2297 14563
rect 2361 14499 2377 14563
rect 2441 14499 2457 14563
rect 2521 14499 2537 14563
rect 2601 14499 2617 14563
rect 2681 14499 2697 14563
rect 2761 14499 2777 14563
rect 2841 14499 2857 14563
rect 2921 14499 2937 14563
rect 3001 14499 3017 14563
rect 3081 14499 3097 14563
rect 3161 14499 3177 14563
rect 3241 14499 3257 14563
rect 3321 14499 3337 14563
rect 3401 14499 3417 14563
rect 3481 14499 3497 14563
rect 3561 14499 3577 14563
rect 3641 14499 3657 14563
rect 3721 14499 3737 14563
rect 3801 14499 3817 14563
rect 3881 14499 3897 14563
rect 3961 14499 3977 14563
rect 4041 14499 4057 14563
rect 4121 14499 4137 14563
rect 4201 14499 4217 14563
rect 4281 14499 4297 14563
rect 4361 14499 4377 14563
rect 4441 14499 4457 14563
rect 4521 14499 4537 14563
rect 4601 14499 4617 14563
rect 4681 14499 4697 14563
rect 4761 14499 4777 14563
rect 4841 14499 4879 14563
rect 99 14482 4879 14499
rect 99 14418 137 14482
rect 201 14418 217 14482
rect 281 14418 297 14482
rect 361 14418 377 14482
rect 441 14418 457 14482
rect 521 14418 537 14482
rect 601 14418 617 14482
rect 681 14418 697 14482
rect 761 14418 777 14482
rect 841 14418 857 14482
rect 921 14418 937 14482
rect 1001 14418 1017 14482
rect 1081 14418 1097 14482
rect 1161 14418 1177 14482
rect 1241 14418 1257 14482
rect 1321 14418 1337 14482
rect 1401 14418 1417 14482
rect 1481 14418 1497 14482
rect 1561 14418 1577 14482
rect 1641 14418 1657 14482
rect 1721 14418 1737 14482
rect 1801 14418 1817 14482
rect 1881 14418 1897 14482
rect 1961 14418 1977 14482
rect 2041 14418 2057 14482
rect 2121 14418 2137 14482
rect 2201 14418 2217 14482
rect 2281 14418 2297 14482
rect 2361 14418 2377 14482
rect 2441 14418 2457 14482
rect 2521 14418 2537 14482
rect 2601 14418 2617 14482
rect 2681 14418 2697 14482
rect 2761 14418 2777 14482
rect 2841 14418 2857 14482
rect 2921 14418 2937 14482
rect 3001 14418 3017 14482
rect 3081 14418 3097 14482
rect 3161 14418 3177 14482
rect 3241 14418 3257 14482
rect 3321 14418 3337 14482
rect 3401 14418 3417 14482
rect 3481 14418 3497 14482
rect 3561 14418 3577 14482
rect 3641 14418 3657 14482
rect 3721 14418 3737 14482
rect 3801 14418 3817 14482
rect 3881 14418 3897 14482
rect 3961 14418 3977 14482
rect 4041 14418 4057 14482
rect 4121 14418 4137 14482
rect 4201 14418 4217 14482
rect 4281 14418 4297 14482
rect 4361 14418 4377 14482
rect 4441 14418 4457 14482
rect 4521 14418 4537 14482
rect 4601 14418 4617 14482
rect 4681 14418 4697 14482
rect 4761 14418 4777 14482
rect 4841 14418 4879 14482
rect 99 14401 4879 14418
rect 99 14337 137 14401
rect 201 14337 217 14401
rect 281 14337 297 14401
rect 361 14337 377 14401
rect 441 14337 457 14401
rect 521 14337 537 14401
rect 601 14337 617 14401
rect 681 14337 697 14401
rect 761 14337 777 14401
rect 841 14337 857 14401
rect 921 14337 937 14401
rect 1001 14337 1017 14401
rect 1081 14337 1097 14401
rect 1161 14337 1177 14401
rect 1241 14337 1257 14401
rect 1321 14337 1337 14401
rect 1401 14337 1417 14401
rect 1481 14337 1497 14401
rect 1561 14337 1577 14401
rect 1641 14337 1657 14401
rect 1721 14337 1737 14401
rect 1801 14337 1817 14401
rect 1881 14337 1897 14401
rect 1961 14337 1977 14401
rect 2041 14337 2057 14401
rect 2121 14337 2137 14401
rect 2201 14337 2217 14401
rect 2281 14337 2297 14401
rect 2361 14337 2377 14401
rect 2441 14337 2457 14401
rect 2521 14337 2537 14401
rect 2601 14337 2617 14401
rect 2681 14337 2697 14401
rect 2761 14337 2777 14401
rect 2841 14337 2857 14401
rect 2921 14337 2937 14401
rect 3001 14337 3017 14401
rect 3081 14337 3097 14401
rect 3161 14337 3177 14401
rect 3241 14337 3257 14401
rect 3321 14337 3337 14401
rect 3401 14337 3417 14401
rect 3481 14337 3497 14401
rect 3561 14337 3577 14401
rect 3641 14337 3657 14401
rect 3721 14337 3737 14401
rect 3801 14337 3817 14401
rect 3881 14337 3897 14401
rect 3961 14337 3977 14401
rect 4041 14337 4057 14401
rect 4121 14337 4137 14401
rect 4201 14337 4217 14401
rect 4281 14337 4297 14401
rect 4361 14337 4377 14401
rect 4441 14337 4457 14401
rect 4521 14337 4537 14401
rect 4601 14337 4617 14401
rect 4681 14337 4697 14401
rect 4761 14337 4777 14401
rect 4841 14337 4879 14401
rect 99 14320 4879 14337
rect 99 14256 137 14320
rect 201 14256 217 14320
rect 281 14256 297 14320
rect 361 14256 377 14320
rect 441 14256 457 14320
rect 521 14256 537 14320
rect 601 14256 617 14320
rect 681 14256 697 14320
rect 761 14256 777 14320
rect 841 14256 857 14320
rect 921 14256 937 14320
rect 1001 14256 1017 14320
rect 1081 14256 1097 14320
rect 1161 14256 1177 14320
rect 1241 14256 1257 14320
rect 1321 14256 1337 14320
rect 1401 14256 1417 14320
rect 1481 14256 1497 14320
rect 1561 14256 1577 14320
rect 1641 14256 1657 14320
rect 1721 14256 1737 14320
rect 1801 14256 1817 14320
rect 1881 14256 1897 14320
rect 1961 14256 1977 14320
rect 2041 14256 2057 14320
rect 2121 14256 2137 14320
rect 2201 14256 2217 14320
rect 2281 14256 2297 14320
rect 2361 14256 2377 14320
rect 2441 14256 2457 14320
rect 2521 14256 2537 14320
rect 2601 14256 2617 14320
rect 2681 14256 2697 14320
rect 2761 14256 2777 14320
rect 2841 14256 2857 14320
rect 2921 14256 2937 14320
rect 3001 14256 3017 14320
rect 3081 14256 3097 14320
rect 3161 14256 3177 14320
rect 3241 14256 3257 14320
rect 3321 14256 3337 14320
rect 3401 14256 3417 14320
rect 3481 14256 3497 14320
rect 3561 14256 3577 14320
rect 3641 14256 3657 14320
rect 3721 14256 3737 14320
rect 3801 14256 3817 14320
rect 3881 14256 3897 14320
rect 3961 14256 3977 14320
rect 4041 14256 4057 14320
rect 4121 14256 4137 14320
rect 4201 14256 4217 14320
rect 4281 14256 4297 14320
rect 4361 14256 4377 14320
rect 4441 14256 4457 14320
rect 4521 14256 4537 14320
rect 4601 14256 4617 14320
rect 4681 14256 4697 14320
rect 4761 14256 4777 14320
rect 4841 14256 4879 14320
rect 99 14239 4879 14256
rect 99 14175 137 14239
rect 201 14175 217 14239
rect 281 14175 297 14239
rect 361 14175 377 14239
rect 441 14175 457 14239
rect 521 14175 537 14239
rect 601 14175 617 14239
rect 681 14175 697 14239
rect 761 14175 777 14239
rect 841 14175 857 14239
rect 921 14175 937 14239
rect 1001 14175 1017 14239
rect 1081 14175 1097 14239
rect 1161 14175 1177 14239
rect 1241 14175 1257 14239
rect 1321 14175 1337 14239
rect 1401 14175 1417 14239
rect 1481 14175 1497 14239
rect 1561 14175 1577 14239
rect 1641 14175 1657 14239
rect 1721 14175 1737 14239
rect 1801 14175 1817 14239
rect 1881 14175 1897 14239
rect 1961 14175 1977 14239
rect 2041 14175 2057 14239
rect 2121 14175 2137 14239
rect 2201 14175 2217 14239
rect 2281 14175 2297 14239
rect 2361 14175 2377 14239
rect 2441 14175 2457 14239
rect 2521 14175 2537 14239
rect 2601 14175 2617 14239
rect 2681 14175 2697 14239
rect 2761 14175 2777 14239
rect 2841 14175 2857 14239
rect 2921 14175 2937 14239
rect 3001 14175 3017 14239
rect 3081 14175 3097 14239
rect 3161 14175 3177 14239
rect 3241 14175 3257 14239
rect 3321 14175 3337 14239
rect 3401 14175 3417 14239
rect 3481 14175 3497 14239
rect 3561 14175 3577 14239
rect 3641 14175 3657 14239
rect 3721 14175 3737 14239
rect 3801 14175 3817 14239
rect 3881 14175 3897 14239
rect 3961 14175 3977 14239
rect 4041 14175 4057 14239
rect 4121 14175 4137 14239
rect 4201 14175 4217 14239
rect 4281 14175 4297 14239
rect 4361 14175 4377 14239
rect 4441 14175 4457 14239
rect 4521 14175 4537 14239
rect 4601 14175 4617 14239
rect 4681 14175 4697 14239
rect 4761 14175 4777 14239
rect 4841 14175 4879 14239
rect 99 14158 4879 14175
rect 99 14094 137 14158
rect 201 14094 217 14158
rect 281 14094 297 14158
rect 361 14094 377 14158
rect 441 14094 457 14158
rect 521 14094 537 14158
rect 601 14094 617 14158
rect 681 14094 697 14158
rect 761 14094 777 14158
rect 841 14094 857 14158
rect 921 14094 937 14158
rect 1001 14094 1017 14158
rect 1081 14094 1097 14158
rect 1161 14094 1177 14158
rect 1241 14094 1257 14158
rect 1321 14094 1337 14158
rect 1401 14094 1417 14158
rect 1481 14094 1497 14158
rect 1561 14094 1577 14158
rect 1641 14094 1657 14158
rect 1721 14094 1737 14158
rect 1801 14094 1817 14158
rect 1881 14094 1897 14158
rect 1961 14094 1977 14158
rect 2041 14094 2057 14158
rect 2121 14094 2137 14158
rect 2201 14094 2217 14158
rect 2281 14094 2297 14158
rect 2361 14094 2377 14158
rect 2441 14094 2457 14158
rect 2521 14094 2537 14158
rect 2601 14094 2617 14158
rect 2681 14094 2697 14158
rect 2761 14094 2777 14158
rect 2841 14094 2857 14158
rect 2921 14094 2937 14158
rect 3001 14094 3017 14158
rect 3081 14094 3097 14158
rect 3161 14094 3177 14158
rect 3241 14094 3257 14158
rect 3321 14094 3337 14158
rect 3401 14094 3417 14158
rect 3481 14094 3497 14158
rect 3561 14094 3577 14158
rect 3641 14094 3657 14158
rect 3721 14094 3737 14158
rect 3801 14094 3817 14158
rect 3881 14094 3897 14158
rect 3961 14094 3977 14158
rect 4041 14094 4057 14158
rect 4121 14094 4137 14158
rect 4201 14094 4217 14158
rect 4281 14094 4297 14158
rect 4361 14094 4377 14158
rect 4441 14094 4457 14158
rect 4521 14094 4537 14158
rect 4601 14094 4617 14158
rect 4681 14094 4697 14158
rect 4761 14094 4777 14158
rect 4841 14094 4879 14158
rect 99 14077 4879 14094
rect 99 14013 137 14077
rect 201 14013 217 14077
rect 281 14013 297 14077
rect 361 14013 377 14077
rect 441 14013 457 14077
rect 521 14013 537 14077
rect 601 14013 617 14077
rect 681 14013 697 14077
rect 761 14013 777 14077
rect 841 14013 857 14077
rect 921 14013 937 14077
rect 1001 14013 1017 14077
rect 1081 14013 1097 14077
rect 1161 14013 1177 14077
rect 1241 14013 1257 14077
rect 1321 14013 1337 14077
rect 1401 14013 1417 14077
rect 1481 14013 1497 14077
rect 1561 14013 1577 14077
rect 1641 14013 1657 14077
rect 1721 14013 1737 14077
rect 1801 14013 1817 14077
rect 1881 14013 1897 14077
rect 1961 14013 1977 14077
rect 2041 14013 2057 14077
rect 2121 14013 2137 14077
rect 2201 14013 2217 14077
rect 2281 14013 2297 14077
rect 2361 14013 2377 14077
rect 2441 14013 2457 14077
rect 2521 14013 2537 14077
rect 2601 14013 2617 14077
rect 2681 14013 2697 14077
rect 2761 14013 2777 14077
rect 2841 14013 2857 14077
rect 2921 14013 2937 14077
rect 3001 14013 3017 14077
rect 3081 14013 3097 14077
rect 3161 14013 3177 14077
rect 3241 14013 3257 14077
rect 3321 14013 3337 14077
rect 3401 14013 3417 14077
rect 3481 14013 3497 14077
rect 3561 14013 3577 14077
rect 3641 14013 3657 14077
rect 3721 14013 3737 14077
rect 3801 14013 3817 14077
rect 3881 14013 3897 14077
rect 3961 14013 3977 14077
rect 4041 14013 4057 14077
rect 4121 14013 4137 14077
rect 4201 14013 4217 14077
rect 4281 14013 4297 14077
rect 4361 14013 4377 14077
rect 4441 14013 4457 14077
rect 4521 14013 4537 14077
rect 4601 14013 4617 14077
rect 4681 14013 4697 14077
rect 4761 14013 4777 14077
rect 4841 14013 4879 14077
rect 99 14007 4879 14013
tri 10078 18037 10125 18084 se
rect 10125 18037 10143 18084
rect 10078 14742 10143 18037
rect 14847 14742 14858 18086
rect 10078 14725 14858 14742
rect 10078 14661 10143 14725
rect 10207 14661 10223 14725
rect 10287 14661 10303 14725
rect 10367 14661 10383 14725
rect 10447 14661 10463 14725
rect 10527 14661 10543 14725
rect 10607 14661 10623 14725
rect 10687 14661 10703 14725
rect 10767 14661 10783 14725
rect 10847 14661 10863 14725
rect 10927 14661 10943 14725
rect 11007 14661 11023 14725
rect 11087 14661 11103 14725
rect 11167 14661 11183 14725
rect 11247 14661 11263 14725
rect 11327 14661 11343 14725
rect 11407 14661 11423 14725
rect 11487 14661 11503 14725
rect 11567 14661 11583 14725
rect 11647 14661 11663 14725
rect 11727 14661 11743 14725
rect 11807 14661 11823 14725
rect 11887 14661 11903 14725
rect 11967 14661 11983 14725
rect 12047 14661 12063 14725
rect 12127 14661 12143 14725
rect 12207 14661 12223 14725
rect 12287 14661 12303 14725
rect 12367 14661 12383 14725
rect 12447 14661 12463 14725
rect 12527 14661 12543 14725
rect 12607 14661 12623 14725
rect 12687 14661 12703 14725
rect 12767 14661 12783 14725
rect 12847 14661 12863 14725
rect 12927 14661 12943 14725
rect 13007 14661 13023 14725
rect 13087 14661 13103 14725
rect 13167 14661 13183 14725
rect 13247 14661 13263 14725
rect 13327 14661 13343 14725
rect 13407 14661 13423 14725
rect 13487 14661 13503 14725
rect 13567 14661 13583 14725
rect 13647 14661 13663 14725
rect 13727 14661 13743 14725
rect 13807 14661 13823 14725
rect 13887 14661 13903 14725
rect 13967 14661 13983 14725
rect 14047 14661 14063 14725
rect 14127 14661 14143 14725
rect 14207 14661 14223 14725
rect 14287 14661 14303 14725
rect 14367 14661 14383 14725
rect 14447 14661 14463 14725
rect 14527 14661 14543 14725
rect 14607 14661 14623 14725
rect 14687 14661 14703 14725
rect 14767 14661 14783 14725
rect 14847 14661 14858 14725
rect 10078 14644 14858 14661
rect 10078 14580 10143 14644
rect 10207 14580 10223 14644
rect 10287 14580 10303 14644
rect 10367 14580 10383 14644
rect 10447 14580 10463 14644
rect 10527 14580 10543 14644
rect 10607 14580 10623 14644
rect 10687 14580 10703 14644
rect 10767 14580 10783 14644
rect 10847 14580 10863 14644
rect 10927 14580 10943 14644
rect 11007 14580 11023 14644
rect 11087 14580 11103 14644
rect 11167 14580 11183 14644
rect 11247 14580 11263 14644
rect 11327 14580 11343 14644
rect 11407 14580 11423 14644
rect 11487 14580 11503 14644
rect 11567 14580 11583 14644
rect 11647 14580 11663 14644
rect 11727 14580 11743 14644
rect 11807 14580 11823 14644
rect 11887 14580 11903 14644
rect 11967 14580 11983 14644
rect 12047 14580 12063 14644
rect 12127 14580 12143 14644
rect 12207 14580 12223 14644
rect 12287 14580 12303 14644
rect 12367 14580 12383 14644
rect 12447 14580 12463 14644
rect 12527 14580 12543 14644
rect 12607 14580 12623 14644
rect 12687 14580 12703 14644
rect 12767 14580 12783 14644
rect 12847 14580 12863 14644
rect 12927 14580 12943 14644
rect 13007 14580 13023 14644
rect 13087 14580 13103 14644
rect 13167 14580 13183 14644
rect 13247 14580 13263 14644
rect 13327 14580 13343 14644
rect 13407 14580 13423 14644
rect 13487 14580 13503 14644
rect 13567 14580 13583 14644
rect 13647 14580 13663 14644
rect 13727 14580 13743 14644
rect 13807 14580 13823 14644
rect 13887 14580 13903 14644
rect 13967 14580 13983 14644
rect 14047 14580 14063 14644
rect 14127 14580 14143 14644
rect 14207 14580 14223 14644
rect 14287 14580 14303 14644
rect 14367 14580 14383 14644
rect 14447 14580 14463 14644
rect 14527 14580 14543 14644
rect 14607 14580 14623 14644
rect 14687 14580 14703 14644
rect 14767 14580 14783 14644
rect 14847 14580 14858 14644
rect 10078 14563 14858 14580
rect 10078 14499 10143 14563
rect 10207 14499 10223 14563
rect 10287 14499 10303 14563
rect 10367 14499 10383 14563
rect 10447 14499 10463 14563
rect 10527 14499 10543 14563
rect 10607 14499 10623 14563
rect 10687 14499 10703 14563
rect 10767 14499 10783 14563
rect 10847 14499 10863 14563
rect 10927 14499 10943 14563
rect 11007 14499 11023 14563
rect 11087 14499 11103 14563
rect 11167 14499 11183 14563
rect 11247 14499 11263 14563
rect 11327 14499 11343 14563
rect 11407 14499 11423 14563
rect 11487 14499 11503 14563
rect 11567 14499 11583 14563
rect 11647 14499 11663 14563
rect 11727 14499 11743 14563
rect 11807 14499 11823 14563
rect 11887 14499 11903 14563
rect 11967 14499 11983 14563
rect 12047 14499 12063 14563
rect 12127 14499 12143 14563
rect 12207 14499 12223 14563
rect 12287 14499 12303 14563
rect 12367 14499 12383 14563
rect 12447 14499 12463 14563
rect 12527 14499 12543 14563
rect 12607 14499 12623 14563
rect 12687 14499 12703 14563
rect 12767 14499 12783 14563
rect 12847 14499 12863 14563
rect 12927 14499 12943 14563
rect 13007 14499 13023 14563
rect 13087 14499 13103 14563
rect 13167 14499 13183 14563
rect 13247 14499 13263 14563
rect 13327 14499 13343 14563
rect 13407 14499 13423 14563
rect 13487 14499 13503 14563
rect 13567 14499 13583 14563
rect 13647 14499 13663 14563
rect 13727 14499 13743 14563
rect 13807 14499 13823 14563
rect 13887 14499 13903 14563
rect 13967 14499 13983 14563
rect 14047 14499 14063 14563
rect 14127 14499 14143 14563
rect 14207 14499 14223 14563
rect 14287 14499 14303 14563
rect 14367 14499 14383 14563
rect 14447 14499 14463 14563
rect 14527 14499 14543 14563
rect 14607 14499 14623 14563
rect 14687 14499 14703 14563
rect 14767 14499 14783 14563
rect 14847 14499 14858 14563
rect 10078 14482 14858 14499
rect 10078 14418 10143 14482
rect 10207 14418 10223 14482
rect 10287 14418 10303 14482
rect 10367 14418 10383 14482
rect 10447 14418 10463 14482
rect 10527 14418 10543 14482
rect 10607 14418 10623 14482
rect 10687 14418 10703 14482
rect 10767 14418 10783 14482
rect 10847 14418 10863 14482
rect 10927 14418 10943 14482
rect 11007 14418 11023 14482
rect 11087 14418 11103 14482
rect 11167 14418 11183 14482
rect 11247 14418 11263 14482
rect 11327 14418 11343 14482
rect 11407 14418 11423 14482
rect 11487 14418 11503 14482
rect 11567 14418 11583 14482
rect 11647 14418 11663 14482
rect 11727 14418 11743 14482
rect 11807 14418 11823 14482
rect 11887 14418 11903 14482
rect 11967 14418 11983 14482
rect 12047 14418 12063 14482
rect 12127 14418 12143 14482
rect 12207 14418 12223 14482
rect 12287 14418 12303 14482
rect 12367 14418 12383 14482
rect 12447 14418 12463 14482
rect 12527 14418 12543 14482
rect 12607 14418 12623 14482
rect 12687 14418 12703 14482
rect 12767 14418 12783 14482
rect 12847 14418 12863 14482
rect 12927 14418 12943 14482
rect 13007 14418 13023 14482
rect 13087 14418 13103 14482
rect 13167 14418 13183 14482
rect 13247 14418 13263 14482
rect 13327 14418 13343 14482
rect 13407 14418 13423 14482
rect 13487 14418 13503 14482
rect 13567 14418 13583 14482
rect 13647 14418 13663 14482
rect 13727 14418 13743 14482
rect 13807 14418 13823 14482
rect 13887 14418 13903 14482
rect 13967 14418 13983 14482
rect 14047 14418 14063 14482
rect 14127 14418 14143 14482
rect 14207 14418 14223 14482
rect 14287 14418 14303 14482
rect 14367 14418 14383 14482
rect 14447 14418 14463 14482
rect 14527 14418 14543 14482
rect 14607 14418 14623 14482
rect 14687 14418 14703 14482
rect 14767 14418 14783 14482
rect 14847 14418 14858 14482
rect 10078 14401 14858 14418
rect 10078 14337 10143 14401
rect 10207 14337 10223 14401
rect 10287 14337 10303 14401
rect 10367 14337 10383 14401
rect 10447 14337 10463 14401
rect 10527 14337 10543 14401
rect 10607 14337 10623 14401
rect 10687 14337 10703 14401
rect 10767 14337 10783 14401
rect 10847 14337 10863 14401
rect 10927 14337 10943 14401
rect 11007 14337 11023 14401
rect 11087 14337 11103 14401
rect 11167 14337 11183 14401
rect 11247 14337 11263 14401
rect 11327 14337 11343 14401
rect 11407 14337 11423 14401
rect 11487 14337 11503 14401
rect 11567 14337 11583 14401
rect 11647 14337 11663 14401
rect 11727 14337 11743 14401
rect 11807 14337 11823 14401
rect 11887 14337 11903 14401
rect 11967 14337 11983 14401
rect 12047 14337 12063 14401
rect 12127 14337 12143 14401
rect 12207 14337 12223 14401
rect 12287 14337 12303 14401
rect 12367 14337 12383 14401
rect 12447 14337 12463 14401
rect 12527 14337 12543 14401
rect 12607 14337 12623 14401
rect 12687 14337 12703 14401
rect 12767 14337 12783 14401
rect 12847 14337 12863 14401
rect 12927 14337 12943 14401
rect 13007 14337 13023 14401
rect 13087 14337 13103 14401
rect 13167 14337 13183 14401
rect 13247 14337 13263 14401
rect 13327 14337 13343 14401
rect 13407 14337 13423 14401
rect 13487 14337 13503 14401
rect 13567 14337 13583 14401
rect 13647 14337 13663 14401
rect 13727 14337 13743 14401
rect 13807 14337 13823 14401
rect 13887 14337 13903 14401
rect 13967 14337 13983 14401
rect 14047 14337 14063 14401
rect 14127 14337 14143 14401
rect 14207 14337 14223 14401
rect 14287 14337 14303 14401
rect 14367 14337 14383 14401
rect 14447 14337 14463 14401
rect 14527 14337 14543 14401
rect 14607 14337 14623 14401
rect 14687 14337 14703 14401
rect 14767 14337 14783 14401
rect 14847 14337 14858 14401
rect 10078 14320 14858 14337
rect 10078 14256 10143 14320
rect 10207 14256 10223 14320
rect 10287 14256 10303 14320
rect 10367 14256 10383 14320
rect 10447 14256 10463 14320
rect 10527 14256 10543 14320
rect 10607 14256 10623 14320
rect 10687 14256 10703 14320
rect 10767 14256 10783 14320
rect 10847 14256 10863 14320
rect 10927 14256 10943 14320
rect 11007 14256 11023 14320
rect 11087 14256 11103 14320
rect 11167 14256 11183 14320
rect 11247 14256 11263 14320
rect 11327 14256 11343 14320
rect 11407 14256 11423 14320
rect 11487 14256 11503 14320
rect 11567 14256 11583 14320
rect 11647 14256 11663 14320
rect 11727 14256 11743 14320
rect 11807 14256 11823 14320
rect 11887 14256 11903 14320
rect 11967 14256 11983 14320
rect 12047 14256 12063 14320
rect 12127 14256 12143 14320
rect 12207 14256 12223 14320
rect 12287 14256 12303 14320
rect 12367 14256 12383 14320
rect 12447 14256 12463 14320
rect 12527 14256 12543 14320
rect 12607 14256 12623 14320
rect 12687 14256 12703 14320
rect 12767 14256 12783 14320
rect 12847 14256 12863 14320
rect 12927 14256 12943 14320
rect 13007 14256 13023 14320
rect 13087 14256 13103 14320
rect 13167 14256 13183 14320
rect 13247 14256 13263 14320
rect 13327 14256 13343 14320
rect 13407 14256 13423 14320
rect 13487 14256 13503 14320
rect 13567 14256 13583 14320
rect 13647 14256 13663 14320
rect 13727 14256 13743 14320
rect 13807 14256 13823 14320
rect 13887 14256 13903 14320
rect 13967 14256 13983 14320
rect 14047 14256 14063 14320
rect 14127 14256 14143 14320
rect 14207 14256 14223 14320
rect 14287 14256 14303 14320
rect 14367 14256 14383 14320
rect 14447 14256 14463 14320
rect 14527 14256 14543 14320
rect 14607 14256 14623 14320
rect 14687 14256 14703 14320
rect 14767 14256 14783 14320
rect 14847 14256 14858 14320
rect 10078 14239 14858 14256
rect 10078 14175 10143 14239
rect 10207 14175 10223 14239
rect 10287 14175 10303 14239
rect 10367 14175 10383 14239
rect 10447 14175 10463 14239
rect 10527 14175 10543 14239
rect 10607 14175 10623 14239
rect 10687 14175 10703 14239
rect 10767 14175 10783 14239
rect 10847 14175 10863 14239
rect 10927 14175 10943 14239
rect 11007 14175 11023 14239
rect 11087 14175 11103 14239
rect 11167 14175 11183 14239
rect 11247 14175 11263 14239
rect 11327 14175 11343 14239
rect 11407 14175 11423 14239
rect 11487 14175 11503 14239
rect 11567 14175 11583 14239
rect 11647 14175 11663 14239
rect 11727 14175 11743 14239
rect 11807 14175 11823 14239
rect 11887 14175 11903 14239
rect 11967 14175 11983 14239
rect 12047 14175 12063 14239
rect 12127 14175 12143 14239
rect 12207 14175 12223 14239
rect 12287 14175 12303 14239
rect 12367 14175 12383 14239
rect 12447 14175 12463 14239
rect 12527 14175 12543 14239
rect 12607 14175 12623 14239
rect 12687 14175 12703 14239
rect 12767 14175 12783 14239
rect 12847 14175 12863 14239
rect 12927 14175 12943 14239
rect 13007 14175 13023 14239
rect 13087 14175 13103 14239
rect 13167 14175 13183 14239
rect 13247 14175 13263 14239
rect 13327 14175 13343 14239
rect 13407 14175 13423 14239
rect 13487 14175 13503 14239
rect 13567 14175 13583 14239
rect 13647 14175 13663 14239
rect 13727 14175 13743 14239
rect 13807 14175 13823 14239
rect 13887 14175 13903 14239
rect 13967 14175 13983 14239
rect 14047 14175 14063 14239
rect 14127 14175 14143 14239
rect 14207 14175 14223 14239
rect 14287 14175 14303 14239
rect 14367 14175 14383 14239
rect 14447 14175 14463 14239
rect 14527 14175 14543 14239
rect 14607 14175 14623 14239
rect 14687 14175 14703 14239
rect 14767 14175 14783 14239
rect 14847 14175 14858 14239
rect 10078 14158 14858 14175
rect 10078 14094 10143 14158
rect 10207 14094 10223 14158
rect 10287 14094 10303 14158
rect 10367 14094 10383 14158
rect 10447 14094 10463 14158
rect 10527 14094 10543 14158
rect 10607 14094 10623 14158
rect 10687 14094 10703 14158
rect 10767 14094 10783 14158
rect 10847 14094 10863 14158
rect 10927 14094 10943 14158
rect 11007 14094 11023 14158
rect 11087 14094 11103 14158
rect 11167 14094 11183 14158
rect 11247 14094 11263 14158
rect 11327 14094 11343 14158
rect 11407 14094 11423 14158
rect 11487 14094 11503 14158
rect 11567 14094 11583 14158
rect 11647 14094 11663 14158
rect 11727 14094 11743 14158
rect 11807 14094 11823 14158
rect 11887 14094 11903 14158
rect 11967 14094 11983 14158
rect 12047 14094 12063 14158
rect 12127 14094 12143 14158
rect 12207 14094 12223 14158
rect 12287 14094 12303 14158
rect 12367 14094 12383 14158
rect 12447 14094 12463 14158
rect 12527 14094 12543 14158
rect 12607 14094 12623 14158
rect 12687 14094 12703 14158
rect 12767 14094 12783 14158
rect 12847 14094 12863 14158
rect 12927 14094 12943 14158
rect 13007 14094 13023 14158
rect 13087 14094 13103 14158
rect 13167 14094 13183 14158
rect 13247 14094 13263 14158
rect 13327 14094 13343 14158
rect 13407 14094 13423 14158
rect 13487 14094 13503 14158
rect 13567 14094 13583 14158
rect 13647 14094 13663 14158
rect 13727 14094 13743 14158
rect 13807 14094 13823 14158
rect 13887 14094 13903 14158
rect 13967 14094 13983 14158
rect 14047 14094 14063 14158
rect 14127 14094 14143 14158
rect 14207 14094 14223 14158
rect 14287 14094 14303 14158
rect 14367 14094 14383 14158
rect 14447 14094 14463 14158
rect 14527 14094 14543 14158
rect 14607 14094 14623 14158
rect 14687 14094 14703 14158
rect 14767 14094 14783 14158
rect 14847 14094 14858 14158
rect 10078 14077 14858 14094
rect 10078 14013 10143 14077
rect 10207 14013 10223 14077
rect 10287 14013 10303 14077
rect 10367 14013 10383 14077
rect 10447 14013 10463 14077
rect 10527 14013 10543 14077
rect 10607 14013 10623 14077
rect 10687 14013 10703 14077
rect 10767 14013 10783 14077
rect 10847 14013 10863 14077
rect 10927 14013 10943 14077
rect 11007 14013 11023 14077
rect 11087 14013 11103 14077
rect 11167 14013 11183 14077
rect 11247 14013 11263 14077
rect 11327 14013 11343 14077
rect 11407 14013 11423 14077
rect 11487 14013 11503 14077
rect 11567 14013 11583 14077
rect 11647 14013 11663 14077
rect 11727 14013 11743 14077
rect 11807 14013 11823 14077
rect 11887 14013 11903 14077
rect 11967 14013 11983 14077
rect 12047 14013 12063 14077
rect 12127 14013 12143 14077
rect 12207 14013 12223 14077
rect 12287 14013 12303 14077
rect 12367 14013 12383 14077
rect 12447 14013 12463 14077
rect 12527 14013 12543 14077
rect 12607 14013 12623 14077
rect 12687 14013 12703 14077
rect 12767 14013 12783 14077
rect 12847 14013 12863 14077
rect 12927 14013 12943 14077
rect 13007 14013 13023 14077
rect 13087 14013 13103 14077
rect 13167 14013 13183 14077
rect 13247 14013 13263 14077
rect 13327 14013 13343 14077
rect 13407 14013 13423 14077
rect 13487 14013 13503 14077
rect 13567 14013 13583 14077
rect 13647 14013 13663 14077
rect 13727 14013 13743 14077
rect 13807 14013 13823 14077
rect 13887 14013 13903 14077
rect 13967 14013 13983 14077
rect 14047 14013 14063 14077
rect 14127 14013 14143 14077
rect 14207 14013 14223 14077
rect 14287 14013 14303 14077
rect 14367 14013 14383 14077
rect 14447 14013 14463 14077
rect 14527 14013 14543 14077
rect 14607 14013 14623 14077
rect 14687 14013 14703 14077
rect 14767 14013 14783 14077
rect 14847 14013 14858 14077
rect 10078 14007 14858 14013
rect 99 13704 4879 13706
rect 99 13640 105 13704
rect 169 13640 186 13704
rect 250 13640 267 13704
rect 331 13640 348 13704
rect 412 13640 429 13704
rect 493 13640 510 13704
rect 574 13640 591 13704
rect 655 13640 672 13704
rect 736 13640 753 13704
rect 817 13640 834 13704
rect 898 13640 915 13704
rect 979 13640 996 13704
rect 1060 13640 1077 13704
rect 1141 13640 1158 13704
rect 1222 13640 1239 13704
rect 1303 13640 1320 13704
rect 1384 13640 1401 13704
rect 1465 13640 1482 13704
rect 1546 13640 1563 13704
rect 1627 13640 1644 13704
rect 1708 13640 1725 13704
rect 1789 13640 1806 13704
rect 1870 13640 1887 13704
rect 1951 13640 1968 13704
rect 2032 13640 2049 13704
rect 2113 13640 2130 13704
rect 2194 13640 2211 13704
rect 2275 13640 2292 13704
rect 2356 13640 2373 13704
rect 2437 13640 2454 13704
rect 2518 13640 2535 13704
rect 2599 13640 2616 13704
rect 2680 13640 2697 13704
rect 2761 13640 2778 13704
rect 2842 13640 2859 13704
rect 2923 13640 2940 13704
rect 3004 13640 3021 13704
rect 3085 13640 3102 13704
rect 3166 13640 3183 13704
rect 3247 13640 3264 13704
rect 3328 13640 3345 13704
rect 3409 13640 3426 13704
rect 3490 13640 3507 13704
rect 3571 13640 3588 13704
rect 3652 13640 3669 13704
rect 3733 13640 3750 13704
rect 3814 13640 3831 13704
rect 3895 13640 3912 13704
rect 3976 13640 3993 13704
rect 4057 13640 4074 13704
rect 4138 13640 4155 13704
rect 4219 13640 4236 13704
rect 4300 13640 4317 13704
rect 4381 13640 4399 13704
rect 4463 13640 4481 13704
rect 4545 13640 4563 13704
rect 4627 13640 4645 13704
rect 4709 13640 4727 13704
rect 4791 13640 4809 13704
rect 4873 13640 4879 13704
rect 99 13622 4879 13640
rect 99 13558 105 13622
rect 169 13558 186 13622
rect 250 13558 267 13622
rect 331 13558 348 13622
rect 412 13558 429 13622
rect 493 13558 510 13622
rect 574 13558 591 13622
rect 655 13558 672 13622
rect 736 13558 753 13622
rect 817 13558 834 13622
rect 898 13558 915 13622
rect 979 13558 996 13622
rect 1060 13558 1077 13622
rect 1141 13558 1158 13622
rect 1222 13558 1239 13622
rect 1303 13558 1320 13622
rect 1384 13558 1401 13622
rect 1465 13558 1482 13622
rect 1546 13558 1563 13622
rect 1627 13558 1644 13622
rect 1708 13558 1725 13622
rect 1789 13558 1806 13622
rect 1870 13558 1887 13622
rect 1951 13558 1968 13622
rect 2032 13558 2049 13622
rect 2113 13558 2130 13622
rect 2194 13558 2211 13622
rect 2275 13558 2292 13622
rect 2356 13558 2373 13622
rect 2437 13558 2454 13622
rect 2518 13558 2535 13622
rect 2599 13558 2616 13622
rect 2680 13558 2697 13622
rect 2761 13558 2778 13622
rect 2842 13558 2859 13622
rect 2923 13558 2940 13622
rect 3004 13558 3021 13622
rect 3085 13558 3102 13622
rect 3166 13558 3183 13622
rect 3247 13558 3264 13622
rect 3328 13558 3345 13622
rect 3409 13558 3426 13622
rect 3490 13558 3507 13622
rect 3571 13558 3588 13622
rect 3652 13558 3669 13622
rect 3733 13558 3750 13622
rect 3814 13558 3831 13622
rect 3895 13558 3912 13622
rect 3976 13558 3993 13622
rect 4057 13558 4074 13622
rect 4138 13558 4155 13622
rect 4219 13558 4236 13622
rect 4300 13558 4317 13622
rect 4381 13558 4399 13622
rect 4463 13558 4481 13622
rect 4545 13558 4563 13622
rect 4627 13558 4645 13622
rect 4709 13558 4727 13622
rect 4791 13558 4809 13622
rect 4873 13558 4879 13622
rect 99 13540 4879 13558
rect 99 13476 105 13540
rect 169 13476 186 13540
rect 250 13476 267 13540
rect 331 13476 348 13540
rect 412 13476 429 13540
rect 493 13476 510 13540
rect 574 13476 591 13540
rect 655 13476 672 13540
rect 736 13476 753 13540
rect 817 13476 834 13540
rect 898 13476 915 13540
rect 979 13476 996 13540
rect 1060 13476 1077 13540
rect 1141 13476 1158 13540
rect 1222 13476 1239 13540
rect 1303 13476 1320 13540
rect 1384 13476 1401 13540
rect 1465 13476 1482 13540
rect 1546 13476 1563 13540
rect 1627 13476 1644 13540
rect 1708 13476 1725 13540
rect 1789 13476 1806 13540
rect 1870 13476 1887 13540
rect 1951 13476 1968 13540
rect 2032 13476 2049 13540
rect 2113 13476 2130 13540
rect 2194 13476 2211 13540
rect 2275 13476 2292 13540
rect 2356 13476 2373 13540
rect 2437 13476 2454 13540
rect 2518 13476 2535 13540
rect 2599 13476 2616 13540
rect 2680 13476 2697 13540
rect 2761 13476 2778 13540
rect 2842 13476 2859 13540
rect 2923 13476 2940 13540
rect 3004 13476 3021 13540
rect 3085 13476 3102 13540
rect 3166 13476 3183 13540
rect 3247 13476 3264 13540
rect 3328 13476 3345 13540
rect 3409 13476 3426 13540
rect 3490 13476 3507 13540
rect 3571 13476 3588 13540
rect 3652 13476 3669 13540
rect 3733 13476 3750 13540
rect 3814 13476 3831 13540
rect 3895 13476 3912 13540
rect 3976 13476 3993 13540
rect 4057 13476 4074 13540
rect 4138 13476 4155 13540
rect 4219 13476 4236 13540
rect 4300 13476 4317 13540
rect 4381 13476 4399 13540
rect 4463 13476 4481 13540
rect 4545 13476 4563 13540
rect 4627 13476 4645 13540
rect 4709 13476 4727 13540
rect 4791 13476 4809 13540
rect 4873 13476 4879 13540
rect 99 13458 4879 13476
rect 99 13394 105 13458
rect 169 13394 186 13458
rect 250 13394 267 13458
rect 331 13394 348 13458
rect 412 13394 429 13458
rect 493 13394 510 13458
rect 574 13394 591 13458
rect 655 13394 672 13458
rect 736 13394 753 13458
rect 817 13394 834 13458
rect 898 13394 915 13458
rect 979 13394 996 13458
rect 1060 13394 1077 13458
rect 1141 13394 1158 13458
rect 1222 13394 1239 13458
rect 1303 13394 1320 13458
rect 1384 13394 1401 13458
rect 1465 13394 1482 13458
rect 1546 13394 1563 13458
rect 1627 13394 1644 13458
rect 1708 13394 1725 13458
rect 1789 13394 1806 13458
rect 1870 13394 1887 13458
rect 1951 13394 1968 13458
rect 2032 13394 2049 13458
rect 2113 13394 2130 13458
rect 2194 13394 2211 13458
rect 2275 13394 2292 13458
rect 2356 13394 2373 13458
rect 2437 13394 2454 13458
rect 2518 13394 2535 13458
rect 2599 13394 2616 13458
rect 2680 13394 2697 13458
rect 2761 13394 2778 13458
rect 2842 13394 2859 13458
rect 2923 13394 2940 13458
rect 3004 13394 3021 13458
rect 3085 13394 3102 13458
rect 3166 13394 3183 13458
rect 3247 13394 3264 13458
rect 3328 13394 3345 13458
rect 3409 13394 3426 13458
rect 3490 13394 3507 13458
rect 3571 13394 3588 13458
rect 3652 13394 3669 13458
rect 3733 13394 3750 13458
rect 3814 13394 3831 13458
rect 3895 13394 3912 13458
rect 3976 13394 3993 13458
rect 4057 13394 4074 13458
rect 4138 13394 4155 13458
rect 4219 13394 4236 13458
rect 4300 13394 4317 13458
rect 4381 13394 4399 13458
rect 4463 13394 4481 13458
rect 4545 13394 4563 13458
rect 4627 13394 4645 13458
rect 4709 13394 4727 13458
rect 4791 13394 4809 13458
rect 4873 13394 4879 13458
rect 99 13376 4879 13394
rect 99 13312 105 13376
rect 169 13312 186 13376
rect 250 13312 267 13376
rect 331 13312 348 13376
rect 412 13312 429 13376
rect 493 13312 510 13376
rect 574 13312 591 13376
rect 655 13312 672 13376
rect 736 13312 753 13376
rect 817 13312 834 13376
rect 898 13312 915 13376
rect 979 13312 996 13376
rect 1060 13312 1077 13376
rect 1141 13312 1158 13376
rect 1222 13312 1239 13376
rect 1303 13312 1320 13376
rect 1384 13312 1401 13376
rect 1465 13312 1482 13376
rect 1546 13312 1563 13376
rect 1627 13312 1644 13376
rect 1708 13312 1725 13376
rect 1789 13312 1806 13376
rect 1870 13312 1887 13376
rect 1951 13312 1968 13376
rect 2032 13312 2049 13376
rect 2113 13312 2130 13376
rect 2194 13312 2211 13376
rect 2275 13312 2292 13376
rect 2356 13312 2373 13376
rect 2437 13312 2454 13376
rect 2518 13312 2535 13376
rect 2599 13312 2616 13376
rect 2680 13312 2697 13376
rect 2761 13312 2778 13376
rect 2842 13312 2859 13376
rect 2923 13312 2940 13376
rect 3004 13312 3021 13376
rect 3085 13312 3102 13376
rect 3166 13312 3183 13376
rect 3247 13312 3264 13376
rect 3328 13312 3345 13376
rect 3409 13312 3426 13376
rect 3490 13312 3507 13376
rect 3571 13312 3588 13376
rect 3652 13312 3669 13376
rect 3733 13312 3750 13376
rect 3814 13312 3831 13376
rect 3895 13312 3912 13376
rect 3976 13312 3993 13376
rect 4057 13312 4074 13376
rect 4138 13312 4155 13376
rect 4219 13312 4236 13376
rect 4300 13312 4317 13376
rect 4381 13312 4399 13376
rect 4463 13312 4481 13376
rect 4545 13312 4563 13376
rect 4627 13312 4645 13376
rect 4709 13312 4727 13376
rect 4791 13312 4809 13376
rect 4873 13312 4879 13376
rect 99 13294 4879 13312
rect 99 13230 105 13294
rect 169 13230 186 13294
rect 250 13230 267 13294
rect 331 13230 348 13294
rect 412 13230 429 13294
rect 493 13230 510 13294
rect 574 13230 591 13294
rect 655 13230 672 13294
rect 736 13230 753 13294
rect 817 13230 834 13294
rect 898 13230 915 13294
rect 979 13230 996 13294
rect 1060 13230 1077 13294
rect 1141 13230 1158 13294
rect 1222 13230 1239 13294
rect 1303 13230 1320 13294
rect 1384 13230 1401 13294
rect 1465 13230 1482 13294
rect 1546 13230 1563 13294
rect 1627 13230 1644 13294
rect 1708 13230 1725 13294
rect 1789 13230 1806 13294
rect 1870 13230 1887 13294
rect 1951 13230 1968 13294
rect 2032 13230 2049 13294
rect 2113 13230 2130 13294
rect 2194 13230 2211 13294
rect 2275 13230 2292 13294
rect 2356 13230 2373 13294
rect 2437 13230 2454 13294
rect 2518 13230 2535 13294
rect 2599 13230 2616 13294
rect 2680 13230 2697 13294
rect 2761 13230 2778 13294
rect 2842 13230 2859 13294
rect 2923 13230 2940 13294
rect 3004 13230 3021 13294
rect 3085 13230 3102 13294
rect 3166 13230 3183 13294
rect 3247 13230 3264 13294
rect 3328 13230 3345 13294
rect 3409 13230 3426 13294
rect 3490 13230 3507 13294
rect 3571 13230 3588 13294
rect 3652 13230 3669 13294
rect 3733 13230 3750 13294
rect 3814 13230 3831 13294
rect 3895 13230 3912 13294
rect 3976 13230 3993 13294
rect 4057 13230 4074 13294
rect 4138 13230 4155 13294
rect 4219 13230 4236 13294
rect 4300 13230 4317 13294
rect 4381 13230 4399 13294
rect 4463 13230 4481 13294
rect 4545 13230 4563 13294
rect 4627 13230 4645 13294
rect 4709 13230 4727 13294
rect 4791 13230 4809 13294
rect 4873 13230 4879 13294
rect 99 13212 4879 13230
rect 99 13148 105 13212
rect 169 13148 186 13212
rect 250 13148 267 13212
rect 331 13148 348 13212
rect 412 13148 429 13212
rect 493 13148 510 13212
rect 574 13148 591 13212
rect 655 13148 672 13212
rect 736 13148 753 13212
rect 817 13148 834 13212
rect 898 13148 915 13212
rect 979 13148 996 13212
rect 1060 13148 1077 13212
rect 1141 13148 1158 13212
rect 1222 13148 1239 13212
rect 1303 13148 1320 13212
rect 1384 13148 1401 13212
rect 1465 13148 1482 13212
rect 1546 13148 1563 13212
rect 1627 13148 1644 13212
rect 1708 13148 1725 13212
rect 1789 13148 1806 13212
rect 1870 13148 1887 13212
rect 1951 13148 1968 13212
rect 2032 13148 2049 13212
rect 2113 13148 2130 13212
rect 2194 13148 2211 13212
rect 2275 13148 2292 13212
rect 2356 13148 2373 13212
rect 2437 13148 2454 13212
rect 2518 13148 2535 13212
rect 2599 13148 2616 13212
rect 2680 13148 2697 13212
rect 2761 13148 2778 13212
rect 2842 13148 2859 13212
rect 2923 13148 2940 13212
rect 3004 13148 3021 13212
rect 3085 13148 3102 13212
rect 3166 13148 3183 13212
rect 3247 13148 3264 13212
rect 3328 13148 3345 13212
rect 3409 13148 3426 13212
rect 3490 13148 3507 13212
rect 3571 13148 3588 13212
rect 3652 13148 3669 13212
rect 3733 13148 3750 13212
rect 3814 13148 3831 13212
rect 3895 13148 3912 13212
rect 3976 13148 3993 13212
rect 4057 13148 4074 13212
rect 4138 13148 4155 13212
rect 4219 13148 4236 13212
rect 4300 13148 4317 13212
rect 4381 13148 4399 13212
rect 4463 13148 4481 13212
rect 4545 13148 4563 13212
rect 4627 13148 4645 13212
rect 4709 13148 4727 13212
rect 4791 13148 4809 13212
rect 4873 13148 4879 13212
rect 99 13130 4879 13148
rect 99 13066 105 13130
rect 169 13066 186 13130
rect 250 13066 267 13130
rect 331 13066 348 13130
rect 412 13066 429 13130
rect 493 13066 510 13130
rect 574 13066 591 13130
rect 655 13066 672 13130
rect 736 13066 753 13130
rect 817 13066 834 13130
rect 898 13066 915 13130
rect 979 13066 996 13130
rect 1060 13066 1077 13130
rect 1141 13066 1158 13130
rect 1222 13066 1239 13130
rect 1303 13066 1320 13130
rect 1384 13066 1401 13130
rect 1465 13066 1482 13130
rect 1546 13066 1563 13130
rect 1627 13066 1644 13130
rect 1708 13066 1725 13130
rect 1789 13066 1806 13130
rect 1870 13066 1887 13130
rect 1951 13066 1968 13130
rect 2032 13066 2049 13130
rect 2113 13066 2130 13130
rect 2194 13066 2211 13130
rect 2275 13066 2292 13130
rect 2356 13066 2373 13130
rect 2437 13066 2454 13130
rect 2518 13066 2535 13130
rect 2599 13066 2616 13130
rect 2680 13066 2697 13130
rect 2761 13066 2778 13130
rect 2842 13066 2859 13130
rect 2923 13066 2940 13130
rect 3004 13066 3021 13130
rect 3085 13066 3102 13130
rect 3166 13066 3183 13130
rect 3247 13066 3264 13130
rect 3328 13066 3345 13130
rect 3409 13066 3426 13130
rect 3490 13066 3507 13130
rect 3571 13066 3588 13130
rect 3652 13066 3669 13130
rect 3733 13066 3750 13130
rect 3814 13066 3831 13130
rect 3895 13066 3912 13130
rect 3976 13066 3993 13130
rect 4057 13066 4074 13130
rect 4138 13066 4155 13130
rect 4219 13066 4236 13130
rect 4300 13066 4317 13130
rect 4381 13066 4399 13130
rect 4463 13066 4481 13130
rect 4545 13066 4563 13130
rect 4627 13066 4645 13130
rect 4709 13066 4727 13130
rect 4791 13066 4809 13130
rect 4873 13066 4879 13130
rect 99 13048 4879 13066
rect 99 12984 105 13048
rect 169 12984 186 13048
rect 250 12984 267 13048
rect 331 12984 348 13048
rect 412 12984 429 13048
rect 493 12984 510 13048
rect 574 12984 591 13048
rect 655 12984 672 13048
rect 736 12984 753 13048
rect 817 12984 834 13048
rect 898 12984 915 13048
rect 979 12984 996 13048
rect 1060 12984 1077 13048
rect 1141 12984 1158 13048
rect 1222 12984 1239 13048
rect 1303 12984 1320 13048
rect 1384 12984 1401 13048
rect 1465 12984 1482 13048
rect 1546 12984 1563 13048
rect 1627 12984 1644 13048
rect 1708 12984 1725 13048
rect 1789 12984 1806 13048
rect 1870 12984 1887 13048
rect 1951 12984 1968 13048
rect 2032 12984 2049 13048
rect 2113 12984 2130 13048
rect 2194 12984 2211 13048
rect 2275 12984 2292 13048
rect 2356 12984 2373 13048
rect 2437 12984 2454 13048
rect 2518 12984 2535 13048
rect 2599 12984 2616 13048
rect 2680 12984 2697 13048
rect 2761 12984 2778 13048
rect 2842 12984 2859 13048
rect 2923 12984 2940 13048
rect 3004 12984 3021 13048
rect 3085 12984 3102 13048
rect 3166 12984 3183 13048
rect 3247 12984 3264 13048
rect 3328 12984 3345 13048
rect 3409 12984 3426 13048
rect 3490 12984 3507 13048
rect 3571 12984 3588 13048
rect 3652 12984 3669 13048
rect 3733 12984 3750 13048
rect 3814 12984 3831 13048
rect 3895 12984 3912 13048
rect 3976 12984 3993 13048
rect 4057 12984 4074 13048
rect 4138 12984 4155 13048
rect 4219 12984 4236 13048
rect 4300 12984 4317 13048
rect 4381 12984 4399 13048
rect 4463 12984 4481 13048
rect 4545 12984 4563 13048
rect 4627 12984 4645 13048
rect 4709 12984 4727 13048
rect 4791 12984 4809 13048
rect 4873 12984 4879 13048
rect 99 12966 4879 12984
rect 99 12902 105 12966
rect 169 12902 186 12966
rect 250 12902 267 12966
rect 331 12902 348 12966
rect 412 12902 429 12966
rect 493 12902 510 12966
rect 574 12902 591 12966
rect 655 12902 672 12966
rect 736 12902 753 12966
rect 817 12902 834 12966
rect 898 12902 915 12966
rect 979 12902 996 12966
rect 1060 12902 1077 12966
rect 1141 12902 1158 12966
rect 1222 12902 1239 12966
rect 1303 12902 1320 12966
rect 1384 12902 1401 12966
rect 1465 12902 1482 12966
rect 1546 12902 1563 12966
rect 1627 12902 1644 12966
rect 1708 12902 1725 12966
rect 1789 12902 1806 12966
rect 1870 12902 1887 12966
rect 1951 12902 1968 12966
rect 2032 12902 2049 12966
rect 2113 12902 2130 12966
rect 2194 12902 2211 12966
rect 2275 12902 2292 12966
rect 2356 12902 2373 12966
rect 2437 12902 2454 12966
rect 2518 12902 2535 12966
rect 2599 12902 2616 12966
rect 2680 12902 2697 12966
rect 2761 12902 2778 12966
rect 2842 12902 2859 12966
rect 2923 12902 2940 12966
rect 3004 12902 3021 12966
rect 3085 12902 3102 12966
rect 3166 12902 3183 12966
rect 3247 12902 3264 12966
rect 3328 12902 3345 12966
rect 3409 12902 3426 12966
rect 3490 12902 3507 12966
rect 3571 12902 3588 12966
rect 3652 12902 3669 12966
rect 3733 12902 3750 12966
rect 3814 12902 3831 12966
rect 3895 12902 3912 12966
rect 3976 12902 3993 12966
rect 4057 12902 4074 12966
rect 4138 12902 4155 12966
rect 4219 12902 4236 12966
rect 4300 12902 4317 12966
rect 4381 12902 4399 12966
rect 4463 12902 4481 12966
rect 4545 12902 4563 12966
rect 4627 12902 4645 12966
rect 4709 12902 4727 12966
rect 4791 12902 4809 12966
rect 4873 12902 4879 12966
rect 99 12884 4879 12902
rect 99 12820 105 12884
rect 169 12820 186 12884
rect 250 12820 267 12884
rect 331 12820 348 12884
rect 412 12820 429 12884
rect 493 12820 510 12884
rect 574 12820 591 12884
rect 655 12820 672 12884
rect 736 12820 753 12884
rect 817 12820 834 12884
rect 898 12820 915 12884
rect 979 12820 996 12884
rect 1060 12820 1077 12884
rect 1141 12820 1158 12884
rect 1222 12820 1239 12884
rect 1303 12820 1320 12884
rect 1384 12820 1401 12884
rect 1465 12820 1482 12884
rect 1546 12820 1563 12884
rect 1627 12820 1644 12884
rect 1708 12820 1725 12884
rect 1789 12820 1806 12884
rect 1870 12820 1887 12884
rect 1951 12820 1968 12884
rect 2032 12820 2049 12884
rect 2113 12820 2130 12884
rect 2194 12820 2211 12884
rect 2275 12820 2292 12884
rect 2356 12820 2373 12884
rect 2437 12820 2454 12884
rect 2518 12820 2535 12884
rect 2599 12820 2616 12884
rect 2680 12820 2697 12884
rect 2761 12820 2778 12884
rect 2842 12820 2859 12884
rect 2923 12820 2940 12884
rect 3004 12820 3021 12884
rect 3085 12820 3102 12884
rect 3166 12820 3183 12884
rect 3247 12820 3264 12884
rect 3328 12820 3345 12884
rect 3409 12820 3426 12884
rect 3490 12820 3507 12884
rect 3571 12820 3588 12884
rect 3652 12820 3669 12884
rect 3733 12820 3750 12884
rect 3814 12820 3831 12884
rect 3895 12820 3912 12884
rect 3976 12820 3993 12884
rect 4057 12820 4074 12884
rect 4138 12820 4155 12884
rect 4219 12820 4236 12884
rect 4300 12820 4317 12884
rect 4381 12820 4399 12884
rect 4463 12820 4481 12884
rect 4545 12820 4563 12884
rect 4627 12820 4645 12884
rect 4709 12820 4727 12884
rect 4791 12820 4809 12884
rect 4873 12820 4879 12884
rect 99 12818 4879 12820
rect 10078 13704 14858 13706
rect 10078 13640 10084 13704
rect 10148 13640 10165 13704
rect 10229 13640 10246 13704
rect 10310 13640 10327 13704
rect 10391 13640 10408 13704
rect 10472 13640 10489 13704
rect 10553 13640 10570 13704
rect 10634 13640 10651 13704
rect 10715 13640 10732 13704
rect 10796 13640 10813 13704
rect 10877 13640 10894 13704
rect 10958 13640 10975 13704
rect 11039 13640 11056 13704
rect 11120 13640 11137 13704
rect 11201 13640 11218 13704
rect 11282 13640 11299 13704
rect 11363 13640 11380 13704
rect 11444 13640 11461 13704
rect 11525 13640 11542 13704
rect 11606 13640 11623 13704
rect 11687 13640 11704 13704
rect 11768 13640 11785 13704
rect 11849 13640 11866 13704
rect 11930 13640 11947 13704
rect 12011 13640 12028 13704
rect 12092 13640 12109 13704
rect 12173 13640 12190 13704
rect 12254 13640 12271 13704
rect 12335 13640 12352 13704
rect 12416 13640 12433 13704
rect 12497 13640 12514 13704
rect 12578 13640 12595 13704
rect 12659 13640 12676 13704
rect 12740 13640 12757 13704
rect 12821 13640 12838 13704
rect 12902 13640 12919 13704
rect 12983 13640 13000 13704
rect 13064 13640 13081 13704
rect 13145 13640 13162 13704
rect 13226 13640 13243 13704
rect 13307 13640 13324 13704
rect 13388 13640 13405 13704
rect 13469 13640 13486 13704
rect 13550 13640 13567 13704
rect 13631 13640 13648 13704
rect 13712 13640 13729 13704
rect 13793 13640 13810 13704
rect 13874 13640 13891 13704
rect 13955 13640 13972 13704
rect 14036 13640 14053 13704
rect 14117 13640 14134 13704
rect 14198 13640 14215 13704
rect 14279 13640 14296 13704
rect 14360 13640 14378 13704
rect 14442 13640 14460 13704
rect 14524 13640 14542 13704
rect 14606 13640 14624 13704
rect 14688 13640 14706 13704
rect 14770 13640 14788 13704
rect 14852 13640 14858 13704
rect 10078 13622 14858 13640
rect 10078 13558 10084 13622
rect 10148 13558 10165 13622
rect 10229 13558 10246 13622
rect 10310 13558 10327 13622
rect 10391 13558 10408 13622
rect 10472 13558 10489 13622
rect 10553 13558 10570 13622
rect 10634 13558 10651 13622
rect 10715 13558 10732 13622
rect 10796 13558 10813 13622
rect 10877 13558 10894 13622
rect 10958 13558 10975 13622
rect 11039 13558 11056 13622
rect 11120 13558 11137 13622
rect 11201 13558 11218 13622
rect 11282 13558 11299 13622
rect 11363 13558 11380 13622
rect 11444 13558 11461 13622
rect 11525 13558 11542 13622
rect 11606 13558 11623 13622
rect 11687 13558 11704 13622
rect 11768 13558 11785 13622
rect 11849 13558 11866 13622
rect 11930 13558 11947 13622
rect 12011 13558 12028 13622
rect 12092 13558 12109 13622
rect 12173 13558 12190 13622
rect 12254 13558 12271 13622
rect 12335 13558 12352 13622
rect 12416 13558 12433 13622
rect 12497 13558 12514 13622
rect 12578 13558 12595 13622
rect 12659 13558 12676 13622
rect 12740 13558 12757 13622
rect 12821 13558 12838 13622
rect 12902 13558 12919 13622
rect 12983 13558 13000 13622
rect 13064 13558 13081 13622
rect 13145 13558 13162 13622
rect 13226 13558 13243 13622
rect 13307 13558 13324 13622
rect 13388 13558 13405 13622
rect 13469 13558 13486 13622
rect 13550 13558 13567 13622
rect 13631 13558 13648 13622
rect 13712 13558 13729 13622
rect 13793 13558 13810 13622
rect 13874 13558 13891 13622
rect 13955 13558 13972 13622
rect 14036 13558 14053 13622
rect 14117 13558 14134 13622
rect 14198 13558 14215 13622
rect 14279 13558 14296 13622
rect 14360 13558 14378 13622
rect 14442 13558 14460 13622
rect 14524 13558 14542 13622
rect 14606 13558 14624 13622
rect 14688 13558 14706 13622
rect 14770 13558 14788 13622
rect 14852 13558 14858 13622
rect 10078 13540 14858 13558
rect 10078 13476 10084 13540
rect 10148 13476 10165 13540
rect 10229 13476 10246 13540
rect 10310 13476 10327 13540
rect 10391 13476 10408 13540
rect 10472 13476 10489 13540
rect 10553 13476 10570 13540
rect 10634 13476 10651 13540
rect 10715 13476 10732 13540
rect 10796 13476 10813 13540
rect 10877 13476 10894 13540
rect 10958 13476 10975 13540
rect 11039 13476 11056 13540
rect 11120 13476 11137 13540
rect 11201 13476 11218 13540
rect 11282 13476 11299 13540
rect 11363 13476 11380 13540
rect 11444 13476 11461 13540
rect 11525 13476 11542 13540
rect 11606 13476 11623 13540
rect 11687 13476 11704 13540
rect 11768 13476 11785 13540
rect 11849 13476 11866 13540
rect 11930 13476 11947 13540
rect 12011 13476 12028 13540
rect 12092 13476 12109 13540
rect 12173 13476 12190 13540
rect 12254 13476 12271 13540
rect 12335 13476 12352 13540
rect 12416 13476 12433 13540
rect 12497 13476 12514 13540
rect 12578 13476 12595 13540
rect 12659 13476 12676 13540
rect 12740 13476 12757 13540
rect 12821 13476 12838 13540
rect 12902 13476 12919 13540
rect 12983 13476 13000 13540
rect 13064 13476 13081 13540
rect 13145 13476 13162 13540
rect 13226 13476 13243 13540
rect 13307 13476 13324 13540
rect 13388 13476 13405 13540
rect 13469 13476 13486 13540
rect 13550 13476 13567 13540
rect 13631 13476 13648 13540
rect 13712 13476 13729 13540
rect 13793 13476 13810 13540
rect 13874 13476 13891 13540
rect 13955 13476 13972 13540
rect 14036 13476 14053 13540
rect 14117 13476 14134 13540
rect 14198 13476 14215 13540
rect 14279 13476 14296 13540
rect 14360 13476 14378 13540
rect 14442 13476 14460 13540
rect 14524 13476 14542 13540
rect 14606 13476 14624 13540
rect 14688 13476 14706 13540
rect 14770 13476 14788 13540
rect 14852 13476 14858 13540
rect 10078 13458 14858 13476
rect 10078 13394 10084 13458
rect 10148 13394 10165 13458
rect 10229 13394 10246 13458
rect 10310 13394 10327 13458
rect 10391 13394 10408 13458
rect 10472 13394 10489 13458
rect 10553 13394 10570 13458
rect 10634 13394 10651 13458
rect 10715 13394 10732 13458
rect 10796 13394 10813 13458
rect 10877 13394 10894 13458
rect 10958 13394 10975 13458
rect 11039 13394 11056 13458
rect 11120 13394 11137 13458
rect 11201 13394 11218 13458
rect 11282 13394 11299 13458
rect 11363 13394 11380 13458
rect 11444 13394 11461 13458
rect 11525 13394 11542 13458
rect 11606 13394 11623 13458
rect 11687 13394 11704 13458
rect 11768 13394 11785 13458
rect 11849 13394 11866 13458
rect 11930 13394 11947 13458
rect 12011 13394 12028 13458
rect 12092 13394 12109 13458
rect 12173 13394 12190 13458
rect 12254 13394 12271 13458
rect 12335 13394 12352 13458
rect 12416 13394 12433 13458
rect 12497 13394 12514 13458
rect 12578 13394 12595 13458
rect 12659 13394 12676 13458
rect 12740 13394 12757 13458
rect 12821 13394 12838 13458
rect 12902 13394 12919 13458
rect 12983 13394 13000 13458
rect 13064 13394 13081 13458
rect 13145 13394 13162 13458
rect 13226 13394 13243 13458
rect 13307 13394 13324 13458
rect 13388 13394 13405 13458
rect 13469 13394 13486 13458
rect 13550 13394 13567 13458
rect 13631 13394 13648 13458
rect 13712 13394 13729 13458
rect 13793 13394 13810 13458
rect 13874 13394 13891 13458
rect 13955 13394 13972 13458
rect 14036 13394 14053 13458
rect 14117 13394 14134 13458
rect 14198 13394 14215 13458
rect 14279 13394 14296 13458
rect 14360 13394 14378 13458
rect 14442 13394 14460 13458
rect 14524 13394 14542 13458
rect 14606 13394 14624 13458
rect 14688 13394 14706 13458
rect 14770 13394 14788 13458
rect 14852 13394 14858 13458
rect 10078 13376 14858 13394
rect 10078 13312 10084 13376
rect 10148 13312 10165 13376
rect 10229 13312 10246 13376
rect 10310 13312 10327 13376
rect 10391 13312 10408 13376
rect 10472 13312 10489 13376
rect 10553 13312 10570 13376
rect 10634 13312 10651 13376
rect 10715 13312 10732 13376
rect 10796 13312 10813 13376
rect 10877 13312 10894 13376
rect 10958 13312 10975 13376
rect 11039 13312 11056 13376
rect 11120 13312 11137 13376
rect 11201 13312 11218 13376
rect 11282 13312 11299 13376
rect 11363 13312 11380 13376
rect 11444 13312 11461 13376
rect 11525 13312 11542 13376
rect 11606 13312 11623 13376
rect 11687 13312 11704 13376
rect 11768 13312 11785 13376
rect 11849 13312 11866 13376
rect 11930 13312 11947 13376
rect 12011 13312 12028 13376
rect 12092 13312 12109 13376
rect 12173 13312 12190 13376
rect 12254 13312 12271 13376
rect 12335 13312 12352 13376
rect 12416 13312 12433 13376
rect 12497 13312 12514 13376
rect 12578 13312 12595 13376
rect 12659 13312 12676 13376
rect 12740 13312 12757 13376
rect 12821 13312 12838 13376
rect 12902 13312 12919 13376
rect 12983 13312 13000 13376
rect 13064 13312 13081 13376
rect 13145 13312 13162 13376
rect 13226 13312 13243 13376
rect 13307 13312 13324 13376
rect 13388 13312 13405 13376
rect 13469 13312 13486 13376
rect 13550 13312 13567 13376
rect 13631 13312 13648 13376
rect 13712 13312 13729 13376
rect 13793 13312 13810 13376
rect 13874 13312 13891 13376
rect 13955 13312 13972 13376
rect 14036 13312 14053 13376
rect 14117 13312 14134 13376
rect 14198 13312 14215 13376
rect 14279 13312 14296 13376
rect 14360 13312 14378 13376
rect 14442 13312 14460 13376
rect 14524 13312 14542 13376
rect 14606 13312 14624 13376
rect 14688 13312 14706 13376
rect 14770 13312 14788 13376
rect 14852 13312 14858 13376
rect 10078 13294 14858 13312
rect 10078 13230 10084 13294
rect 10148 13230 10165 13294
rect 10229 13230 10246 13294
rect 10310 13230 10327 13294
rect 10391 13230 10408 13294
rect 10472 13230 10489 13294
rect 10553 13230 10570 13294
rect 10634 13230 10651 13294
rect 10715 13230 10732 13294
rect 10796 13230 10813 13294
rect 10877 13230 10894 13294
rect 10958 13230 10975 13294
rect 11039 13230 11056 13294
rect 11120 13230 11137 13294
rect 11201 13230 11218 13294
rect 11282 13230 11299 13294
rect 11363 13230 11380 13294
rect 11444 13230 11461 13294
rect 11525 13230 11542 13294
rect 11606 13230 11623 13294
rect 11687 13230 11704 13294
rect 11768 13230 11785 13294
rect 11849 13230 11866 13294
rect 11930 13230 11947 13294
rect 12011 13230 12028 13294
rect 12092 13230 12109 13294
rect 12173 13230 12190 13294
rect 12254 13230 12271 13294
rect 12335 13230 12352 13294
rect 12416 13230 12433 13294
rect 12497 13230 12514 13294
rect 12578 13230 12595 13294
rect 12659 13230 12676 13294
rect 12740 13230 12757 13294
rect 12821 13230 12838 13294
rect 12902 13230 12919 13294
rect 12983 13230 13000 13294
rect 13064 13230 13081 13294
rect 13145 13230 13162 13294
rect 13226 13230 13243 13294
rect 13307 13230 13324 13294
rect 13388 13230 13405 13294
rect 13469 13230 13486 13294
rect 13550 13230 13567 13294
rect 13631 13230 13648 13294
rect 13712 13230 13729 13294
rect 13793 13230 13810 13294
rect 13874 13230 13891 13294
rect 13955 13230 13972 13294
rect 14036 13230 14053 13294
rect 14117 13230 14134 13294
rect 14198 13230 14215 13294
rect 14279 13230 14296 13294
rect 14360 13230 14378 13294
rect 14442 13230 14460 13294
rect 14524 13230 14542 13294
rect 14606 13230 14624 13294
rect 14688 13230 14706 13294
rect 14770 13230 14788 13294
rect 14852 13230 14858 13294
rect 10078 13212 14858 13230
rect 10078 13148 10084 13212
rect 10148 13148 10165 13212
rect 10229 13148 10246 13212
rect 10310 13148 10327 13212
rect 10391 13148 10408 13212
rect 10472 13148 10489 13212
rect 10553 13148 10570 13212
rect 10634 13148 10651 13212
rect 10715 13148 10732 13212
rect 10796 13148 10813 13212
rect 10877 13148 10894 13212
rect 10958 13148 10975 13212
rect 11039 13148 11056 13212
rect 11120 13148 11137 13212
rect 11201 13148 11218 13212
rect 11282 13148 11299 13212
rect 11363 13148 11380 13212
rect 11444 13148 11461 13212
rect 11525 13148 11542 13212
rect 11606 13148 11623 13212
rect 11687 13148 11704 13212
rect 11768 13148 11785 13212
rect 11849 13148 11866 13212
rect 11930 13148 11947 13212
rect 12011 13148 12028 13212
rect 12092 13148 12109 13212
rect 12173 13148 12190 13212
rect 12254 13148 12271 13212
rect 12335 13148 12352 13212
rect 12416 13148 12433 13212
rect 12497 13148 12514 13212
rect 12578 13148 12595 13212
rect 12659 13148 12676 13212
rect 12740 13148 12757 13212
rect 12821 13148 12838 13212
rect 12902 13148 12919 13212
rect 12983 13148 13000 13212
rect 13064 13148 13081 13212
rect 13145 13148 13162 13212
rect 13226 13148 13243 13212
rect 13307 13148 13324 13212
rect 13388 13148 13405 13212
rect 13469 13148 13486 13212
rect 13550 13148 13567 13212
rect 13631 13148 13648 13212
rect 13712 13148 13729 13212
rect 13793 13148 13810 13212
rect 13874 13148 13891 13212
rect 13955 13148 13972 13212
rect 14036 13148 14053 13212
rect 14117 13148 14134 13212
rect 14198 13148 14215 13212
rect 14279 13148 14296 13212
rect 14360 13148 14378 13212
rect 14442 13148 14460 13212
rect 14524 13148 14542 13212
rect 14606 13148 14624 13212
rect 14688 13148 14706 13212
rect 14770 13148 14788 13212
rect 14852 13148 14858 13212
rect 10078 13130 14858 13148
rect 10078 13066 10084 13130
rect 10148 13066 10165 13130
rect 10229 13066 10246 13130
rect 10310 13066 10327 13130
rect 10391 13066 10408 13130
rect 10472 13066 10489 13130
rect 10553 13066 10570 13130
rect 10634 13066 10651 13130
rect 10715 13066 10732 13130
rect 10796 13066 10813 13130
rect 10877 13066 10894 13130
rect 10958 13066 10975 13130
rect 11039 13066 11056 13130
rect 11120 13066 11137 13130
rect 11201 13066 11218 13130
rect 11282 13066 11299 13130
rect 11363 13066 11380 13130
rect 11444 13066 11461 13130
rect 11525 13066 11542 13130
rect 11606 13066 11623 13130
rect 11687 13066 11704 13130
rect 11768 13066 11785 13130
rect 11849 13066 11866 13130
rect 11930 13066 11947 13130
rect 12011 13066 12028 13130
rect 12092 13066 12109 13130
rect 12173 13066 12190 13130
rect 12254 13066 12271 13130
rect 12335 13066 12352 13130
rect 12416 13066 12433 13130
rect 12497 13066 12514 13130
rect 12578 13066 12595 13130
rect 12659 13066 12676 13130
rect 12740 13066 12757 13130
rect 12821 13066 12838 13130
rect 12902 13066 12919 13130
rect 12983 13066 13000 13130
rect 13064 13066 13081 13130
rect 13145 13066 13162 13130
rect 13226 13066 13243 13130
rect 13307 13066 13324 13130
rect 13388 13066 13405 13130
rect 13469 13066 13486 13130
rect 13550 13066 13567 13130
rect 13631 13066 13648 13130
rect 13712 13066 13729 13130
rect 13793 13066 13810 13130
rect 13874 13066 13891 13130
rect 13955 13066 13972 13130
rect 14036 13066 14053 13130
rect 14117 13066 14134 13130
rect 14198 13066 14215 13130
rect 14279 13066 14296 13130
rect 14360 13066 14378 13130
rect 14442 13066 14460 13130
rect 14524 13066 14542 13130
rect 14606 13066 14624 13130
rect 14688 13066 14706 13130
rect 14770 13066 14788 13130
rect 14852 13066 14858 13130
rect 10078 13048 14858 13066
rect 10078 12984 10084 13048
rect 10148 12984 10165 13048
rect 10229 12984 10246 13048
rect 10310 12984 10327 13048
rect 10391 12984 10408 13048
rect 10472 12984 10489 13048
rect 10553 12984 10570 13048
rect 10634 12984 10651 13048
rect 10715 12984 10732 13048
rect 10796 12984 10813 13048
rect 10877 12984 10894 13048
rect 10958 12984 10975 13048
rect 11039 12984 11056 13048
rect 11120 12984 11137 13048
rect 11201 12984 11218 13048
rect 11282 12984 11299 13048
rect 11363 12984 11380 13048
rect 11444 12984 11461 13048
rect 11525 12984 11542 13048
rect 11606 12984 11623 13048
rect 11687 12984 11704 13048
rect 11768 12984 11785 13048
rect 11849 12984 11866 13048
rect 11930 12984 11947 13048
rect 12011 12984 12028 13048
rect 12092 12984 12109 13048
rect 12173 12984 12190 13048
rect 12254 12984 12271 13048
rect 12335 12984 12352 13048
rect 12416 12984 12433 13048
rect 12497 12984 12514 13048
rect 12578 12984 12595 13048
rect 12659 12984 12676 13048
rect 12740 12984 12757 13048
rect 12821 12984 12838 13048
rect 12902 12984 12919 13048
rect 12983 12984 13000 13048
rect 13064 12984 13081 13048
rect 13145 12984 13162 13048
rect 13226 12984 13243 13048
rect 13307 12984 13324 13048
rect 13388 12984 13405 13048
rect 13469 12984 13486 13048
rect 13550 12984 13567 13048
rect 13631 12984 13648 13048
rect 13712 12984 13729 13048
rect 13793 12984 13810 13048
rect 13874 12984 13891 13048
rect 13955 12984 13972 13048
rect 14036 12984 14053 13048
rect 14117 12984 14134 13048
rect 14198 12984 14215 13048
rect 14279 12984 14296 13048
rect 14360 12984 14378 13048
rect 14442 12984 14460 13048
rect 14524 12984 14542 13048
rect 14606 12984 14624 13048
rect 14688 12984 14706 13048
rect 14770 12984 14788 13048
rect 14852 12984 14858 13048
rect 10078 12966 14858 12984
rect 10078 12902 10084 12966
rect 10148 12902 10165 12966
rect 10229 12902 10246 12966
rect 10310 12902 10327 12966
rect 10391 12902 10408 12966
rect 10472 12902 10489 12966
rect 10553 12902 10570 12966
rect 10634 12902 10651 12966
rect 10715 12902 10732 12966
rect 10796 12902 10813 12966
rect 10877 12902 10894 12966
rect 10958 12902 10975 12966
rect 11039 12902 11056 12966
rect 11120 12902 11137 12966
rect 11201 12902 11218 12966
rect 11282 12902 11299 12966
rect 11363 12902 11380 12966
rect 11444 12902 11461 12966
rect 11525 12902 11542 12966
rect 11606 12902 11623 12966
rect 11687 12902 11704 12966
rect 11768 12902 11785 12966
rect 11849 12902 11866 12966
rect 11930 12902 11947 12966
rect 12011 12902 12028 12966
rect 12092 12902 12109 12966
rect 12173 12902 12190 12966
rect 12254 12902 12271 12966
rect 12335 12902 12352 12966
rect 12416 12902 12433 12966
rect 12497 12902 12514 12966
rect 12578 12902 12595 12966
rect 12659 12902 12676 12966
rect 12740 12902 12757 12966
rect 12821 12902 12838 12966
rect 12902 12902 12919 12966
rect 12983 12902 13000 12966
rect 13064 12902 13081 12966
rect 13145 12902 13162 12966
rect 13226 12902 13243 12966
rect 13307 12902 13324 12966
rect 13388 12902 13405 12966
rect 13469 12902 13486 12966
rect 13550 12902 13567 12966
rect 13631 12902 13648 12966
rect 13712 12902 13729 12966
rect 13793 12902 13810 12966
rect 13874 12902 13891 12966
rect 13955 12902 13972 12966
rect 14036 12902 14053 12966
rect 14117 12902 14134 12966
rect 14198 12902 14215 12966
rect 14279 12902 14296 12966
rect 14360 12902 14378 12966
rect 14442 12902 14460 12966
rect 14524 12902 14542 12966
rect 14606 12902 14624 12966
rect 14688 12902 14706 12966
rect 14770 12902 14788 12966
rect 14852 12902 14858 12966
rect 10078 12884 14858 12902
rect 10078 12820 10084 12884
rect 10148 12820 10165 12884
rect 10229 12820 10246 12884
rect 10310 12820 10327 12884
rect 10391 12820 10408 12884
rect 10472 12820 10489 12884
rect 10553 12820 10570 12884
rect 10634 12820 10651 12884
rect 10715 12820 10732 12884
rect 10796 12820 10813 12884
rect 10877 12820 10894 12884
rect 10958 12820 10975 12884
rect 11039 12820 11056 12884
rect 11120 12820 11137 12884
rect 11201 12820 11218 12884
rect 11282 12820 11299 12884
rect 11363 12820 11380 12884
rect 11444 12820 11461 12884
rect 11525 12820 11542 12884
rect 11606 12820 11623 12884
rect 11687 12820 11704 12884
rect 11768 12820 11785 12884
rect 11849 12820 11866 12884
rect 11930 12820 11947 12884
rect 12011 12820 12028 12884
rect 12092 12820 12109 12884
rect 12173 12820 12190 12884
rect 12254 12820 12271 12884
rect 12335 12820 12352 12884
rect 12416 12820 12433 12884
rect 12497 12820 12514 12884
rect 12578 12820 12595 12884
rect 12659 12820 12676 12884
rect 12740 12820 12757 12884
rect 12821 12820 12838 12884
rect 12902 12820 12919 12884
rect 12983 12820 13000 12884
rect 13064 12820 13081 12884
rect 13145 12820 13162 12884
rect 13226 12820 13243 12884
rect 13307 12820 13324 12884
rect 13388 12820 13405 12884
rect 13469 12820 13486 12884
rect 13550 12820 13567 12884
rect 13631 12820 13648 12884
rect 13712 12820 13729 12884
rect 13793 12820 13810 12884
rect 13874 12820 13891 12884
rect 13955 12820 13972 12884
rect 14036 12820 14053 12884
rect 14117 12820 14134 12884
rect 14198 12820 14215 12884
rect 14279 12820 14296 12884
rect 14360 12820 14378 12884
rect 14442 12820 14460 12884
rect 14524 12820 14542 12884
rect 14606 12820 14624 12884
rect 14688 12820 14706 12884
rect 14770 12820 14788 12884
rect 14852 12820 14858 12884
rect 10078 12818 14858 12820
rect 99 4884 4879 4886
rect 99 4820 105 4884
rect 169 4820 186 4884
rect 250 4820 267 4884
rect 331 4820 348 4884
rect 412 4820 429 4884
rect 493 4820 510 4884
rect 574 4820 591 4884
rect 655 4820 672 4884
rect 736 4820 753 4884
rect 817 4820 834 4884
rect 898 4820 915 4884
rect 979 4820 996 4884
rect 1060 4820 1077 4884
rect 1141 4820 1158 4884
rect 1222 4820 1239 4884
rect 1303 4820 1320 4884
rect 1384 4820 1401 4884
rect 1465 4820 1482 4884
rect 1546 4820 1563 4884
rect 1627 4820 1644 4884
rect 1708 4820 1725 4884
rect 1789 4820 1806 4884
rect 1870 4820 1887 4884
rect 1951 4820 1968 4884
rect 2032 4820 2049 4884
rect 2113 4820 2130 4884
rect 2194 4820 2211 4884
rect 2275 4820 2292 4884
rect 2356 4820 2373 4884
rect 2437 4820 2454 4884
rect 2518 4820 2535 4884
rect 2599 4820 2616 4884
rect 2680 4820 2697 4884
rect 2761 4820 2778 4884
rect 2842 4820 2859 4884
rect 2923 4820 2940 4884
rect 3004 4820 3021 4884
rect 3085 4820 3102 4884
rect 3166 4820 3183 4884
rect 3247 4820 3264 4884
rect 3328 4820 3345 4884
rect 3409 4820 3426 4884
rect 3490 4820 3507 4884
rect 3571 4820 3588 4884
rect 3652 4820 3669 4884
rect 3733 4820 3750 4884
rect 3814 4820 3831 4884
rect 3895 4820 3912 4884
rect 3976 4820 3993 4884
rect 4057 4820 4074 4884
rect 4138 4820 4155 4884
rect 4219 4820 4236 4884
rect 4300 4820 4317 4884
rect 4381 4820 4399 4884
rect 4463 4820 4481 4884
rect 4545 4820 4563 4884
rect 4627 4820 4645 4884
rect 4709 4820 4727 4884
rect 4791 4820 4809 4884
rect 4873 4820 4879 4884
rect 99 4798 4879 4820
rect 99 4734 105 4798
rect 169 4734 186 4798
rect 250 4734 267 4798
rect 331 4734 348 4798
rect 412 4734 429 4798
rect 493 4734 510 4798
rect 574 4734 591 4798
rect 655 4734 672 4798
rect 736 4734 753 4798
rect 817 4734 834 4798
rect 898 4734 915 4798
rect 979 4734 996 4798
rect 1060 4734 1077 4798
rect 1141 4734 1158 4798
rect 1222 4734 1239 4798
rect 1303 4734 1320 4798
rect 1384 4734 1401 4798
rect 1465 4734 1482 4798
rect 1546 4734 1563 4798
rect 1627 4734 1644 4798
rect 1708 4734 1725 4798
rect 1789 4734 1806 4798
rect 1870 4734 1887 4798
rect 1951 4734 1968 4798
rect 2032 4734 2049 4798
rect 2113 4734 2130 4798
rect 2194 4734 2211 4798
rect 2275 4734 2292 4798
rect 2356 4734 2373 4798
rect 2437 4734 2454 4798
rect 2518 4734 2535 4798
rect 2599 4734 2616 4798
rect 2680 4734 2697 4798
rect 2761 4734 2778 4798
rect 2842 4734 2859 4798
rect 2923 4734 2940 4798
rect 3004 4734 3021 4798
rect 3085 4734 3102 4798
rect 3166 4734 3183 4798
rect 3247 4734 3264 4798
rect 3328 4734 3345 4798
rect 3409 4734 3426 4798
rect 3490 4734 3507 4798
rect 3571 4734 3588 4798
rect 3652 4734 3669 4798
rect 3733 4734 3750 4798
rect 3814 4734 3831 4798
rect 3895 4734 3912 4798
rect 3976 4734 3993 4798
rect 4057 4734 4074 4798
rect 4138 4734 4155 4798
rect 4219 4734 4236 4798
rect 4300 4734 4317 4798
rect 4381 4734 4399 4798
rect 4463 4734 4481 4798
rect 4545 4734 4563 4798
rect 4627 4734 4645 4798
rect 4709 4734 4727 4798
rect 4791 4734 4809 4798
rect 4873 4734 4879 4798
rect 99 4712 4879 4734
rect 99 4648 105 4712
rect 169 4648 186 4712
rect 250 4648 267 4712
rect 331 4648 348 4712
rect 412 4648 429 4712
rect 493 4648 510 4712
rect 574 4648 591 4712
rect 655 4648 672 4712
rect 736 4648 753 4712
rect 817 4648 834 4712
rect 898 4648 915 4712
rect 979 4648 996 4712
rect 1060 4648 1077 4712
rect 1141 4648 1158 4712
rect 1222 4648 1239 4712
rect 1303 4648 1320 4712
rect 1384 4648 1401 4712
rect 1465 4648 1482 4712
rect 1546 4648 1563 4712
rect 1627 4648 1644 4712
rect 1708 4648 1725 4712
rect 1789 4648 1806 4712
rect 1870 4648 1887 4712
rect 1951 4648 1968 4712
rect 2032 4648 2049 4712
rect 2113 4648 2130 4712
rect 2194 4648 2211 4712
rect 2275 4648 2292 4712
rect 2356 4648 2373 4712
rect 2437 4648 2454 4712
rect 2518 4648 2535 4712
rect 2599 4648 2616 4712
rect 2680 4648 2697 4712
rect 2761 4648 2778 4712
rect 2842 4648 2859 4712
rect 2923 4648 2940 4712
rect 3004 4648 3021 4712
rect 3085 4648 3102 4712
rect 3166 4648 3183 4712
rect 3247 4648 3264 4712
rect 3328 4648 3345 4712
rect 3409 4648 3426 4712
rect 3490 4648 3507 4712
rect 3571 4648 3588 4712
rect 3652 4648 3669 4712
rect 3733 4648 3750 4712
rect 3814 4648 3831 4712
rect 3895 4648 3912 4712
rect 3976 4648 3993 4712
rect 4057 4648 4074 4712
rect 4138 4648 4155 4712
rect 4219 4648 4236 4712
rect 4300 4648 4317 4712
rect 4381 4648 4399 4712
rect 4463 4648 4481 4712
rect 4545 4648 4563 4712
rect 4627 4648 4645 4712
rect 4709 4648 4727 4712
rect 4791 4648 4809 4712
rect 4873 4648 4879 4712
rect 99 4626 4879 4648
rect 99 4562 105 4626
rect 169 4562 186 4626
rect 250 4562 267 4626
rect 331 4562 348 4626
rect 412 4562 429 4626
rect 493 4562 510 4626
rect 574 4562 591 4626
rect 655 4562 672 4626
rect 736 4562 753 4626
rect 817 4562 834 4626
rect 898 4562 915 4626
rect 979 4562 996 4626
rect 1060 4562 1077 4626
rect 1141 4562 1158 4626
rect 1222 4562 1239 4626
rect 1303 4562 1320 4626
rect 1384 4562 1401 4626
rect 1465 4562 1482 4626
rect 1546 4562 1563 4626
rect 1627 4562 1644 4626
rect 1708 4562 1725 4626
rect 1789 4562 1806 4626
rect 1870 4562 1887 4626
rect 1951 4562 1968 4626
rect 2032 4562 2049 4626
rect 2113 4562 2130 4626
rect 2194 4562 2211 4626
rect 2275 4562 2292 4626
rect 2356 4562 2373 4626
rect 2437 4562 2454 4626
rect 2518 4562 2535 4626
rect 2599 4562 2616 4626
rect 2680 4562 2697 4626
rect 2761 4562 2778 4626
rect 2842 4562 2859 4626
rect 2923 4562 2940 4626
rect 3004 4562 3021 4626
rect 3085 4562 3102 4626
rect 3166 4562 3183 4626
rect 3247 4562 3264 4626
rect 3328 4562 3345 4626
rect 3409 4562 3426 4626
rect 3490 4562 3507 4626
rect 3571 4562 3588 4626
rect 3652 4562 3669 4626
rect 3733 4562 3750 4626
rect 3814 4562 3831 4626
rect 3895 4562 3912 4626
rect 3976 4562 3993 4626
rect 4057 4562 4074 4626
rect 4138 4562 4155 4626
rect 4219 4562 4236 4626
rect 4300 4562 4317 4626
rect 4381 4562 4399 4626
rect 4463 4562 4481 4626
rect 4545 4562 4563 4626
rect 4627 4562 4645 4626
rect 4709 4562 4727 4626
rect 4791 4562 4809 4626
rect 4873 4562 4879 4626
rect 99 4540 4879 4562
rect 99 4476 105 4540
rect 169 4476 186 4540
rect 250 4476 267 4540
rect 331 4476 348 4540
rect 412 4476 429 4540
rect 493 4476 510 4540
rect 574 4476 591 4540
rect 655 4476 672 4540
rect 736 4476 753 4540
rect 817 4476 834 4540
rect 898 4476 915 4540
rect 979 4476 996 4540
rect 1060 4476 1077 4540
rect 1141 4476 1158 4540
rect 1222 4476 1239 4540
rect 1303 4476 1320 4540
rect 1384 4476 1401 4540
rect 1465 4476 1482 4540
rect 1546 4476 1563 4540
rect 1627 4476 1644 4540
rect 1708 4476 1725 4540
rect 1789 4476 1806 4540
rect 1870 4476 1887 4540
rect 1951 4476 1968 4540
rect 2032 4476 2049 4540
rect 2113 4476 2130 4540
rect 2194 4476 2211 4540
rect 2275 4476 2292 4540
rect 2356 4476 2373 4540
rect 2437 4476 2454 4540
rect 2518 4476 2535 4540
rect 2599 4476 2616 4540
rect 2680 4476 2697 4540
rect 2761 4476 2778 4540
rect 2842 4476 2859 4540
rect 2923 4476 2940 4540
rect 3004 4476 3021 4540
rect 3085 4476 3102 4540
rect 3166 4476 3183 4540
rect 3247 4476 3264 4540
rect 3328 4476 3345 4540
rect 3409 4476 3426 4540
rect 3490 4476 3507 4540
rect 3571 4476 3588 4540
rect 3652 4476 3669 4540
rect 3733 4476 3750 4540
rect 3814 4476 3831 4540
rect 3895 4476 3912 4540
rect 3976 4476 3993 4540
rect 4057 4476 4074 4540
rect 4138 4476 4155 4540
rect 4219 4476 4236 4540
rect 4300 4476 4317 4540
rect 4381 4476 4399 4540
rect 4463 4476 4481 4540
rect 4545 4476 4563 4540
rect 4627 4476 4645 4540
rect 4709 4476 4727 4540
rect 4791 4476 4809 4540
rect 4873 4476 4879 4540
rect 99 4454 4879 4476
rect 99 4390 105 4454
rect 169 4390 186 4454
rect 250 4390 267 4454
rect 331 4390 348 4454
rect 412 4390 429 4454
rect 493 4390 510 4454
rect 574 4390 591 4454
rect 655 4390 672 4454
rect 736 4390 753 4454
rect 817 4390 834 4454
rect 898 4390 915 4454
rect 979 4390 996 4454
rect 1060 4390 1077 4454
rect 1141 4390 1158 4454
rect 1222 4390 1239 4454
rect 1303 4390 1320 4454
rect 1384 4390 1401 4454
rect 1465 4390 1482 4454
rect 1546 4390 1563 4454
rect 1627 4390 1644 4454
rect 1708 4390 1725 4454
rect 1789 4390 1806 4454
rect 1870 4390 1887 4454
rect 1951 4390 1968 4454
rect 2032 4390 2049 4454
rect 2113 4390 2130 4454
rect 2194 4390 2211 4454
rect 2275 4390 2292 4454
rect 2356 4390 2373 4454
rect 2437 4390 2454 4454
rect 2518 4390 2535 4454
rect 2599 4390 2616 4454
rect 2680 4390 2697 4454
rect 2761 4390 2778 4454
rect 2842 4390 2859 4454
rect 2923 4390 2940 4454
rect 3004 4390 3021 4454
rect 3085 4390 3102 4454
rect 3166 4390 3183 4454
rect 3247 4390 3264 4454
rect 3328 4390 3345 4454
rect 3409 4390 3426 4454
rect 3490 4390 3507 4454
rect 3571 4390 3588 4454
rect 3652 4390 3669 4454
rect 3733 4390 3750 4454
rect 3814 4390 3831 4454
rect 3895 4390 3912 4454
rect 3976 4390 3993 4454
rect 4057 4390 4074 4454
rect 4138 4390 4155 4454
rect 4219 4390 4236 4454
rect 4300 4390 4317 4454
rect 4381 4390 4399 4454
rect 4463 4390 4481 4454
rect 4545 4390 4563 4454
rect 4627 4390 4645 4454
rect 4709 4390 4727 4454
rect 4791 4390 4809 4454
rect 4873 4390 4879 4454
rect 99 4368 4879 4390
rect 99 4304 105 4368
rect 169 4304 186 4368
rect 250 4304 267 4368
rect 331 4304 348 4368
rect 412 4304 429 4368
rect 493 4304 510 4368
rect 574 4304 591 4368
rect 655 4304 672 4368
rect 736 4304 753 4368
rect 817 4304 834 4368
rect 898 4304 915 4368
rect 979 4304 996 4368
rect 1060 4304 1077 4368
rect 1141 4304 1158 4368
rect 1222 4304 1239 4368
rect 1303 4304 1320 4368
rect 1384 4304 1401 4368
rect 1465 4304 1482 4368
rect 1546 4304 1563 4368
rect 1627 4304 1644 4368
rect 1708 4304 1725 4368
rect 1789 4304 1806 4368
rect 1870 4304 1887 4368
rect 1951 4304 1968 4368
rect 2032 4304 2049 4368
rect 2113 4304 2130 4368
rect 2194 4304 2211 4368
rect 2275 4304 2292 4368
rect 2356 4304 2373 4368
rect 2437 4304 2454 4368
rect 2518 4304 2535 4368
rect 2599 4304 2616 4368
rect 2680 4304 2697 4368
rect 2761 4304 2778 4368
rect 2842 4304 2859 4368
rect 2923 4304 2940 4368
rect 3004 4304 3021 4368
rect 3085 4304 3102 4368
rect 3166 4304 3183 4368
rect 3247 4304 3264 4368
rect 3328 4304 3345 4368
rect 3409 4304 3426 4368
rect 3490 4304 3507 4368
rect 3571 4304 3588 4368
rect 3652 4304 3669 4368
rect 3733 4304 3750 4368
rect 3814 4304 3831 4368
rect 3895 4304 3912 4368
rect 3976 4304 3993 4368
rect 4057 4304 4074 4368
rect 4138 4304 4155 4368
rect 4219 4304 4236 4368
rect 4300 4304 4317 4368
rect 4381 4304 4399 4368
rect 4463 4304 4481 4368
rect 4545 4304 4563 4368
rect 4627 4304 4645 4368
rect 4709 4304 4727 4368
rect 4791 4304 4809 4368
rect 4873 4304 4879 4368
rect 99 4282 4879 4304
rect 99 4218 105 4282
rect 169 4218 186 4282
rect 250 4218 267 4282
rect 331 4218 348 4282
rect 412 4218 429 4282
rect 493 4218 510 4282
rect 574 4218 591 4282
rect 655 4218 672 4282
rect 736 4218 753 4282
rect 817 4218 834 4282
rect 898 4218 915 4282
rect 979 4218 996 4282
rect 1060 4218 1077 4282
rect 1141 4218 1158 4282
rect 1222 4218 1239 4282
rect 1303 4218 1320 4282
rect 1384 4218 1401 4282
rect 1465 4218 1482 4282
rect 1546 4218 1563 4282
rect 1627 4218 1644 4282
rect 1708 4218 1725 4282
rect 1789 4218 1806 4282
rect 1870 4218 1887 4282
rect 1951 4218 1968 4282
rect 2032 4218 2049 4282
rect 2113 4218 2130 4282
rect 2194 4218 2211 4282
rect 2275 4218 2292 4282
rect 2356 4218 2373 4282
rect 2437 4218 2454 4282
rect 2518 4218 2535 4282
rect 2599 4218 2616 4282
rect 2680 4218 2697 4282
rect 2761 4218 2778 4282
rect 2842 4218 2859 4282
rect 2923 4218 2940 4282
rect 3004 4218 3021 4282
rect 3085 4218 3102 4282
rect 3166 4218 3183 4282
rect 3247 4218 3264 4282
rect 3328 4218 3345 4282
rect 3409 4218 3426 4282
rect 3490 4218 3507 4282
rect 3571 4218 3588 4282
rect 3652 4218 3669 4282
rect 3733 4218 3750 4282
rect 3814 4218 3831 4282
rect 3895 4218 3912 4282
rect 3976 4218 3993 4282
rect 4057 4218 4074 4282
rect 4138 4218 4155 4282
rect 4219 4218 4236 4282
rect 4300 4218 4317 4282
rect 4381 4218 4399 4282
rect 4463 4218 4481 4282
rect 4545 4218 4563 4282
rect 4627 4218 4645 4282
rect 4709 4218 4727 4282
rect 4791 4218 4809 4282
rect 4873 4218 4879 4282
rect 99 4196 4879 4218
rect 99 4132 105 4196
rect 169 4132 186 4196
rect 250 4132 267 4196
rect 331 4132 348 4196
rect 412 4132 429 4196
rect 493 4132 510 4196
rect 574 4132 591 4196
rect 655 4132 672 4196
rect 736 4132 753 4196
rect 817 4132 834 4196
rect 898 4132 915 4196
rect 979 4132 996 4196
rect 1060 4132 1077 4196
rect 1141 4132 1158 4196
rect 1222 4132 1239 4196
rect 1303 4132 1320 4196
rect 1384 4132 1401 4196
rect 1465 4132 1482 4196
rect 1546 4132 1563 4196
rect 1627 4132 1644 4196
rect 1708 4132 1725 4196
rect 1789 4132 1806 4196
rect 1870 4132 1887 4196
rect 1951 4132 1968 4196
rect 2032 4132 2049 4196
rect 2113 4132 2130 4196
rect 2194 4132 2211 4196
rect 2275 4132 2292 4196
rect 2356 4132 2373 4196
rect 2437 4132 2454 4196
rect 2518 4132 2535 4196
rect 2599 4132 2616 4196
rect 2680 4132 2697 4196
rect 2761 4132 2778 4196
rect 2842 4132 2859 4196
rect 2923 4132 2940 4196
rect 3004 4132 3021 4196
rect 3085 4132 3102 4196
rect 3166 4132 3183 4196
rect 3247 4132 3264 4196
rect 3328 4132 3345 4196
rect 3409 4132 3426 4196
rect 3490 4132 3507 4196
rect 3571 4132 3588 4196
rect 3652 4132 3669 4196
rect 3733 4132 3750 4196
rect 3814 4132 3831 4196
rect 3895 4132 3912 4196
rect 3976 4132 3993 4196
rect 4057 4132 4074 4196
rect 4138 4132 4155 4196
rect 4219 4132 4236 4196
rect 4300 4132 4317 4196
rect 4381 4132 4399 4196
rect 4463 4132 4481 4196
rect 4545 4132 4563 4196
rect 4627 4132 4645 4196
rect 4709 4132 4727 4196
rect 4791 4132 4809 4196
rect 4873 4132 4879 4196
rect 99 4110 4879 4132
rect 99 4046 105 4110
rect 169 4046 186 4110
rect 250 4046 267 4110
rect 331 4046 348 4110
rect 412 4046 429 4110
rect 493 4046 510 4110
rect 574 4046 591 4110
rect 655 4046 672 4110
rect 736 4046 753 4110
rect 817 4046 834 4110
rect 898 4046 915 4110
rect 979 4046 996 4110
rect 1060 4046 1077 4110
rect 1141 4046 1158 4110
rect 1222 4046 1239 4110
rect 1303 4046 1320 4110
rect 1384 4046 1401 4110
rect 1465 4046 1482 4110
rect 1546 4046 1563 4110
rect 1627 4046 1644 4110
rect 1708 4046 1725 4110
rect 1789 4046 1806 4110
rect 1870 4046 1887 4110
rect 1951 4046 1968 4110
rect 2032 4046 2049 4110
rect 2113 4046 2130 4110
rect 2194 4046 2211 4110
rect 2275 4046 2292 4110
rect 2356 4046 2373 4110
rect 2437 4046 2454 4110
rect 2518 4046 2535 4110
rect 2599 4046 2616 4110
rect 2680 4046 2697 4110
rect 2761 4046 2778 4110
rect 2842 4046 2859 4110
rect 2923 4046 2940 4110
rect 3004 4046 3021 4110
rect 3085 4046 3102 4110
rect 3166 4046 3183 4110
rect 3247 4046 3264 4110
rect 3328 4046 3345 4110
rect 3409 4046 3426 4110
rect 3490 4046 3507 4110
rect 3571 4046 3588 4110
rect 3652 4046 3669 4110
rect 3733 4046 3750 4110
rect 3814 4046 3831 4110
rect 3895 4046 3912 4110
rect 3976 4046 3993 4110
rect 4057 4046 4074 4110
rect 4138 4046 4155 4110
rect 4219 4046 4236 4110
rect 4300 4046 4317 4110
rect 4381 4046 4399 4110
rect 4463 4046 4481 4110
rect 4545 4046 4563 4110
rect 4627 4046 4645 4110
rect 4709 4046 4727 4110
rect 4791 4046 4809 4110
rect 4873 4046 4879 4110
rect 99 4024 4879 4046
rect 99 3960 105 4024
rect 169 3960 186 4024
rect 250 3960 267 4024
rect 331 3960 348 4024
rect 412 3960 429 4024
rect 493 3960 510 4024
rect 574 3960 591 4024
rect 655 3960 672 4024
rect 736 3960 753 4024
rect 817 3960 834 4024
rect 898 3960 915 4024
rect 979 3960 996 4024
rect 1060 3960 1077 4024
rect 1141 3960 1158 4024
rect 1222 3960 1239 4024
rect 1303 3960 1320 4024
rect 1384 3960 1401 4024
rect 1465 3960 1482 4024
rect 1546 3960 1563 4024
rect 1627 3960 1644 4024
rect 1708 3960 1725 4024
rect 1789 3960 1806 4024
rect 1870 3960 1887 4024
rect 1951 3960 1968 4024
rect 2032 3960 2049 4024
rect 2113 3960 2130 4024
rect 2194 3960 2211 4024
rect 2275 3960 2292 4024
rect 2356 3960 2373 4024
rect 2437 3960 2454 4024
rect 2518 3960 2535 4024
rect 2599 3960 2616 4024
rect 2680 3960 2697 4024
rect 2761 3960 2778 4024
rect 2842 3960 2859 4024
rect 2923 3960 2940 4024
rect 3004 3960 3021 4024
rect 3085 3960 3102 4024
rect 3166 3960 3183 4024
rect 3247 3960 3264 4024
rect 3328 3960 3345 4024
rect 3409 3960 3426 4024
rect 3490 3960 3507 4024
rect 3571 3960 3588 4024
rect 3652 3960 3669 4024
rect 3733 3960 3750 4024
rect 3814 3960 3831 4024
rect 3895 3960 3912 4024
rect 3976 3960 3993 4024
rect 4057 3960 4074 4024
rect 4138 3960 4155 4024
rect 4219 3960 4236 4024
rect 4300 3960 4317 4024
rect 4381 3960 4399 4024
rect 4463 3960 4481 4024
rect 4545 3960 4563 4024
rect 4627 3960 4645 4024
rect 4709 3960 4727 4024
rect 4791 3960 4809 4024
rect 4873 3960 4879 4024
rect 99 3958 4879 3960
rect 10078 4884 14858 4886
rect 10078 4820 10084 4884
rect 10148 4820 10165 4884
rect 10229 4820 10246 4884
rect 10310 4820 10327 4884
rect 10391 4820 10408 4884
rect 10472 4820 10489 4884
rect 10553 4820 10570 4884
rect 10634 4820 10651 4884
rect 10715 4820 10732 4884
rect 10796 4820 10813 4884
rect 10877 4820 10894 4884
rect 10958 4820 10975 4884
rect 11039 4820 11056 4884
rect 11120 4820 11137 4884
rect 11201 4820 11218 4884
rect 11282 4820 11299 4884
rect 11363 4820 11380 4884
rect 11444 4820 11461 4884
rect 11525 4820 11542 4884
rect 11606 4820 11623 4884
rect 11687 4820 11704 4884
rect 11768 4820 11785 4884
rect 11849 4820 11866 4884
rect 11930 4820 11947 4884
rect 12011 4820 12028 4884
rect 12092 4820 12109 4884
rect 12173 4820 12190 4884
rect 12254 4820 12271 4884
rect 12335 4820 12352 4884
rect 12416 4820 12433 4884
rect 12497 4820 12514 4884
rect 12578 4820 12595 4884
rect 12659 4820 12676 4884
rect 12740 4820 12757 4884
rect 12821 4820 12838 4884
rect 12902 4820 12919 4884
rect 12983 4820 13000 4884
rect 13064 4820 13081 4884
rect 13145 4820 13162 4884
rect 13226 4820 13243 4884
rect 13307 4820 13324 4884
rect 13388 4820 13405 4884
rect 13469 4820 13486 4884
rect 13550 4820 13567 4884
rect 13631 4820 13648 4884
rect 13712 4820 13729 4884
rect 13793 4820 13810 4884
rect 13874 4820 13891 4884
rect 13955 4820 13972 4884
rect 14036 4820 14053 4884
rect 14117 4820 14134 4884
rect 14198 4820 14215 4884
rect 14279 4820 14296 4884
rect 14360 4820 14378 4884
rect 14442 4820 14460 4884
rect 14524 4820 14542 4884
rect 14606 4820 14624 4884
rect 14688 4820 14706 4884
rect 14770 4820 14788 4884
rect 14852 4820 14858 4884
rect 10078 4798 14858 4820
rect 10078 4734 10084 4798
rect 10148 4734 10165 4798
rect 10229 4734 10246 4798
rect 10310 4734 10327 4798
rect 10391 4734 10408 4798
rect 10472 4734 10489 4798
rect 10553 4734 10570 4798
rect 10634 4734 10651 4798
rect 10715 4734 10732 4798
rect 10796 4734 10813 4798
rect 10877 4734 10894 4798
rect 10958 4734 10975 4798
rect 11039 4734 11056 4798
rect 11120 4734 11137 4798
rect 11201 4734 11218 4798
rect 11282 4734 11299 4798
rect 11363 4734 11380 4798
rect 11444 4734 11461 4798
rect 11525 4734 11542 4798
rect 11606 4734 11623 4798
rect 11687 4734 11704 4798
rect 11768 4734 11785 4798
rect 11849 4734 11866 4798
rect 11930 4734 11947 4798
rect 12011 4734 12028 4798
rect 12092 4734 12109 4798
rect 12173 4734 12190 4798
rect 12254 4734 12271 4798
rect 12335 4734 12352 4798
rect 12416 4734 12433 4798
rect 12497 4734 12514 4798
rect 12578 4734 12595 4798
rect 12659 4734 12676 4798
rect 12740 4734 12757 4798
rect 12821 4734 12838 4798
rect 12902 4734 12919 4798
rect 12983 4734 13000 4798
rect 13064 4734 13081 4798
rect 13145 4734 13162 4798
rect 13226 4734 13243 4798
rect 13307 4734 13324 4798
rect 13388 4734 13405 4798
rect 13469 4734 13486 4798
rect 13550 4734 13567 4798
rect 13631 4734 13648 4798
rect 13712 4734 13729 4798
rect 13793 4734 13810 4798
rect 13874 4734 13891 4798
rect 13955 4734 13972 4798
rect 14036 4734 14053 4798
rect 14117 4734 14134 4798
rect 14198 4734 14215 4798
rect 14279 4734 14296 4798
rect 14360 4734 14378 4798
rect 14442 4734 14460 4798
rect 14524 4734 14542 4798
rect 14606 4734 14624 4798
rect 14688 4734 14706 4798
rect 14770 4734 14788 4798
rect 14852 4734 14858 4798
rect 10078 4712 14858 4734
rect 10078 4648 10084 4712
rect 10148 4648 10165 4712
rect 10229 4648 10246 4712
rect 10310 4648 10327 4712
rect 10391 4648 10408 4712
rect 10472 4648 10489 4712
rect 10553 4648 10570 4712
rect 10634 4648 10651 4712
rect 10715 4648 10732 4712
rect 10796 4648 10813 4712
rect 10877 4648 10894 4712
rect 10958 4648 10975 4712
rect 11039 4648 11056 4712
rect 11120 4648 11137 4712
rect 11201 4648 11218 4712
rect 11282 4648 11299 4712
rect 11363 4648 11380 4712
rect 11444 4648 11461 4712
rect 11525 4648 11542 4712
rect 11606 4648 11623 4712
rect 11687 4648 11704 4712
rect 11768 4648 11785 4712
rect 11849 4648 11866 4712
rect 11930 4648 11947 4712
rect 12011 4648 12028 4712
rect 12092 4648 12109 4712
rect 12173 4648 12190 4712
rect 12254 4648 12271 4712
rect 12335 4648 12352 4712
rect 12416 4648 12433 4712
rect 12497 4648 12514 4712
rect 12578 4648 12595 4712
rect 12659 4648 12676 4712
rect 12740 4648 12757 4712
rect 12821 4648 12838 4712
rect 12902 4648 12919 4712
rect 12983 4648 13000 4712
rect 13064 4648 13081 4712
rect 13145 4648 13162 4712
rect 13226 4648 13243 4712
rect 13307 4648 13324 4712
rect 13388 4648 13405 4712
rect 13469 4648 13486 4712
rect 13550 4648 13567 4712
rect 13631 4648 13648 4712
rect 13712 4648 13729 4712
rect 13793 4648 13810 4712
rect 13874 4648 13891 4712
rect 13955 4648 13972 4712
rect 14036 4648 14053 4712
rect 14117 4648 14134 4712
rect 14198 4648 14215 4712
rect 14279 4648 14296 4712
rect 14360 4648 14378 4712
rect 14442 4648 14460 4712
rect 14524 4648 14542 4712
rect 14606 4648 14624 4712
rect 14688 4648 14706 4712
rect 14770 4648 14788 4712
rect 14852 4648 14858 4712
rect 10078 4626 14858 4648
rect 10078 4562 10084 4626
rect 10148 4562 10165 4626
rect 10229 4562 10246 4626
rect 10310 4562 10327 4626
rect 10391 4562 10408 4626
rect 10472 4562 10489 4626
rect 10553 4562 10570 4626
rect 10634 4562 10651 4626
rect 10715 4562 10732 4626
rect 10796 4562 10813 4626
rect 10877 4562 10894 4626
rect 10958 4562 10975 4626
rect 11039 4562 11056 4626
rect 11120 4562 11137 4626
rect 11201 4562 11218 4626
rect 11282 4562 11299 4626
rect 11363 4562 11380 4626
rect 11444 4562 11461 4626
rect 11525 4562 11542 4626
rect 11606 4562 11623 4626
rect 11687 4562 11704 4626
rect 11768 4562 11785 4626
rect 11849 4562 11866 4626
rect 11930 4562 11947 4626
rect 12011 4562 12028 4626
rect 12092 4562 12109 4626
rect 12173 4562 12190 4626
rect 12254 4562 12271 4626
rect 12335 4562 12352 4626
rect 12416 4562 12433 4626
rect 12497 4562 12514 4626
rect 12578 4562 12595 4626
rect 12659 4562 12676 4626
rect 12740 4562 12757 4626
rect 12821 4562 12838 4626
rect 12902 4562 12919 4626
rect 12983 4562 13000 4626
rect 13064 4562 13081 4626
rect 13145 4562 13162 4626
rect 13226 4562 13243 4626
rect 13307 4562 13324 4626
rect 13388 4562 13405 4626
rect 13469 4562 13486 4626
rect 13550 4562 13567 4626
rect 13631 4562 13648 4626
rect 13712 4562 13729 4626
rect 13793 4562 13810 4626
rect 13874 4562 13891 4626
rect 13955 4562 13972 4626
rect 14036 4562 14053 4626
rect 14117 4562 14134 4626
rect 14198 4562 14215 4626
rect 14279 4562 14296 4626
rect 14360 4562 14378 4626
rect 14442 4562 14460 4626
rect 14524 4562 14542 4626
rect 14606 4562 14624 4626
rect 14688 4562 14706 4626
rect 14770 4562 14788 4626
rect 14852 4562 14858 4626
rect 10078 4540 14858 4562
rect 10078 4476 10084 4540
rect 10148 4476 10165 4540
rect 10229 4476 10246 4540
rect 10310 4476 10327 4540
rect 10391 4476 10408 4540
rect 10472 4476 10489 4540
rect 10553 4476 10570 4540
rect 10634 4476 10651 4540
rect 10715 4476 10732 4540
rect 10796 4476 10813 4540
rect 10877 4476 10894 4540
rect 10958 4476 10975 4540
rect 11039 4476 11056 4540
rect 11120 4476 11137 4540
rect 11201 4476 11218 4540
rect 11282 4476 11299 4540
rect 11363 4476 11380 4540
rect 11444 4476 11461 4540
rect 11525 4476 11542 4540
rect 11606 4476 11623 4540
rect 11687 4476 11704 4540
rect 11768 4476 11785 4540
rect 11849 4476 11866 4540
rect 11930 4476 11947 4540
rect 12011 4476 12028 4540
rect 12092 4476 12109 4540
rect 12173 4476 12190 4540
rect 12254 4476 12271 4540
rect 12335 4476 12352 4540
rect 12416 4476 12433 4540
rect 12497 4476 12514 4540
rect 12578 4476 12595 4540
rect 12659 4476 12676 4540
rect 12740 4476 12757 4540
rect 12821 4476 12838 4540
rect 12902 4476 12919 4540
rect 12983 4476 13000 4540
rect 13064 4476 13081 4540
rect 13145 4476 13162 4540
rect 13226 4476 13243 4540
rect 13307 4476 13324 4540
rect 13388 4476 13405 4540
rect 13469 4476 13486 4540
rect 13550 4476 13567 4540
rect 13631 4476 13648 4540
rect 13712 4476 13729 4540
rect 13793 4476 13810 4540
rect 13874 4476 13891 4540
rect 13955 4476 13972 4540
rect 14036 4476 14053 4540
rect 14117 4476 14134 4540
rect 14198 4476 14215 4540
rect 14279 4476 14296 4540
rect 14360 4476 14378 4540
rect 14442 4476 14460 4540
rect 14524 4476 14542 4540
rect 14606 4476 14624 4540
rect 14688 4476 14706 4540
rect 14770 4476 14788 4540
rect 14852 4476 14858 4540
rect 10078 4454 14858 4476
rect 10078 4390 10084 4454
rect 10148 4390 10165 4454
rect 10229 4390 10246 4454
rect 10310 4390 10327 4454
rect 10391 4390 10408 4454
rect 10472 4390 10489 4454
rect 10553 4390 10570 4454
rect 10634 4390 10651 4454
rect 10715 4390 10732 4454
rect 10796 4390 10813 4454
rect 10877 4390 10894 4454
rect 10958 4390 10975 4454
rect 11039 4390 11056 4454
rect 11120 4390 11137 4454
rect 11201 4390 11218 4454
rect 11282 4390 11299 4454
rect 11363 4390 11380 4454
rect 11444 4390 11461 4454
rect 11525 4390 11542 4454
rect 11606 4390 11623 4454
rect 11687 4390 11704 4454
rect 11768 4390 11785 4454
rect 11849 4390 11866 4454
rect 11930 4390 11947 4454
rect 12011 4390 12028 4454
rect 12092 4390 12109 4454
rect 12173 4390 12190 4454
rect 12254 4390 12271 4454
rect 12335 4390 12352 4454
rect 12416 4390 12433 4454
rect 12497 4390 12514 4454
rect 12578 4390 12595 4454
rect 12659 4390 12676 4454
rect 12740 4390 12757 4454
rect 12821 4390 12838 4454
rect 12902 4390 12919 4454
rect 12983 4390 13000 4454
rect 13064 4390 13081 4454
rect 13145 4390 13162 4454
rect 13226 4390 13243 4454
rect 13307 4390 13324 4454
rect 13388 4390 13405 4454
rect 13469 4390 13486 4454
rect 13550 4390 13567 4454
rect 13631 4390 13648 4454
rect 13712 4390 13729 4454
rect 13793 4390 13810 4454
rect 13874 4390 13891 4454
rect 13955 4390 13972 4454
rect 14036 4390 14053 4454
rect 14117 4390 14134 4454
rect 14198 4390 14215 4454
rect 14279 4390 14296 4454
rect 14360 4390 14378 4454
rect 14442 4390 14460 4454
rect 14524 4390 14542 4454
rect 14606 4390 14624 4454
rect 14688 4390 14706 4454
rect 14770 4390 14788 4454
rect 14852 4390 14858 4454
rect 10078 4368 14858 4390
rect 10078 4304 10084 4368
rect 10148 4304 10165 4368
rect 10229 4304 10246 4368
rect 10310 4304 10327 4368
rect 10391 4304 10408 4368
rect 10472 4304 10489 4368
rect 10553 4304 10570 4368
rect 10634 4304 10651 4368
rect 10715 4304 10732 4368
rect 10796 4304 10813 4368
rect 10877 4304 10894 4368
rect 10958 4304 10975 4368
rect 11039 4304 11056 4368
rect 11120 4304 11137 4368
rect 11201 4304 11218 4368
rect 11282 4304 11299 4368
rect 11363 4304 11380 4368
rect 11444 4304 11461 4368
rect 11525 4304 11542 4368
rect 11606 4304 11623 4368
rect 11687 4304 11704 4368
rect 11768 4304 11785 4368
rect 11849 4304 11866 4368
rect 11930 4304 11947 4368
rect 12011 4304 12028 4368
rect 12092 4304 12109 4368
rect 12173 4304 12190 4368
rect 12254 4304 12271 4368
rect 12335 4304 12352 4368
rect 12416 4304 12433 4368
rect 12497 4304 12514 4368
rect 12578 4304 12595 4368
rect 12659 4304 12676 4368
rect 12740 4304 12757 4368
rect 12821 4304 12838 4368
rect 12902 4304 12919 4368
rect 12983 4304 13000 4368
rect 13064 4304 13081 4368
rect 13145 4304 13162 4368
rect 13226 4304 13243 4368
rect 13307 4304 13324 4368
rect 13388 4304 13405 4368
rect 13469 4304 13486 4368
rect 13550 4304 13567 4368
rect 13631 4304 13648 4368
rect 13712 4304 13729 4368
rect 13793 4304 13810 4368
rect 13874 4304 13891 4368
rect 13955 4304 13972 4368
rect 14036 4304 14053 4368
rect 14117 4304 14134 4368
rect 14198 4304 14215 4368
rect 14279 4304 14296 4368
rect 14360 4304 14378 4368
rect 14442 4304 14460 4368
rect 14524 4304 14542 4368
rect 14606 4304 14624 4368
rect 14688 4304 14706 4368
rect 14770 4304 14788 4368
rect 14852 4304 14858 4368
rect 10078 4282 14858 4304
rect 10078 4218 10084 4282
rect 10148 4218 10165 4282
rect 10229 4218 10246 4282
rect 10310 4218 10327 4282
rect 10391 4218 10408 4282
rect 10472 4218 10489 4282
rect 10553 4218 10570 4282
rect 10634 4218 10651 4282
rect 10715 4218 10732 4282
rect 10796 4218 10813 4282
rect 10877 4218 10894 4282
rect 10958 4218 10975 4282
rect 11039 4218 11056 4282
rect 11120 4218 11137 4282
rect 11201 4218 11218 4282
rect 11282 4218 11299 4282
rect 11363 4218 11380 4282
rect 11444 4218 11461 4282
rect 11525 4218 11542 4282
rect 11606 4218 11623 4282
rect 11687 4218 11704 4282
rect 11768 4218 11785 4282
rect 11849 4218 11866 4282
rect 11930 4218 11947 4282
rect 12011 4218 12028 4282
rect 12092 4218 12109 4282
rect 12173 4218 12190 4282
rect 12254 4218 12271 4282
rect 12335 4218 12352 4282
rect 12416 4218 12433 4282
rect 12497 4218 12514 4282
rect 12578 4218 12595 4282
rect 12659 4218 12676 4282
rect 12740 4218 12757 4282
rect 12821 4218 12838 4282
rect 12902 4218 12919 4282
rect 12983 4218 13000 4282
rect 13064 4218 13081 4282
rect 13145 4218 13162 4282
rect 13226 4218 13243 4282
rect 13307 4218 13324 4282
rect 13388 4218 13405 4282
rect 13469 4218 13486 4282
rect 13550 4218 13567 4282
rect 13631 4218 13648 4282
rect 13712 4218 13729 4282
rect 13793 4218 13810 4282
rect 13874 4218 13891 4282
rect 13955 4218 13972 4282
rect 14036 4218 14053 4282
rect 14117 4218 14134 4282
rect 14198 4218 14215 4282
rect 14279 4218 14296 4282
rect 14360 4218 14378 4282
rect 14442 4218 14460 4282
rect 14524 4218 14542 4282
rect 14606 4218 14624 4282
rect 14688 4218 14706 4282
rect 14770 4218 14788 4282
rect 14852 4218 14858 4282
rect 10078 4196 14858 4218
rect 10078 4132 10084 4196
rect 10148 4132 10165 4196
rect 10229 4132 10246 4196
rect 10310 4132 10327 4196
rect 10391 4132 10408 4196
rect 10472 4132 10489 4196
rect 10553 4132 10570 4196
rect 10634 4132 10651 4196
rect 10715 4132 10732 4196
rect 10796 4132 10813 4196
rect 10877 4132 10894 4196
rect 10958 4132 10975 4196
rect 11039 4132 11056 4196
rect 11120 4132 11137 4196
rect 11201 4132 11218 4196
rect 11282 4132 11299 4196
rect 11363 4132 11380 4196
rect 11444 4132 11461 4196
rect 11525 4132 11542 4196
rect 11606 4132 11623 4196
rect 11687 4132 11704 4196
rect 11768 4132 11785 4196
rect 11849 4132 11866 4196
rect 11930 4132 11947 4196
rect 12011 4132 12028 4196
rect 12092 4132 12109 4196
rect 12173 4132 12190 4196
rect 12254 4132 12271 4196
rect 12335 4132 12352 4196
rect 12416 4132 12433 4196
rect 12497 4132 12514 4196
rect 12578 4132 12595 4196
rect 12659 4132 12676 4196
rect 12740 4132 12757 4196
rect 12821 4132 12838 4196
rect 12902 4132 12919 4196
rect 12983 4132 13000 4196
rect 13064 4132 13081 4196
rect 13145 4132 13162 4196
rect 13226 4132 13243 4196
rect 13307 4132 13324 4196
rect 13388 4132 13405 4196
rect 13469 4132 13486 4196
rect 13550 4132 13567 4196
rect 13631 4132 13648 4196
rect 13712 4132 13729 4196
rect 13793 4132 13810 4196
rect 13874 4132 13891 4196
rect 13955 4132 13972 4196
rect 14036 4132 14053 4196
rect 14117 4132 14134 4196
rect 14198 4132 14215 4196
rect 14279 4132 14296 4196
rect 14360 4132 14378 4196
rect 14442 4132 14460 4196
rect 14524 4132 14542 4196
rect 14606 4132 14624 4196
rect 14688 4132 14706 4196
rect 14770 4132 14788 4196
rect 14852 4132 14858 4196
rect 10078 4110 14858 4132
rect 10078 4046 10084 4110
rect 10148 4046 10165 4110
rect 10229 4046 10246 4110
rect 10310 4046 10327 4110
rect 10391 4046 10408 4110
rect 10472 4046 10489 4110
rect 10553 4046 10570 4110
rect 10634 4046 10651 4110
rect 10715 4046 10732 4110
rect 10796 4046 10813 4110
rect 10877 4046 10894 4110
rect 10958 4046 10975 4110
rect 11039 4046 11056 4110
rect 11120 4046 11137 4110
rect 11201 4046 11218 4110
rect 11282 4046 11299 4110
rect 11363 4046 11380 4110
rect 11444 4046 11461 4110
rect 11525 4046 11542 4110
rect 11606 4046 11623 4110
rect 11687 4046 11704 4110
rect 11768 4046 11785 4110
rect 11849 4046 11866 4110
rect 11930 4046 11947 4110
rect 12011 4046 12028 4110
rect 12092 4046 12109 4110
rect 12173 4046 12190 4110
rect 12254 4046 12271 4110
rect 12335 4046 12352 4110
rect 12416 4046 12433 4110
rect 12497 4046 12514 4110
rect 12578 4046 12595 4110
rect 12659 4046 12676 4110
rect 12740 4046 12757 4110
rect 12821 4046 12838 4110
rect 12902 4046 12919 4110
rect 12983 4046 13000 4110
rect 13064 4046 13081 4110
rect 13145 4046 13162 4110
rect 13226 4046 13243 4110
rect 13307 4046 13324 4110
rect 13388 4046 13405 4110
rect 13469 4046 13486 4110
rect 13550 4046 13567 4110
rect 13631 4046 13648 4110
rect 13712 4046 13729 4110
rect 13793 4046 13810 4110
rect 13874 4046 13891 4110
rect 13955 4046 13972 4110
rect 14036 4046 14053 4110
rect 14117 4046 14134 4110
rect 14198 4046 14215 4110
rect 14279 4046 14296 4110
rect 14360 4046 14378 4110
rect 14442 4046 14460 4110
rect 14524 4046 14542 4110
rect 14606 4046 14624 4110
rect 14688 4046 14706 4110
rect 14770 4046 14788 4110
rect 14852 4046 14858 4110
rect 10078 4024 14858 4046
rect 10078 3960 10084 4024
rect 10148 3960 10165 4024
rect 10229 3960 10246 4024
rect 10310 3960 10327 4024
rect 10391 3960 10408 4024
rect 10472 3960 10489 4024
rect 10553 3960 10570 4024
rect 10634 3960 10651 4024
rect 10715 3960 10732 4024
rect 10796 3960 10813 4024
rect 10877 3960 10894 4024
rect 10958 3960 10975 4024
rect 11039 3960 11056 4024
rect 11120 3960 11137 4024
rect 11201 3960 11218 4024
rect 11282 3960 11299 4024
rect 11363 3960 11380 4024
rect 11444 3960 11461 4024
rect 11525 3960 11542 4024
rect 11606 3960 11623 4024
rect 11687 3960 11704 4024
rect 11768 3960 11785 4024
rect 11849 3960 11866 4024
rect 11930 3960 11947 4024
rect 12011 3960 12028 4024
rect 12092 3960 12109 4024
rect 12173 3960 12190 4024
rect 12254 3960 12271 4024
rect 12335 3960 12352 4024
rect 12416 3960 12433 4024
rect 12497 3960 12514 4024
rect 12578 3960 12595 4024
rect 12659 3960 12676 4024
rect 12740 3960 12757 4024
rect 12821 3960 12838 4024
rect 12902 3960 12919 4024
rect 12983 3960 13000 4024
rect 13064 3960 13081 4024
rect 13145 3960 13162 4024
rect 13226 3960 13243 4024
rect 13307 3960 13324 4024
rect 13388 3960 13405 4024
rect 13469 3960 13486 4024
rect 13550 3960 13567 4024
rect 13631 3960 13648 4024
rect 13712 3960 13729 4024
rect 13793 3960 13810 4024
rect 13874 3960 13891 4024
rect 13955 3960 13972 4024
rect 14036 3960 14053 4024
rect 14117 3960 14134 4024
rect 14198 3960 14215 4024
rect 14279 3960 14296 4024
rect 14360 3960 14378 4024
rect 14442 3960 14460 4024
rect 14524 3960 14542 4024
rect 14606 3960 14624 4024
rect 14688 3960 14706 4024
rect 14770 3960 14788 4024
rect 14852 3960 14858 4024
rect 10078 3958 14858 3960
<< via3 >>
rect 162 18886 226 18950
rect 243 18886 307 18950
rect 324 18886 388 18950
rect 405 18886 469 18950
rect 486 18886 550 18950
rect 567 18886 631 18950
rect 648 18886 712 18950
rect 729 18886 793 18950
rect 810 18886 874 18950
rect 891 18886 955 18950
rect 972 18886 1036 18950
rect 1053 18886 1117 18950
rect 1134 18886 1198 18950
rect 1215 18886 1279 18950
rect 1296 18886 1360 18950
rect 1377 18886 1441 18950
rect 1458 18886 1522 18950
rect 1539 18886 1603 18950
rect 1620 18886 1684 18950
rect 1701 18886 1765 18950
rect 1782 18886 1846 18950
rect 1863 18886 1927 18950
rect 1944 18886 2008 18950
rect 2025 18886 2089 18950
rect 2106 18886 2170 18950
rect 2187 18886 2251 18950
rect 2268 18886 2332 18950
rect 2349 18886 2413 18950
rect 2430 18886 2494 18950
rect 2511 18886 2575 18950
rect 2592 18886 2656 18950
rect 2673 18886 2737 18950
rect 2754 18886 2818 18950
rect 2835 18886 2899 18950
rect 2916 18886 2980 18950
rect 2997 18886 3061 18950
rect 3078 18886 3142 18950
rect 3159 18886 3223 18950
rect 3240 18886 3304 18950
rect 3321 18886 3385 18950
rect 3402 18886 3466 18950
rect 3483 18886 3547 18950
rect 3563 18886 3627 18950
rect 3643 18886 3707 18950
rect 3723 18886 3787 18950
rect 3803 18886 3867 18950
rect 3883 18886 3947 18950
rect 162 18802 226 18866
rect 243 18802 307 18866
rect 324 18802 388 18866
rect 405 18802 469 18866
rect 486 18802 550 18866
rect 567 18802 631 18866
rect 648 18802 712 18866
rect 729 18802 793 18866
rect 810 18802 874 18866
rect 891 18802 955 18866
rect 972 18802 1036 18866
rect 1053 18802 1117 18866
rect 1134 18802 1198 18866
rect 1215 18802 1279 18866
rect 1296 18802 1360 18866
rect 1377 18802 1441 18866
rect 1458 18802 1522 18866
rect 1539 18802 1603 18866
rect 1620 18802 1684 18866
rect 1701 18802 1765 18866
rect 1782 18802 1846 18866
rect 1863 18802 1927 18866
rect 1944 18802 2008 18866
rect 2025 18802 2089 18866
rect 2106 18802 2170 18866
rect 2187 18802 2251 18866
rect 2268 18802 2332 18866
rect 2349 18802 2413 18866
rect 2430 18802 2494 18866
rect 2511 18802 2575 18866
rect 2592 18802 2656 18866
rect 2673 18802 2737 18866
rect 2754 18802 2818 18866
rect 2835 18802 2899 18866
rect 2916 18802 2980 18866
rect 2997 18802 3061 18866
rect 3078 18802 3142 18866
rect 3159 18802 3223 18866
rect 3240 18802 3304 18866
rect 3321 18802 3385 18866
rect 3402 18802 3466 18866
rect 3483 18802 3547 18866
rect 3563 18802 3627 18866
rect 3643 18802 3707 18866
rect 3723 18802 3787 18866
rect 3803 18802 3867 18866
rect 3883 18802 3947 18866
rect 162 18718 226 18782
rect 243 18718 307 18782
rect 324 18718 388 18782
rect 405 18718 469 18782
rect 486 18718 550 18782
rect 567 18718 631 18782
rect 648 18718 712 18782
rect 729 18718 793 18782
rect 810 18718 874 18782
rect 891 18718 955 18782
rect 972 18718 1036 18782
rect 1053 18718 1117 18782
rect 1134 18718 1198 18782
rect 1215 18718 1279 18782
rect 1296 18718 1360 18782
rect 1377 18718 1441 18782
rect 1458 18718 1522 18782
rect 1539 18718 1603 18782
rect 1620 18718 1684 18782
rect 1701 18718 1765 18782
rect 1782 18718 1846 18782
rect 1863 18718 1927 18782
rect 1944 18718 2008 18782
rect 2025 18718 2089 18782
rect 2106 18718 2170 18782
rect 2187 18718 2251 18782
rect 2268 18718 2332 18782
rect 2349 18718 2413 18782
rect 2430 18718 2494 18782
rect 2511 18718 2575 18782
rect 2592 18718 2656 18782
rect 2673 18718 2737 18782
rect 2754 18718 2818 18782
rect 2835 18718 2899 18782
rect 2916 18718 2980 18782
rect 2997 18718 3061 18782
rect 3078 18718 3142 18782
rect 3159 18718 3223 18782
rect 3240 18718 3304 18782
rect 3321 18718 3385 18782
rect 3402 18718 3466 18782
rect 3483 18718 3547 18782
rect 3563 18718 3627 18782
rect 3643 18718 3707 18782
rect 3723 18718 3787 18782
rect 3803 18718 3867 18782
rect 3883 18718 3947 18782
rect 11065 18886 11129 18950
rect 11145 18886 11209 18950
rect 11225 18886 11289 18950
rect 11305 18886 11369 18950
rect 11385 18886 11449 18950
rect 11465 18886 11529 18950
rect 11546 18886 11610 18950
rect 11627 18886 11691 18950
rect 11708 18886 11772 18950
rect 11789 18886 11853 18950
rect 11870 18886 11934 18950
rect 11951 18886 12015 18950
rect 12032 18886 12096 18950
rect 12113 18886 12177 18950
rect 12194 18886 12258 18950
rect 12275 18886 12339 18950
rect 12356 18886 12420 18950
rect 12437 18886 12501 18950
rect 12518 18886 12582 18950
rect 12599 18886 12663 18950
rect 12680 18886 12744 18950
rect 12761 18886 12825 18950
rect 12842 18886 12906 18950
rect 12923 18886 12987 18950
rect 13004 18886 13068 18950
rect 13085 18886 13149 18950
rect 13166 18886 13230 18950
rect 13247 18886 13311 18950
rect 13328 18886 13392 18950
rect 13409 18886 13473 18950
rect 13490 18886 13554 18950
rect 13571 18886 13635 18950
rect 13652 18886 13716 18950
rect 13733 18886 13797 18950
rect 13814 18886 13878 18950
rect 13895 18886 13959 18950
rect 13976 18886 14040 18950
rect 14057 18886 14121 18950
rect 14138 18886 14202 18950
rect 14219 18886 14283 18950
rect 14300 18886 14364 18950
rect 14381 18886 14445 18950
rect 14462 18886 14526 18950
rect 14543 18886 14607 18950
rect 14624 18886 14688 18950
rect 14705 18886 14769 18950
rect 14786 18886 14850 18950
rect 11065 18802 11129 18866
rect 11145 18802 11209 18866
rect 11225 18802 11289 18866
rect 11305 18802 11369 18866
rect 11385 18802 11449 18866
rect 11465 18802 11529 18866
rect 11546 18802 11610 18866
rect 11627 18802 11691 18866
rect 11708 18802 11772 18866
rect 11789 18802 11853 18866
rect 11870 18802 11934 18866
rect 11951 18802 12015 18866
rect 12032 18802 12096 18866
rect 12113 18802 12177 18866
rect 12194 18802 12258 18866
rect 12275 18802 12339 18866
rect 12356 18802 12420 18866
rect 12437 18802 12501 18866
rect 12518 18802 12582 18866
rect 12599 18802 12663 18866
rect 12680 18802 12744 18866
rect 12761 18802 12825 18866
rect 12842 18802 12906 18866
rect 12923 18802 12987 18866
rect 13004 18802 13068 18866
rect 13085 18802 13149 18866
rect 13166 18802 13230 18866
rect 13247 18802 13311 18866
rect 13328 18802 13392 18866
rect 13409 18802 13473 18866
rect 13490 18802 13554 18866
rect 13571 18802 13635 18866
rect 13652 18802 13716 18866
rect 13733 18802 13797 18866
rect 13814 18802 13878 18866
rect 13895 18802 13959 18866
rect 13976 18802 14040 18866
rect 14057 18802 14121 18866
rect 14138 18802 14202 18866
rect 14219 18802 14283 18866
rect 14300 18802 14364 18866
rect 14381 18802 14445 18866
rect 14462 18802 14526 18866
rect 14543 18802 14607 18866
rect 14624 18802 14688 18866
rect 14705 18802 14769 18866
rect 14786 18802 14850 18866
rect 3994 18701 4058 18765
rect 4124 18701 4188 18765
rect 162 18634 226 18698
rect 243 18634 307 18698
rect 324 18634 388 18698
rect 405 18634 469 18698
rect 486 18634 550 18698
rect 567 18634 631 18698
rect 648 18634 712 18698
rect 729 18634 793 18698
rect 810 18634 874 18698
rect 891 18634 955 18698
rect 972 18634 1036 18698
rect 1053 18634 1117 18698
rect 1134 18634 1198 18698
rect 1215 18634 1279 18698
rect 1296 18634 1360 18698
rect 1377 18634 1441 18698
rect 1458 18634 1522 18698
rect 1539 18634 1603 18698
rect 1620 18634 1684 18698
rect 1701 18634 1765 18698
rect 1782 18634 1846 18698
rect 1863 18634 1927 18698
rect 1944 18634 2008 18698
rect 2025 18634 2089 18698
rect 2106 18634 2170 18698
rect 2187 18634 2251 18698
rect 2268 18634 2332 18698
rect 2349 18634 2413 18698
rect 2430 18634 2494 18698
rect 2511 18634 2575 18698
rect 2592 18634 2656 18698
rect 2673 18634 2737 18698
rect 2754 18634 2818 18698
rect 2835 18634 2899 18698
rect 2916 18634 2980 18698
rect 2997 18634 3061 18698
rect 3078 18634 3142 18698
rect 3159 18634 3223 18698
rect 3240 18634 3304 18698
rect 3321 18634 3385 18698
rect 3402 18634 3466 18698
rect 3483 18634 3547 18698
rect 3563 18634 3627 18698
rect 3643 18634 3707 18698
rect 3723 18634 3787 18698
rect 3803 18634 3867 18698
rect 3883 18634 3947 18698
rect 162 18550 226 18614
rect 243 18550 307 18614
rect 324 18550 388 18614
rect 405 18550 469 18614
rect 486 18550 550 18614
rect 567 18550 631 18614
rect 648 18550 712 18614
rect 729 18550 793 18614
rect 810 18550 874 18614
rect 891 18550 955 18614
rect 972 18550 1036 18614
rect 1053 18550 1117 18614
rect 1134 18550 1198 18614
rect 1215 18550 1279 18614
rect 1296 18550 1360 18614
rect 1377 18550 1441 18614
rect 1458 18550 1522 18614
rect 1539 18550 1603 18614
rect 1620 18550 1684 18614
rect 1701 18550 1765 18614
rect 1782 18550 1846 18614
rect 1863 18550 1927 18614
rect 1944 18550 2008 18614
rect 2025 18550 2089 18614
rect 2106 18550 2170 18614
rect 2187 18550 2251 18614
rect 2268 18550 2332 18614
rect 2349 18550 2413 18614
rect 2430 18550 2494 18614
rect 2511 18550 2575 18614
rect 2592 18550 2656 18614
rect 2673 18550 2737 18614
rect 2754 18550 2818 18614
rect 2835 18550 2899 18614
rect 2916 18550 2980 18614
rect 2997 18550 3061 18614
rect 3078 18550 3142 18614
rect 3159 18550 3223 18614
rect 3240 18550 3304 18614
rect 3321 18550 3385 18614
rect 3402 18550 3466 18614
rect 3483 18550 3547 18614
rect 3563 18550 3627 18614
rect 3643 18550 3707 18614
rect 3723 18550 3787 18614
rect 3803 18550 3867 18614
rect 3883 18550 3947 18614
rect 3994 18579 4058 18643
rect 4124 18579 4188 18643
rect 10824 18701 10888 18765
rect 10954 18701 11018 18765
rect 11065 18718 11129 18782
rect 11145 18718 11209 18782
rect 11225 18718 11289 18782
rect 11305 18718 11369 18782
rect 11385 18718 11449 18782
rect 11465 18718 11529 18782
rect 11546 18718 11610 18782
rect 11627 18718 11691 18782
rect 11708 18718 11772 18782
rect 11789 18718 11853 18782
rect 11870 18718 11934 18782
rect 11951 18718 12015 18782
rect 12032 18718 12096 18782
rect 12113 18718 12177 18782
rect 12194 18718 12258 18782
rect 12275 18718 12339 18782
rect 12356 18718 12420 18782
rect 12437 18718 12501 18782
rect 12518 18718 12582 18782
rect 12599 18718 12663 18782
rect 12680 18718 12744 18782
rect 12761 18718 12825 18782
rect 12842 18718 12906 18782
rect 12923 18718 12987 18782
rect 13004 18718 13068 18782
rect 13085 18718 13149 18782
rect 13166 18718 13230 18782
rect 13247 18718 13311 18782
rect 13328 18718 13392 18782
rect 13409 18718 13473 18782
rect 13490 18718 13554 18782
rect 13571 18718 13635 18782
rect 13652 18718 13716 18782
rect 13733 18718 13797 18782
rect 13814 18718 13878 18782
rect 13895 18718 13959 18782
rect 13976 18718 14040 18782
rect 14057 18718 14121 18782
rect 14138 18718 14202 18782
rect 14219 18718 14283 18782
rect 14300 18718 14364 18782
rect 14381 18718 14445 18782
rect 14462 18718 14526 18782
rect 14543 18718 14607 18782
rect 14624 18718 14688 18782
rect 14705 18718 14769 18782
rect 14786 18718 14850 18782
rect 10824 18579 10888 18643
rect 10954 18579 11018 18643
rect 11065 18634 11129 18698
rect 11145 18634 11209 18698
rect 11225 18634 11289 18698
rect 11305 18634 11369 18698
rect 11385 18634 11449 18698
rect 11465 18634 11529 18698
rect 11546 18634 11610 18698
rect 11627 18634 11691 18698
rect 11708 18634 11772 18698
rect 11789 18634 11853 18698
rect 11870 18634 11934 18698
rect 11951 18634 12015 18698
rect 12032 18634 12096 18698
rect 12113 18634 12177 18698
rect 12194 18634 12258 18698
rect 12275 18634 12339 18698
rect 12356 18634 12420 18698
rect 12437 18634 12501 18698
rect 12518 18634 12582 18698
rect 12599 18634 12663 18698
rect 12680 18634 12744 18698
rect 12761 18634 12825 18698
rect 12842 18634 12906 18698
rect 12923 18634 12987 18698
rect 13004 18634 13068 18698
rect 13085 18634 13149 18698
rect 13166 18634 13230 18698
rect 13247 18634 13311 18698
rect 13328 18634 13392 18698
rect 13409 18634 13473 18698
rect 13490 18634 13554 18698
rect 13571 18634 13635 18698
rect 13652 18634 13716 18698
rect 13733 18634 13797 18698
rect 13814 18634 13878 18698
rect 13895 18634 13959 18698
rect 13976 18634 14040 18698
rect 14057 18634 14121 18698
rect 14138 18634 14202 18698
rect 14219 18634 14283 18698
rect 14300 18634 14364 18698
rect 14381 18634 14445 18698
rect 14462 18634 14526 18698
rect 14543 18634 14607 18698
rect 14624 18634 14688 18698
rect 14705 18634 14769 18698
rect 14786 18634 14850 18698
rect 162 18466 226 18530
rect 243 18466 307 18530
rect 324 18466 388 18530
rect 405 18466 469 18530
rect 486 18466 550 18530
rect 567 18466 631 18530
rect 648 18466 712 18530
rect 729 18466 793 18530
rect 810 18466 874 18530
rect 891 18466 955 18530
rect 972 18466 1036 18530
rect 1053 18466 1117 18530
rect 1134 18466 1198 18530
rect 1215 18466 1279 18530
rect 1296 18466 1360 18530
rect 1377 18466 1441 18530
rect 1458 18466 1522 18530
rect 1539 18466 1603 18530
rect 1620 18466 1684 18530
rect 1701 18466 1765 18530
rect 1782 18466 1846 18530
rect 1863 18466 1927 18530
rect 1944 18466 2008 18530
rect 2025 18466 2089 18530
rect 2106 18466 2170 18530
rect 2187 18466 2251 18530
rect 2268 18466 2332 18530
rect 2349 18466 2413 18530
rect 2430 18466 2494 18530
rect 2511 18466 2575 18530
rect 2592 18466 2656 18530
rect 2673 18466 2737 18530
rect 2754 18466 2818 18530
rect 2835 18466 2899 18530
rect 2916 18466 2980 18530
rect 2997 18466 3061 18530
rect 3078 18466 3142 18530
rect 3159 18466 3223 18530
rect 3240 18466 3304 18530
rect 3321 18466 3385 18530
rect 3402 18466 3466 18530
rect 3483 18466 3547 18530
rect 3563 18466 3627 18530
rect 3643 18466 3707 18530
rect 3723 18466 3787 18530
rect 3803 18466 3867 18530
rect 3883 18466 3947 18530
rect 11065 18550 11129 18614
rect 11145 18550 11209 18614
rect 11225 18550 11289 18614
rect 11305 18550 11369 18614
rect 11385 18550 11449 18614
rect 11465 18550 11529 18614
rect 11546 18550 11610 18614
rect 11627 18550 11691 18614
rect 11708 18550 11772 18614
rect 11789 18550 11853 18614
rect 11870 18550 11934 18614
rect 11951 18550 12015 18614
rect 12032 18550 12096 18614
rect 12113 18550 12177 18614
rect 12194 18550 12258 18614
rect 12275 18550 12339 18614
rect 12356 18550 12420 18614
rect 12437 18550 12501 18614
rect 12518 18550 12582 18614
rect 12599 18550 12663 18614
rect 12680 18550 12744 18614
rect 12761 18550 12825 18614
rect 12842 18550 12906 18614
rect 12923 18550 12987 18614
rect 13004 18550 13068 18614
rect 13085 18550 13149 18614
rect 13166 18550 13230 18614
rect 13247 18550 13311 18614
rect 13328 18550 13392 18614
rect 13409 18550 13473 18614
rect 13490 18550 13554 18614
rect 13571 18550 13635 18614
rect 13652 18550 13716 18614
rect 13733 18550 13797 18614
rect 13814 18550 13878 18614
rect 13895 18550 13959 18614
rect 13976 18550 14040 18614
rect 14057 18550 14121 18614
rect 14138 18550 14202 18614
rect 14219 18550 14283 18614
rect 14300 18550 14364 18614
rect 14381 18550 14445 18614
rect 14462 18550 14526 18614
rect 14543 18550 14607 18614
rect 14624 18550 14688 18614
rect 14705 18550 14769 18614
rect 14786 18550 14850 18614
rect 4016 18448 4080 18512
rect 4129 18448 4193 18512
rect 4242 18448 4306 18512
rect 4355 18448 4419 18512
rect 162 18382 226 18446
rect 243 18382 307 18446
rect 324 18382 388 18446
rect 405 18382 469 18446
rect 486 18382 550 18446
rect 567 18382 631 18446
rect 648 18382 712 18446
rect 729 18382 793 18446
rect 810 18382 874 18446
rect 891 18382 955 18446
rect 972 18382 1036 18446
rect 1053 18382 1117 18446
rect 1134 18382 1198 18446
rect 1215 18382 1279 18446
rect 1296 18382 1360 18446
rect 1377 18382 1441 18446
rect 1458 18382 1522 18446
rect 1539 18382 1603 18446
rect 1620 18382 1684 18446
rect 1701 18382 1765 18446
rect 1782 18382 1846 18446
rect 1863 18382 1927 18446
rect 1944 18382 2008 18446
rect 2025 18382 2089 18446
rect 2106 18382 2170 18446
rect 2187 18382 2251 18446
rect 2268 18382 2332 18446
rect 2349 18382 2413 18446
rect 2430 18382 2494 18446
rect 2511 18382 2575 18446
rect 2592 18382 2656 18446
rect 2673 18382 2737 18446
rect 2754 18382 2818 18446
rect 2835 18382 2899 18446
rect 2916 18382 2980 18446
rect 2997 18382 3061 18446
rect 3078 18382 3142 18446
rect 3159 18382 3223 18446
rect 3240 18382 3304 18446
rect 3321 18382 3385 18446
rect 3402 18382 3466 18446
rect 3483 18382 3547 18446
rect 3563 18382 3627 18446
rect 3643 18382 3707 18446
rect 3723 18382 3787 18446
rect 3803 18382 3867 18446
rect 3883 18382 3947 18446
rect 162 18298 226 18362
rect 243 18298 307 18362
rect 324 18298 388 18362
rect 405 18298 469 18362
rect 486 18298 550 18362
rect 567 18298 631 18362
rect 648 18298 712 18362
rect 729 18298 793 18362
rect 810 18298 874 18362
rect 891 18298 955 18362
rect 972 18298 1036 18362
rect 1053 18298 1117 18362
rect 1134 18298 1198 18362
rect 1215 18298 1279 18362
rect 1296 18298 1360 18362
rect 1377 18298 1441 18362
rect 1458 18298 1522 18362
rect 1539 18298 1603 18362
rect 1620 18298 1684 18362
rect 1701 18298 1765 18362
rect 1782 18298 1846 18362
rect 1863 18298 1927 18362
rect 1944 18298 2008 18362
rect 2025 18298 2089 18362
rect 2106 18298 2170 18362
rect 2187 18298 2251 18362
rect 2268 18298 2332 18362
rect 2349 18298 2413 18362
rect 2430 18298 2494 18362
rect 2511 18298 2575 18362
rect 2592 18298 2656 18362
rect 2673 18298 2737 18362
rect 2754 18298 2818 18362
rect 2835 18298 2899 18362
rect 2916 18298 2980 18362
rect 2997 18298 3061 18362
rect 3078 18298 3142 18362
rect 3159 18298 3223 18362
rect 3240 18298 3304 18362
rect 3321 18298 3385 18362
rect 3402 18298 3466 18362
rect 3483 18298 3547 18362
rect 3563 18298 3627 18362
rect 3643 18298 3707 18362
rect 3723 18298 3787 18362
rect 3803 18298 3867 18362
rect 3883 18298 3947 18362
rect 4016 18346 4080 18410
rect 4129 18346 4193 18410
rect 4242 18346 4306 18410
rect 4355 18346 4419 18410
rect 162 18214 226 18278
rect 243 18214 307 18278
rect 324 18214 388 18278
rect 405 18214 469 18278
rect 486 18214 550 18278
rect 567 18214 631 18278
rect 648 18214 712 18278
rect 729 18214 793 18278
rect 810 18214 874 18278
rect 891 18214 955 18278
rect 972 18214 1036 18278
rect 1053 18214 1117 18278
rect 1134 18214 1198 18278
rect 1215 18214 1279 18278
rect 1296 18214 1360 18278
rect 1377 18214 1441 18278
rect 1458 18214 1522 18278
rect 1539 18214 1603 18278
rect 1620 18214 1684 18278
rect 1701 18214 1765 18278
rect 1782 18214 1846 18278
rect 1863 18214 1927 18278
rect 1944 18214 2008 18278
rect 2025 18214 2089 18278
rect 2106 18214 2170 18278
rect 2187 18214 2251 18278
rect 2268 18214 2332 18278
rect 2349 18214 2413 18278
rect 2430 18214 2494 18278
rect 2511 18214 2575 18278
rect 2592 18214 2656 18278
rect 2673 18214 2737 18278
rect 2754 18214 2818 18278
rect 2835 18214 2899 18278
rect 2916 18214 2980 18278
rect 2997 18214 3061 18278
rect 3078 18214 3142 18278
rect 3159 18214 3223 18278
rect 3240 18214 3304 18278
rect 3321 18214 3385 18278
rect 3402 18214 3466 18278
rect 3483 18214 3547 18278
rect 3563 18214 3627 18278
rect 3643 18214 3707 18278
rect 3723 18214 3787 18278
rect 3803 18214 3867 18278
rect 3883 18214 3947 18278
rect 4016 18244 4080 18308
rect 4129 18244 4193 18308
rect 4242 18244 4306 18308
rect 4355 18244 4419 18308
rect 10593 18448 10657 18512
rect 10706 18448 10770 18512
rect 10819 18448 10883 18512
rect 10932 18448 10996 18512
rect 11065 18466 11129 18530
rect 11145 18466 11209 18530
rect 11225 18466 11289 18530
rect 11305 18466 11369 18530
rect 11385 18466 11449 18530
rect 11465 18466 11529 18530
rect 11546 18466 11610 18530
rect 11627 18466 11691 18530
rect 11708 18466 11772 18530
rect 11789 18466 11853 18530
rect 11870 18466 11934 18530
rect 11951 18466 12015 18530
rect 12032 18466 12096 18530
rect 12113 18466 12177 18530
rect 12194 18466 12258 18530
rect 12275 18466 12339 18530
rect 12356 18466 12420 18530
rect 12437 18466 12501 18530
rect 12518 18466 12582 18530
rect 12599 18466 12663 18530
rect 12680 18466 12744 18530
rect 12761 18466 12825 18530
rect 12842 18466 12906 18530
rect 12923 18466 12987 18530
rect 13004 18466 13068 18530
rect 13085 18466 13149 18530
rect 13166 18466 13230 18530
rect 13247 18466 13311 18530
rect 13328 18466 13392 18530
rect 13409 18466 13473 18530
rect 13490 18466 13554 18530
rect 13571 18466 13635 18530
rect 13652 18466 13716 18530
rect 13733 18466 13797 18530
rect 13814 18466 13878 18530
rect 13895 18466 13959 18530
rect 13976 18466 14040 18530
rect 14057 18466 14121 18530
rect 14138 18466 14202 18530
rect 14219 18466 14283 18530
rect 14300 18466 14364 18530
rect 14381 18466 14445 18530
rect 14462 18466 14526 18530
rect 14543 18466 14607 18530
rect 14624 18466 14688 18530
rect 14705 18466 14769 18530
rect 14786 18466 14850 18530
rect 10593 18346 10657 18410
rect 10706 18346 10770 18410
rect 10819 18346 10883 18410
rect 10932 18346 10996 18410
rect 11065 18382 11129 18446
rect 11145 18382 11209 18446
rect 11225 18382 11289 18446
rect 11305 18382 11369 18446
rect 11385 18382 11449 18446
rect 11465 18382 11529 18446
rect 11546 18382 11610 18446
rect 11627 18382 11691 18446
rect 11708 18382 11772 18446
rect 11789 18382 11853 18446
rect 11870 18382 11934 18446
rect 11951 18382 12015 18446
rect 12032 18382 12096 18446
rect 12113 18382 12177 18446
rect 12194 18382 12258 18446
rect 12275 18382 12339 18446
rect 12356 18382 12420 18446
rect 12437 18382 12501 18446
rect 12518 18382 12582 18446
rect 12599 18382 12663 18446
rect 12680 18382 12744 18446
rect 12761 18382 12825 18446
rect 12842 18382 12906 18446
rect 12923 18382 12987 18446
rect 13004 18382 13068 18446
rect 13085 18382 13149 18446
rect 13166 18382 13230 18446
rect 13247 18382 13311 18446
rect 13328 18382 13392 18446
rect 13409 18382 13473 18446
rect 13490 18382 13554 18446
rect 13571 18382 13635 18446
rect 13652 18382 13716 18446
rect 13733 18382 13797 18446
rect 13814 18382 13878 18446
rect 13895 18382 13959 18446
rect 13976 18382 14040 18446
rect 14057 18382 14121 18446
rect 14138 18382 14202 18446
rect 14219 18382 14283 18446
rect 14300 18382 14364 18446
rect 14381 18382 14445 18446
rect 14462 18382 14526 18446
rect 14543 18382 14607 18446
rect 14624 18382 14688 18446
rect 14705 18382 14769 18446
rect 14786 18382 14850 18446
rect 4478 18233 4542 18297
rect 4598 18233 4662 18297
rect 162 18130 226 18194
rect 243 18130 307 18194
rect 324 18130 388 18194
rect 405 18130 469 18194
rect 486 18130 550 18194
rect 567 18130 631 18194
rect 648 18130 712 18194
rect 729 18130 793 18194
rect 810 18130 874 18194
rect 891 18130 955 18194
rect 972 18130 1036 18194
rect 1053 18130 1117 18194
rect 1134 18130 1198 18194
rect 1215 18130 1279 18194
rect 1296 18130 1360 18194
rect 1377 18130 1441 18194
rect 1458 18130 1522 18194
rect 1539 18130 1603 18194
rect 1620 18130 1684 18194
rect 1701 18130 1765 18194
rect 1782 18130 1846 18194
rect 1863 18130 1927 18194
rect 1944 18130 2008 18194
rect 2025 18130 2089 18194
rect 2106 18130 2170 18194
rect 2187 18130 2251 18194
rect 2268 18130 2332 18194
rect 2349 18130 2413 18194
rect 2430 18130 2494 18194
rect 2511 18130 2575 18194
rect 2592 18130 2656 18194
rect 2673 18130 2737 18194
rect 2754 18130 2818 18194
rect 2835 18130 2899 18194
rect 2916 18130 2980 18194
rect 2997 18130 3061 18194
rect 3078 18130 3142 18194
rect 3159 18130 3223 18194
rect 3240 18130 3304 18194
rect 3321 18130 3385 18194
rect 3402 18130 3466 18194
rect 3483 18130 3547 18194
rect 3563 18130 3627 18194
rect 3643 18130 3707 18194
rect 3723 18130 3787 18194
rect 3803 18130 3867 18194
rect 3883 18130 3947 18194
rect 4016 18142 4080 18206
rect 4129 18142 4193 18206
rect 4242 18142 4306 18206
rect 4355 18142 4419 18206
rect 4478 18119 4542 18183
rect 4598 18119 4662 18183
rect 10350 18233 10414 18297
rect 10470 18233 10534 18297
rect 10593 18244 10657 18308
rect 10706 18244 10770 18308
rect 10819 18244 10883 18308
rect 10932 18244 10996 18308
rect 11065 18298 11129 18362
rect 11145 18298 11209 18362
rect 11225 18298 11289 18362
rect 11305 18298 11369 18362
rect 11385 18298 11449 18362
rect 11465 18298 11529 18362
rect 11546 18298 11610 18362
rect 11627 18298 11691 18362
rect 11708 18298 11772 18362
rect 11789 18298 11853 18362
rect 11870 18298 11934 18362
rect 11951 18298 12015 18362
rect 12032 18298 12096 18362
rect 12113 18298 12177 18362
rect 12194 18298 12258 18362
rect 12275 18298 12339 18362
rect 12356 18298 12420 18362
rect 12437 18298 12501 18362
rect 12518 18298 12582 18362
rect 12599 18298 12663 18362
rect 12680 18298 12744 18362
rect 12761 18298 12825 18362
rect 12842 18298 12906 18362
rect 12923 18298 12987 18362
rect 13004 18298 13068 18362
rect 13085 18298 13149 18362
rect 13166 18298 13230 18362
rect 13247 18298 13311 18362
rect 13328 18298 13392 18362
rect 13409 18298 13473 18362
rect 13490 18298 13554 18362
rect 13571 18298 13635 18362
rect 13652 18298 13716 18362
rect 13733 18298 13797 18362
rect 13814 18298 13878 18362
rect 13895 18298 13959 18362
rect 13976 18298 14040 18362
rect 14057 18298 14121 18362
rect 14138 18298 14202 18362
rect 14219 18298 14283 18362
rect 14300 18298 14364 18362
rect 14381 18298 14445 18362
rect 14462 18298 14526 18362
rect 14543 18298 14607 18362
rect 14624 18298 14688 18362
rect 14705 18298 14769 18362
rect 14786 18298 14850 18362
rect 11065 18214 11129 18278
rect 11145 18214 11209 18278
rect 11225 18214 11289 18278
rect 11305 18214 11369 18278
rect 11385 18214 11449 18278
rect 11465 18214 11529 18278
rect 11546 18214 11610 18278
rect 11627 18214 11691 18278
rect 11708 18214 11772 18278
rect 11789 18214 11853 18278
rect 11870 18214 11934 18278
rect 11951 18214 12015 18278
rect 12032 18214 12096 18278
rect 12113 18214 12177 18278
rect 12194 18214 12258 18278
rect 12275 18214 12339 18278
rect 12356 18214 12420 18278
rect 12437 18214 12501 18278
rect 12518 18214 12582 18278
rect 12599 18214 12663 18278
rect 12680 18214 12744 18278
rect 12761 18214 12825 18278
rect 12842 18214 12906 18278
rect 12923 18214 12987 18278
rect 13004 18214 13068 18278
rect 13085 18214 13149 18278
rect 13166 18214 13230 18278
rect 13247 18214 13311 18278
rect 13328 18214 13392 18278
rect 13409 18214 13473 18278
rect 13490 18214 13554 18278
rect 13571 18214 13635 18278
rect 13652 18214 13716 18278
rect 13733 18214 13797 18278
rect 13814 18214 13878 18278
rect 13895 18214 13959 18278
rect 13976 18214 14040 18278
rect 14057 18214 14121 18278
rect 14138 18214 14202 18278
rect 14219 18214 14283 18278
rect 14300 18214 14364 18278
rect 14381 18214 14445 18278
rect 14462 18214 14526 18278
rect 14543 18214 14607 18278
rect 14624 18214 14688 18278
rect 14705 18214 14769 18278
rect 14786 18214 14850 18278
rect 10350 18119 10414 18183
rect 10470 18119 10534 18183
rect 10593 18142 10657 18206
rect 10706 18142 10770 18206
rect 10819 18142 10883 18206
rect 10932 18142 10996 18206
rect 11065 18130 11129 18194
rect 11145 18130 11209 18194
rect 11225 18130 11289 18194
rect 11305 18130 11369 18194
rect 11385 18130 11449 18194
rect 11465 18130 11529 18194
rect 11546 18130 11610 18194
rect 11627 18130 11691 18194
rect 11708 18130 11772 18194
rect 11789 18130 11853 18194
rect 11870 18130 11934 18194
rect 11951 18130 12015 18194
rect 12032 18130 12096 18194
rect 12113 18130 12177 18194
rect 12194 18130 12258 18194
rect 12275 18130 12339 18194
rect 12356 18130 12420 18194
rect 12437 18130 12501 18194
rect 12518 18130 12582 18194
rect 12599 18130 12663 18194
rect 12680 18130 12744 18194
rect 12761 18130 12825 18194
rect 12842 18130 12906 18194
rect 12923 18130 12987 18194
rect 13004 18130 13068 18194
rect 13085 18130 13149 18194
rect 13166 18130 13230 18194
rect 13247 18130 13311 18194
rect 13328 18130 13392 18194
rect 13409 18130 13473 18194
rect 13490 18130 13554 18194
rect 13571 18130 13635 18194
rect 13652 18130 13716 18194
rect 13733 18130 13797 18194
rect 13814 18130 13878 18194
rect 13895 18130 13959 18194
rect 13976 18130 14040 18194
rect 14057 18130 14121 18194
rect 14138 18130 14202 18194
rect 14219 18130 14283 18194
rect 14300 18130 14364 18194
rect 14381 18130 14445 18194
rect 14462 18130 14526 18194
rect 14543 18130 14607 18194
rect 14624 18130 14688 18194
rect 14705 18130 14769 18194
rect 14786 18130 14850 18194
rect 137 14742 4841 18086
rect 137 14661 201 14725
rect 217 14661 281 14725
rect 297 14661 361 14725
rect 377 14661 441 14725
rect 457 14661 521 14725
rect 537 14661 601 14725
rect 617 14661 681 14725
rect 697 14661 761 14725
rect 777 14661 841 14725
rect 857 14661 921 14725
rect 937 14661 1001 14725
rect 1017 14661 1081 14725
rect 1097 14661 1161 14725
rect 1177 14661 1241 14725
rect 1257 14661 1321 14725
rect 1337 14661 1401 14725
rect 1417 14661 1481 14725
rect 1497 14661 1561 14725
rect 1577 14661 1641 14725
rect 1657 14661 1721 14725
rect 1737 14661 1801 14725
rect 1817 14661 1881 14725
rect 1897 14661 1961 14725
rect 1977 14661 2041 14725
rect 2057 14661 2121 14725
rect 2137 14661 2201 14725
rect 2217 14661 2281 14725
rect 2297 14661 2361 14725
rect 2377 14661 2441 14725
rect 2457 14661 2521 14725
rect 2537 14661 2601 14725
rect 2617 14661 2681 14725
rect 2697 14661 2761 14725
rect 2777 14661 2841 14725
rect 2857 14661 2921 14725
rect 2937 14661 3001 14725
rect 3017 14661 3081 14725
rect 3097 14661 3161 14725
rect 3177 14661 3241 14725
rect 3257 14661 3321 14725
rect 3337 14661 3401 14725
rect 3417 14661 3481 14725
rect 3497 14661 3561 14725
rect 3577 14661 3641 14725
rect 3657 14661 3721 14725
rect 3737 14661 3801 14725
rect 3817 14661 3881 14725
rect 3897 14661 3961 14725
rect 3977 14661 4041 14725
rect 4057 14661 4121 14725
rect 4137 14661 4201 14725
rect 4217 14661 4281 14725
rect 4297 14661 4361 14725
rect 4377 14661 4441 14725
rect 4457 14661 4521 14725
rect 4537 14661 4601 14725
rect 4617 14661 4681 14725
rect 4697 14661 4761 14725
rect 4777 14661 4841 14725
rect 137 14580 201 14644
rect 217 14580 281 14644
rect 297 14580 361 14644
rect 377 14580 441 14644
rect 457 14580 521 14644
rect 537 14580 601 14644
rect 617 14580 681 14644
rect 697 14580 761 14644
rect 777 14580 841 14644
rect 857 14580 921 14644
rect 937 14580 1001 14644
rect 1017 14580 1081 14644
rect 1097 14580 1161 14644
rect 1177 14580 1241 14644
rect 1257 14580 1321 14644
rect 1337 14580 1401 14644
rect 1417 14580 1481 14644
rect 1497 14580 1561 14644
rect 1577 14580 1641 14644
rect 1657 14580 1721 14644
rect 1737 14580 1801 14644
rect 1817 14580 1881 14644
rect 1897 14580 1961 14644
rect 1977 14580 2041 14644
rect 2057 14580 2121 14644
rect 2137 14580 2201 14644
rect 2217 14580 2281 14644
rect 2297 14580 2361 14644
rect 2377 14580 2441 14644
rect 2457 14580 2521 14644
rect 2537 14580 2601 14644
rect 2617 14580 2681 14644
rect 2697 14580 2761 14644
rect 2777 14580 2841 14644
rect 2857 14580 2921 14644
rect 2937 14580 3001 14644
rect 3017 14580 3081 14644
rect 3097 14580 3161 14644
rect 3177 14580 3241 14644
rect 3257 14580 3321 14644
rect 3337 14580 3401 14644
rect 3417 14580 3481 14644
rect 3497 14580 3561 14644
rect 3577 14580 3641 14644
rect 3657 14580 3721 14644
rect 3737 14580 3801 14644
rect 3817 14580 3881 14644
rect 3897 14580 3961 14644
rect 3977 14580 4041 14644
rect 4057 14580 4121 14644
rect 4137 14580 4201 14644
rect 4217 14580 4281 14644
rect 4297 14580 4361 14644
rect 4377 14580 4441 14644
rect 4457 14580 4521 14644
rect 4537 14580 4601 14644
rect 4617 14580 4681 14644
rect 4697 14580 4761 14644
rect 4777 14580 4841 14644
rect 137 14499 201 14563
rect 217 14499 281 14563
rect 297 14499 361 14563
rect 377 14499 441 14563
rect 457 14499 521 14563
rect 537 14499 601 14563
rect 617 14499 681 14563
rect 697 14499 761 14563
rect 777 14499 841 14563
rect 857 14499 921 14563
rect 937 14499 1001 14563
rect 1017 14499 1081 14563
rect 1097 14499 1161 14563
rect 1177 14499 1241 14563
rect 1257 14499 1321 14563
rect 1337 14499 1401 14563
rect 1417 14499 1481 14563
rect 1497 14499 1561 14563
rect 1577 14499 1641 14563
rect 1657 14499 1721 14563
rect 1737 14499 1801 14563
rect 1817 14499 1881 14563
rect 1897 14499 1961 14563
rect 1977 14499 2041 14563
rect 2057 14499 2121 14563
rect 2137 14499 2201 14563
rect 2217 14499 2281 14563
rect 2297 14499 2361 14563
rect 2377 14499 2441 14563
rect 2457 14499 2521 14563
rect 2537 14499 2601 14563
rect 2617 14499 2681 14563
rect 2697 14499 2761 14563
rect 2777 14499 2841 14563
rect 2857 14499 2921 14563
rect 2937 14499 3001 14563
rect 3017 14499 3081 14563
rect 3097 14499 3161 14563
rect 3177 14499 3241 14563
rect 3257 14499 3321 14563
rect 3337 14499 3401 14563
rect 3417 14499 3481 14563
rect 3497 14499 3561 14563
rect 3577 14499 3641 14563
rect 3657 14499 3721 14563
rect 3737 14499 3801 14563
rect 3817 14499 3881 14563
rect 3897 14499 3961 14563
rect 3977 14499 4041 14563
rect 4057 14499 4121 14563
rect 4137 14499 4201 14563
rect 4217 14499 4281 14563
rect 4297 14499 4361 14563
rect 4377 14499 4441 14563
rect 4457 14499 4521 14563
rect 4537 14499 4601 14563
rect 4617 14499 4681 14563
rect 4697 14499 4761 14563
rect 4777 14499 4841 14563
rect 137 14418 201 14482
rect 217 14418 281 14482
rect 297 14418 361 14482
rect 377 14418 441 14482
rect 457 14418 521 14482
rect 537 14418 601 14482
rect 617 14418 681 14482
rect 697 14418 761 14482
rect 777 14418 841 14482
rect 857 14418 921 14482
rect 937 14418 1001 14482
rect 1017 14418 1081 14482
rect 1097 14418 1161 14482
rect 1177 14418 1241 14482
rect 1257 14418 1321 14482
rect 1337 14418 1401 14482
rect 1417 14418 1481 14482
rect 1497 14418 1561 14482
rect 1577 14418 1641 14482
rect 1657 14418 1721 14482
rect 1737 14418 1801 14482
rect 1817 14418 1881 14482
rect 1897 14418 1961 14482
rect 1977 14418 2041 14482
rect 2057 14418 2121 14482
rect 2137 14418 2201 14482
rect 2217 14418 2281 14482
rect 2297 14418 2361 14482
rect 2377 14418 2441 14482
rect 2457 14418 2521 14482
rect 2537 14418 2601 14482
rect 2617 14418 2681 14482
rect 2697 14418 2761 14482
rect 2777 14418 2841 14482
rect 2857 14418 2921 14482
rect 2937 14418 3001 14482
rect 3017 14418 3081 14482
rect 3097 14418 3161 14482
rect 3177 14418 3241 14482
rect 3257 14418 3321 14482
rect 3337 14418 3401 14482
rect 3417 14418 3481 14482
rect 3497 14418 3561 14482
rect 3577 14418 3641 14482
rect 3657 14418 3721 14482
rect 3737 14418 3801 14482
rect 3817 14418 3881 14482
rect 3897 14418 3961 14482
rect 3977 14418 4041 14482
rect 4057 14418 4121 14482
rect 4137 14418 4201 14482
rect 4217 14418 4281 14482
rect 4297 14418 4361 14482
rect 4377 14418 4441 14482
rect 4457 14418 4521 14482
rect 4537 14418 4601 14482
rect 4617 14418 4681 14482
rect 4697 14418 4761 14482
rect 4777 14418 4841 14482
rect 137 14337 201 14401
rect 217 14337 281 14401
rect 297 14337 361 14401
rect 377 14337 441 14401
rect 457 14337 521 14401
rect 537 14337 601 14401
rect 617 14337 681 14401
rect 697 14337 761 14401
rect 777 14337 841 14401
rect 857 14337 921 14401
rect 937 14337 1001 14401
rect 1017 14337 1081 14401
rect 1097 14337 1161 14401
rect 1177 14337 1241 14401
rect 1257 14337 1321 14401
rect 1337 14337 1401 14401
rect 1417 14337 1481 14401
rect 1497 14337 1561 14401
rect 1577 14337 1641 14401
rect 1657 14337 1721 14401
rect 1737 14337 1801 14401
rect 1817 14337 1881 14401
rect 1897 14337 1961 14401
rect 1977 14337 2041 14401
rect 2057 14337 2121 14401
rect 2137 14337 2201 14401
rect 2217 14337 2281 14401
rect 2297 14337 2361 14401
rect 2377 14337 2441 14401
rect 2457 14337 2521 14401
rect 2537 14337 2601 14401
rect 2617 14337 2681 14401
rect 2697 14337 2761 14401
rect 2777 14337 2841 14401
rect 2857 14337 2921 14401
rect 2937 14337 3001 14401
rect 3017 14337 3081 14401
rect 3097 14337 3161 14401
rect 3177 14337 3241 14401
rect 3257 14337 3321 14401
rect 3337 14337 3401 14401
rect 3417 14337 3481 14401
rect 3497 14337 3561 14401
rect 3577 14337 3641 14401
rect 3657 14337 3721 14401
rect 3737 14337 3801 14401
rect 3817 14337 3881 14401
rect 3897 14337 3961 14401
rect 3977 14337 4041 14401
rect 4057 14337 4121 14401
rect 4137 14337 4201 14401
rect 4217 14337 4281 14401
rect 4297 14337 4361 14401
rect 4377 14337 4441 14401
rect 4457 14337 4521 14401
rect 4537 14337 4601 14401
rect 4617 14337 4681 14401
rect 4697 14337 4761 14401
rect 4777 14337 4841 14401
rect 137 14256 201 14320
rect 217 14256 281 14320
rect 297 14256 361 14320
rect 377 14256 441 14320
rect 457 14256 521 14320
rect 537 14256 601 14320
rect 617 14256 681 14320
rect 697 14256 761 14320
rect 777 14256 841 14320
rect 857 14256 921 14320
rect 937 14256 1001 14320
rect 1017 14256 1081 14320
rect 1097 14256 1161 14320
rect 1177 14256 1241 14320
rect 1257 14256 1321 14320
rect 1337 14256 1401 14320
rect 1417 14256 1481 14320
rect 1497 14256 1561 14320
rect 1577 14256 1641 14320
rect 1657 14256 1721 14320
rect 1737 14256 1801 14320
rect 1817 14256 1881 14320
rect 1897 14256 1961 14320
rect 1977 14256 2041 14320
rect 2057 14256 2121 14320
rect 2137 14256 2201 14320
rect 2217 14256 2281 14320
rect 2297 14256 2361 14320
rect 2377 14256 2441 14320
rect 2457 14256 2521 14320
rect 2537 14256 2601 14320
rect 2617 14256 2681 14320
rect 2697 14256 2761 14320
rect 2777 14256 2841 14320
rect 2857 14256 2921 14320
rect 2937 14256 3001 14320
rect 3017 14256 3081 14320
rect 3097 14256 3161 14320
rect 3177 14256 3241 14320
rect 3257 14256 3321 14320
rect 3337 14256 3401 14320
rect 3417 14256 3481 14320
rect 3497 14256 3561 14320
rect 3577 14256 3641 14320
rect 3657 14256 3721 14320
rect 3737 14256 3801 14320
rect 3817 14256 3881 14320
rect 3897 14256 3961 14320
rect 3977 14256 4041 14320
rect 4057 14256 4121 14320
rect 4137 14256 4201 14320
rect 4217 14256 4281 14320
rect 4297 14256 4361 14320
rect 4377 14256 4441 14320
rect 4457 14256 4521 14320
rect 4537 14256 4601 14320
rect 4617 14256 4681 14320
rect 4697 14256 4761 14320
rect 4777 14256 4841 14320
rect 137 14175 201 14239
rect 217 14175 281 14239
rect 297 14175 361 14239
rect 377 14175 441 14239
rect 457 14175 521 14239
rect 537 14175 601 14239
rect 617 14175 681 14239
rect 697 14175 761 14239
rect 777 14175 841 14239
rect 857 14175 921 14239
rect 937 14175 1001 14239
rect 1017 14175 1081 14239
rect 1097 14175 1161 14239
rect 1177 14175 1241 14239
rect 1257 14175 1321 14239
rect 1337 14175 1401 14239
rect 1417 14175 1481 14239
rect 1497 14175 1561 14239
rect 1577 14175 1641 14239
rect 1657 14175 1721 14239
rect 1737 14175 1801 14239
rect 1817 14175 1881 14239
rect 1897 14175 1961 14239
rect 1977 14175 2041 14239
rect 2057 14175 2121 14239
rect 2137 14175 2201 14239
rect 2217 14175 2281 14239
rect 2297 14175 2361 14239
rect 2377 14175 2441 14239
rect 2457 14175 2521 14239
rect 2537 14175 2601 14239
rect 2617 14175 2681 14239
rect 2697 14175 2761 14239
rect 2777 14175 2841 14239
rect 2857 14175 2921 14239
rect 2937 14175 3001 14239
rect 3017 14175 3081 14239
rect 3097 14175 3161 14239
rect 3177 14175 3241 14239
rect 3257 14175 3321 14239
rect 3337 14175 3401 14239
rect 3417 14175 3481 14239
rect 3497 14175 3561 14239
rect 3577 14175 3641 14239
rect 3657 14175 3721 14239
rect 3737 14175 3801 14239
rect 3817 14175 3881 14239
rect 3897 14175 3961 14239
rect 3977 14175 4041 14239
rect 4057 14175 4121 14239
rect 4137 14175 4201 14239
rect 4217 14175 4281 14239
rect 4297 14175 4361 14239
rect 4377 14175 4441 14239
rect 4457 14175 4521 14239
rect 4537 14175 4601 14239
rect 4617 14175 4681 14239
rect 4697 14175 4761 14239
rect 4777 14175 4841 14239
rect 137 14094 201 14158
rect 217 14094 281 14158
rect 297 14094 361 14158
rect 377 14094 441 14158
rect 457 14094 521 14158
rect 537 14094 601 14158
rect 617 14094 681 14158
rect 697 14094 761 14158
rect 777 14094 841 14158
rect 857 14094 921 14158
rect 937 14094 1001 14158
rect 1017 14094 1081 14158
rect 1097 14094 1161 14158
rect 1177 14094 1241 14158
rect 1257 14094 1321 14158
rect 1337 14094 1401 14158
rect 1417 14094 1481 14158
rect 1497 14094 1561 14158
rect 1577 14094 1641 14158
rect 1657 14094 1721 14158
rect 1737 14094 1801 14158
rect 1817 14094 1881 14158
rect 1897 14094 1961 14158
rect 1977 14094 2041 14158
rect 2057 14094 2121 14158
rect 2137 14094 2201 14158
rect 2217 14094 2281 14158
rect 2297 14094 2361 14158
rect 2377 14094 2441 14158
rect 2457 14094 2521 14158
rect 2537 14094 2601 14158
rect 2617 14094 2681 14158
rect 2697 14094 2761 14158
rect 2777 14094 2841 14158
rect 2857 14094 2921 14158
rect 2937 14094 3001 14158
rect 3017 14094 3081 14158
rect 3097 14094 3161 14158
rect 3177 14094 3241 14158
rect 3257 14094 3321 14158
rect 3337 14094 3401 14158
rect 3417 14094 3481 14158
rect 3497 14094 3561 14158
rect 3577 14094 3641 14158
rect 3657 14094 3721 14158
rect 3737 14094 3801 14158
rect 3817 14094 3881 14158
rect 3897 14094 3961 14158
rect 3977 14094 4041 14158
rect 4057 14094 4121 14158
rect 4137 14094 4201 14158
rect 4217 14094 4281 14158
rect 4297 14094 4361 14158
rect 4377 14094 4441 14158
rect 4457 14094 4521 14158
rect 4537 14094 4601 14158
rect 4617 14094 4681 14158
rect 4697 14094 4761 14158
rect 4777 14094 4841 14158
rect 137 14013 201 14077
rect 217 14013 281 14077
rect 297 14013 361 14077
rect 377 14013 441 14077
rect 457 14013 521 14077
rect 537 14013 601 14077
rect 617 14013 681 14077
rect 697 14013 761 14077
rect 777 14013 841 14077
rect 857 14013 921 14077
rect 937 14013 1001 14077
rect 1017 14013 1081 14077
rect 1097 14013 1161 14077
rect 1177 14013 1241 14077
rect 1257 14013 1321 14077
rect 1337 14013 1401 14077
rect 1417 14013 1481 14077
rect 1497 14013 1561 14077
rect 1577 14013 1641 14077
rect 1657 14013 1721 14077
rect 1737 14013 1801 14077
rect 1817 14013 1881 14077
rect 1897 14013 1961 14077
rect 1977 14013 2041 14077
rect 2057 14013 2121 14077
rect 2137 14013 2201 14077
rect 2217 14013 2281 14077
rect 2297 14013 2361 14077
rect 2377 14013 2441 14077
rect 2457 14013 2521 14077
rect 2537 14013 2601 14077
rect 2617 14013 2681 14077
rect 2697 14013 2761 14077
rect 2777 14013 2841 14077
rect 2857 14013 2921 14077
rect 2937 14013 3001 14077
rect 3017 14013 3081 14077
rect 3097 14013 3161 14077
rect 3177 14013 3241 14077
rect 3257 14013 3321 14077
rect 3337 14013 3401 14077
rect 3417 14013 3481 14077
rect 3497 14013 3561 14077
rect 3577 14013 3641 14077
rect 3657 14013 3721 14077
rect 3737 14013 3801 14077
rect 3817 14013 3881 14077
rect 3897 14013 3961 14077
rect 3977 14013 4041 14077
rect 4057 14013 4121 14077
rect 4137 14013 4201 14077
rect 4217 14013 4281 14077
rect 4297 14013 4361 14077
rect 4377 14013 4441 14077
rect 4457 14013 4521 14077
rect 4537 14013 4601 14077
rect 4617 14013 4681 14077
rect 4697 14013 4761 14077
rect 4777 14013 4841 14077
rect 10143 14742 14847 18086
rect 10143 14661 10207 14725
rect 10223 14661 10287 14725
rect 10303 14661 10367 14725
rect 10383 14661 10447 14725
rect 10463 14661 10527 14725
rect 10543 14661 10607 14725
rect 10623 14661 10687 14725
rect 10703 14661 10767 14725
rect 10783 14661 10847 14725
rect 10863 14661 10927 14725
rect 10943 14661 11007 14725
rect 11023 14661 11087 14725
rect 11103 14661 11167 14725
rect 11183 14661 11247 14725
rect 11263 14661 11327 14725
rect 11343 14661 11407 14725
rect 11423 14661 11487 14725
rect 11503 14661 11567 14725
rect 11583 14661 11647 14725
rect 11663 14661 11727 14725
rect 11743 14661 11807 14725
rect 11823 14661 11887 14725
rect 11903 14661 11967 14725
rect 11983 14661 12047 14725
rect 12063 14661 12127 14725
rect 12143 14661 12207 14725
rect 12223 14661 12287 14725
rect 12303 14661 12367 14725
rect 12383 14661 12447 14725
rect 12463 14661 12527 14725
rect 12543 14661 12607 14725
rect 12623 14661 12687 14725
rect 12703 14661 12767 14725
rect 12783 14661 12847 14725
rect 12863 14661 12927 14725
rect 12943 14661 13007 14725
rect 13023 14661 13087 14725
rect 13103 14661 13167 14725
rect 13183 14661 13247 14725
rect 13263 14661 13327 14725
rect 13343 14661 13407 14725
rect 13423 14661 13487 14725
rect 13503 14661 13567 14725
rect 13583 14661 13647 14725
rect 13663 14661 13727 14725
rect 13743 14661 13807 14725
rect 13823 14661 13887 14725
rect 13903 14661 13967 14725
rect 13983 14661 14047 14725
rect 14063 14661 14127 14725
rect 14143 14661 14207 14725
rect 14223 14661 14287 14725
rect 14303 14661 14367 14725
rect 14383 14661 14447 14725
rect 14463 14661 14527 14725
rect 14543 14661 14607 14725
rect 14623 14661 14687 14725
rect 14703 14661 14767 14725
rect 14783 14661 14847 14725
rect 10143 14580 10207 14644
rect 10223 14580 10287 14644
rect 10303 14580 10367 14644
rect 10383 14580 10447 14644
rect 10463 14580 10527 14644
rect 10543 14580 10607 14644
rect 10623 14580 10687 14644
rect 10703 14580 10767 14644
rect 10783 14580 10847 14644
rect 10863 14580 10927 14644
rect 10943 14580 11007 14644
rect 11023 14580 11087 14644
rect 11103 14580 11167 14644
rect 11183 14580 11247 14644
rect 11263 14580 11327 14644
rect 11343 14580 11407 14644
rect 11423 14580 11487 14644
rect 11503 14580 11567 14644
rect 11583 14580 11647 14644
rect 11663 14580 11727 14644
rect 11743 14580 11807 14644
rect 11823 14580 11887 14644
rect 11903 14580 11967 14644
rect 11983 14580 12047 14644
rect 12063 14580 12127 14644
rect 12143 14580 12207 14644
rect 12223 14580 12287 14644
rect 12303 14580 12367 14644
rect 12383 14580 12447 14644
rect 12463 14580 12527 14644
rect 12543 14580 12607 14644
rect 12623 14580 12687 14644
rect 12703 14580 12767 14644
rect 12783 14580 12847 14644
rect 12863 14580 12927 14644
rect 12943 14580 13007 14644
rect 13023 14580 13087 14644
rect 13103 14580 13167 14644
rect 13183 14580 13247 14644
rect 13263 14580 13327 14644
rect 13343 14580 13407 14644
rect 13423 14580 13487 14644
rect 13503 14580 13567 14644
rect 13583 14580 13647 14644
rect 13663 14580 13727 14644
rect 13743 14580 13807 14644
rect 13823 14580 13887 14644
rect 13903 14580 13967 14644
rect 13983 14580 14047 14644
rect 14063 14580 14127 14644
rect 14143 14580 14207 14644
rect 14223 14580 14287 14644
rect 14303 14580 14367 14644
rect 14383 14580 14447 14644
rect 14463 14580 14527 14644
rect 14543 14580 14607 14644
rect 14623 14580 14687 14644
rect 14703 14580 14767 14644
rect 14783 14580 14847 14644
rect 10143 14499 10207 14563
rect 10223 14499 10287 14563
rect 10303 14499 10367 14563
rect 10383 14499 10447 14563
rect 10463 14499 10527 14563
rect 10543 14499 10607 14563
rect 10623 14499 10687 14563
rect 10703 14499 10767 14563
rect 10783 14499 10847 14563
rect 10863 14499 10927 14563
rect 10943 14499 11007 14563
rect 11023 14499 11087 14563
rect 11103 14499 11167 14563
rect 11183 14499 11247 14563
rect 11263 14499 11327 14563
rect 11343 14499 11407 14563
rect 11423 14499 11487 14563
rect 11503 14499 11567 14563
rect 11583 14499 11647 14563
rect 11663 14499 11727 14563
rect 11743 14499 11807 14563
rect 11823 14499 11887 14563
rect 11903 14499 11967 14563
rect 11983 14499 12047 14563
rect 12063 14499 12127 14563
rect 12143 14499 12207 14563
rect 12223 14499 12287 14563
rect 12303 14499 12367 14563
rect 12383 14499 12447 14563
rect 12463 14499 12527 14563
rect 12543 14499 12607 14563
rect 12623 14499 12687 14563
rect 12703 14499 12767 14563
rect 12783 14499 12847 14563
rect 12863 14499 12927 14563
rect 12943 14499 13007 14563
rect 13023 14499 13087 14563
rect 13103 14499 13167 14563
rect 13183 14499 13247 14563
rect 13263 14499 13327 14563
rect 13343 14499 13407 14563
rect 13423 14499 13487 14563
rect 13503 14499 13567 14563
rect 13583 14499 13647 14563
rect 13663 14499 13727 14563
rect 13743 14499 13807 14563
rect 13823 14499 13887 14563
rect 13903 14499 13967 14563
rect 13983 14499 14047 14563
rect 14063 14499 14127 14563
rect 14143 14499 14207 14563
rect 14223 14499 14287 14563
rect 14303 14499 14367 14563
rect 14383 14499 14447 14563
rect 14463 14499 14527 14563
rect 14543 14499 14607 14563
rect 14623 14499 14687 14563
rect 14703 14499 14767 14563
rect 14783 14499 14847 14563
rect 10143 14418 10207 14482
rect 10223 14418 10287 14482
rect 10303 14418 10367 14482
rect 10383 14418 10447 14482
rect 10463 14418 10527 14482
rect 10543 14418 10607 14482
rect 10623 14418 10687 14482
rect 10703 14418 10767 14482
rect 10783 14418 10847 14482
rect 10863 14418 10927 14482
rect 10943 14418 11007 14482
rect 11023 14418 11087 14482
rect 11103 14418 11167 14482
rect 11183 14418 11247 14482
rect 11263 14418 11327 14482
rect 11343 14418 11407 14482
rect 11423 14418 11487 14482
rect 11503 14418 11567 14482
rect 11583 14418 11647 14482
rect 11663 14418 11727 14482
rect 11743 14418 11807 14482
rect 11823 14418 11887 14482
rect 11903 14418 11967 14482
rect 11983 14418 12047 14482
rect 12063 14418 12127 14482
rect 12143 14418 12207 14482
rect 12223 14418 12287 14482
rect 12303 14418 12367 14482
rect 12383 14418 12447 14482
rect 12463 14418 12527 14482
rect 12543 14418 12607 14482
rect 12623 14418 12687 14482
rect 12703 14418 12767 14482
rect 12783 14418 12847 14482
rect 12863 14418 12927 14482
rect 12943 14418 13007 14482
rect 13023 14418 13087 14482
rect 13103 14418 13167 14482
rect 13183 14418 13247 14482
rect 13263 14418 13327 14482
rect 13343 14418 13407 14482
rect 13423 14418 13487 14482
rect 13503 14418 13567 14482
rect 13583 14418 13647 14482
rect 13663 14418 13727 14482
rect 13743 14418 13807 14482
rect 13823 14418 13887 14482
rect 13903 14418 13967 14482
rect 13983 14418 14047 14482
rect 14063 14418 14127 14482
rect 14143 14418 14207 14482
rect 14223 14418 14287 14482
rect 14303 14418 14367 14482
rect 14383 14418 14447 14482
rect 14463 14418 14527 14482
rect 14543 14418 14607 14482
rect 14623 14418 14687 14482
rect 14703 14418 14767 14482
rect 14783 14418 14847 14482
rect 10143 14337 10207 14401
rect 10223 14337 10287 14401
rect 10303 14337 10367 14401
rect 10383 14337 10447 14401
rect 10463 14337 10527 14401
rect 10543 14337 10607 14401
rect 10623 14337 10687 14401
rect 10703 14337 10767 14401
rect 10783 14337 10847 14401
rect 10863 14337 10927 14401
rect 10943 14337 11007 14401
rect 11023 14337 11087 14401
rect 11103 14337 11167 14401
rect 11183 14337 11247 14401
rect 11263 14337 11327 14401
rect 11343 14337 11407 14401
rect 11423 14337 11487 14401
rect 11503 14337 11567 14401
rect 11583 14337 11647 14401
rect 11663 14337 11727 14401
rect 11743 14337 11807 14401
rect 11823 14337 11887 14401
rect 11903 14337 11967 14401
rect 11983 14337 12047 14401
rect 12063 14337 12127 14401
rect 12143 14337 12207 14401
rect 12223 14337 12287 14401
rect 12303 14337 12367 14401
rect 12383 14337 12447 14401
rect 12463 14337 12527 14401
rect 12543 14337 12607 14401
rect 12623 14337 12687 14401
rect 12703 14337 12767 14401
rect 12783 14337 12847 14401
rect 12863 14337 12927 14401
rect 12943 14337 13007 14401
rect 13023 14337 13087 14401
rect 13103 14337 13167 14401
rect 13183 14337 13247 14401
rect 13263 14337 13327 14401
rect 13343 14337 13407 14401
rect 13423 14337 13487 14401
rect 13503 14337 13567 14401
rect 13583 14337 13647 14401
rect 13663 14337 13727 14401
rect 13743 14337 13807 14401
rect 13823 14337 13887 14401
rect 13903 14337 13967 14401
rect 13983 14337 14047 14401
rect 14063 14337 14127 14401
rect 14143 14337 14207 14401
rect 14223 14337 14287 14401
rect 14303 14337 14367 14401
rect 14383 14337 14447 14401
rect 14463 14337 14527 14401
rect 14543 14337 14607 14401
rect 14623 14337 14687 14401
rect 14703 14337 14767 14401
rect 14783 14337 14847 14401
rect 10143 14256 10207 14320
rect 10223 14256 10287 14320
rect 10303 14256 10367 14320
rect 10383 14256 10447 14320
rect 10463 14256 10527 14320
rect 10543 14256 10607 14320
rect 10623 14256 10687 14320
rect 10703 14256 10767 14320
rect 10783 14256 10847 14320
rect 10863 14256 10927 14320
rect 10943 14256 11007 14320
rect 11023 14256 11087 14320
rect 11103 14256 11167 14320
rect 11183 14256 11247 14320
rect 11263 14256 11327 14320
rect 11343 14256 11407 14320
rect 11423 14256 11487 14320
rect 11503 14256 11567 14320
rect 11583 14256 11647 14320
rect 11663 14256 11727 14320
rect 11743 14256 11807 14320
rect 11823 14256 11887 14320
rect 11903 14256 11967 14320
rect 11983 14256 12047 14320
rect 12063 14256 12127 14320
rect 12143 14256 12207 14320
rect 12223 14256 12287 14320
rect 12303 14256 12367 14320
rect 12383 14256 12447 14320
rect 12463 14256 12527 14320
rect 12543 14256 12607 14320
rect 12623 14256 12687 14320
rect 12703 14256 12767 14320
rect 12783 14256 12847 14320
rect 12863 14256 12927 14320
rect 12943 14256 13007 14320
rect 13023 14256 13087 14320
rect 13103 14256 13167 14320
rect 13183 14256 13247 14320
rect 13263 14256 13327 14320
rect 13343 14256 13407 14320
rect 13423 14256 13487 14320
rect 13503 14256 13567 14320
rect 13583 14256 13647 14320
rect 13663 14256 13727 14320
rect 13743 14256 13807 14320
rect 13823 14256 13887 14320
rect 13903 14256 13967 14320
rect 13983 14256 14047 14320
rect 14063 14256 14127 14320
rect 14143 14256 14207 14320
rect 14223 14256 14287 14320
rect 14303 14256 14367 14320
rect 14383 14256 14447 14320
rect 14463 14256 14527 14320
rect 14543 14256 14607 14320
rect 14623 14256 14687 14320
rect 14703 14256 14767 14320
rect 14783 14256 14847 14320
rect 10143 14175 10207 14239
rect 10223 14175 10287 14239
rect 10303 14175 10367 14239
rect 10383 14175 10447 14239
rect 10463 14175 10527 14239
rect 10543 14175 10607 14239
rect 10623 14175 10687 14239
rect 10703 14175 10767 14239
rect 10783 14175 10847 14239
rect 10863 14175 10927 14239
rect 10943 14175 11007 14239
rect 11023 14175 11087 14239
rect 11103 14175 11167 14239
rect 11183 14175 11247 14239
rect 11263 14175 11327 14239
rect 11343 14175 11407 14239
rect 11423 14175 11487 14239
rect 11503 14175 11567 14239
rect 11583 14175 11647 14239
rect 11663 14175 11727 14239
rect 11743 14175 11807 14239
rect 11823 14175 11887 14239
rect 11903 14175 11967 14239
rect 11983 14175 12047 14239
rect 12063 14175 12127 14239
rect 12143 14175 12207 14239
rect 12223 14175 12287 14239
rect 12303 14175 12367 14239
rect 12383 14175 12447 14239
rect 12463 14175 12527 14239
rect 12543 14175 12607 14239
rect 12623 14175 12687 14239
rect 12703 14175 12767 14239
rect 12783 14175 12847 14239
rect 12863 14175 12927 14239
rect 12943 14175 13007 14239
rect 13023 14175 13087 14239
rect 13103 14175 13167 14239
rect 13183 14175 13247 14239
rect 13263 14175 13327 14239
rect 13343 14175 13407 14239
rect 13423 14175 13487 14239
rect 13503 14175 13567 14239
rect 13583 14175 13647 14239
rect 13663 14175 13727 14239
rect 13743 14175 13807 14239
rect 13823 14175 13887 14239
rect 13903 14175 13967 14239
rect 13983 14175 14047 14239
rect 14063 14175 14127 14239
rect 14143 14175 14207 14239
rect 14223 14175 14287 14239
rect 14303 14175 14367 14239
rect 14383 14175 14447 14239
rect 14463 14175 14527 14239
rect 14543 14175 14607 14239
rect 14623 14175 14687 14239
rect 14703 14175 14767 14239
rect 14783 14175 14847 14239
rect 10143 14094 10207 14158
rect 10223 14094 10287 14158
rect 10303 14094 10367 14158
rect 10383 14094 10447 14158
rect 10463 14094 10527 14158
rect 10543 14094 10607 14158
rect 10623 14094 10687 14158
rect 10703 14094 10767 14158
rect 10783 14094 10847 14158
rect 10863 14094 10927 14158
rect 10943 14094 11007 14158
rect 11023 14094 11087 14158
rect 11103 14094 11167 14158
rect 11183 14094 11247 14158
rect 11263 14094 11327 14158
rect 11343 14094 11407 14158
rect 11423 14094 11487 14158
rect 11503 14094 11567 14158
rect 11583 14094 11647 14158
rect 11663 14094 11727 14158
rect 11743 14094 11807 14158
rect 11823 14094 11887 14158
rect 11903 14094 11967 14158
rect 11983 14094 12047 14158
rect 12063 14094 12127 14158
rect 12143 14094 12207 14158
rect 12223 14094 12287 14158
rect 12303 14094 12367 14158
rect 12383 14094 12447 14158
rect 12463 14094 12527 14158
rect 12543 14094 12607 14158
rect 12623 14094 12687 14158
rect 12703 14094 12767 14158
rect 12783 14094 12847 14158
rect 12863 14094 12927 14158
rect 12943 14094 13007 14158
rect 13023 14094 13087 14158
rect 13103 14094 13167 14158
rect 13183 14094 13247 14158
rect 13263 14094 13327 14158
rect 13343 14094 13407 14158
rect 13423 14094 13487 14158
rect 13503 14094 13567 14158
rect 13583 14094 13647 14158
rect 13663 14094 13727 14158
rect 13743 14094 13807 14158
rect 13823 14094 13887 14158
rect 13903 14094 13967 14158
rect 13983 14094 14047 14158
rect 14063 14094 14127 14158
rect 14143 14094 14207 14158
rect 14223 14094 14287 14158
rect 14303 14094 14367 14158
rect 14383 14094 14447 14158
rect 14463 14094 14527 14158
rect 14543 14094 14607 14158
rect 14623 14094 14687 14158
rect 14703 14094 14767 14158
rect 14783 14094 14847 14158
rect 10143 14013 10207 14077
rect 10223 14013 10287 14077
rect 10303 14013 10367 14077
rect 10383 14013 10447 14077
rect 10463 14013 10527 14077
rect 10543 14013 10607 14077
rect 10623 14013 10687 14077
rect 10703 14013 10767 14077
rect 10783 14013 10847 14077
rect 10863 14013 10927 14077
rect 10943 14013 11007 14077
rect 11023 14013 11087 14077
rect 11103 14013 11167 14077
rect 11183 14013 11247 14077
rect 11263 14013 11327 14077
rect 11343 14013 11407 14077
rect 11423 14013 11487 14077
rect 11503 14013 11567 14077
rect 11583 14013 11647 14077
rect 11663 14013 11727 14077
rect 11743 14013 11807 14077
rect 11823 14013 11887 14077
rect 11903 14013 11967 14077
rect 11983 14013 12047 14077
rect 12063 14013 12127 14077
rect 12143 14013 12207 14077
rect 12223 14013 12287 14077
rect 12303 14013 12367 14077
rect 12383 14013 12447 14077
rect 12463 14013 12527 14077
rect 12543 14013 12607 14077
rect 12623 14013 12687 14077
rect 12703 14013 12767 14077
rect 12783 14013 12847 14077
rect 12863 14013 12927 14077
rect 12943 14013 13007 14077
rect 13023 14013 13087 14077
rect 13103 14013 13167 14077
rect 13183 14013 13247 14077
rect 13263 14013 13327 14077
rect 13343 14013 13407 14077
rect 13423 14013 13487 14077
rect 13503 14013 13567 14077
rect 13583 14013 13647 14077
rect 13663 14013 13727 14077
rect 13743 14013 13807 14077
rect 13823 14013 13887 14077
rect 13903 14013 13967 14077
rect 13983 14013 14047 14077
rect 14063 14013 14127 14077
rect 14143 14013 14207 14077
rect 14223 14013 14287 14077
rect 14303 14013 14367 14077
rect 14383 14013 14447 14077
rect 14463 14013 14527 14077
rect 14543 14013 14607 14077
rect 14623 14013 14687 14077
rect 14703 14013 14767 14077
rect 14783 14013 14847 14077
rect 105 13640 169 13704
rect 186 13640 250 13704
rect 267 13640 331 13704
rect 348 13640 412 13704
rect 429 13640 493 13704
rect 510 13640 574 13704
rect 591 13640 655 13704
rect 672 13640 736 13704
rect 753 13640 817 13704
rect 834 13640 898 13704
rect 915 13640 979 13704
rect 996 13640 1060 13704
rect 1077 13640 1141 13704
rect 1158 13640 1222 13704
rect 1239 13640 1303 13704
rect 1320 13640 1384 13704
rect 1401 13640 1465 13704
rect 1482 13640 1546 13704
rect 1563 13640 1627 13704
rect 1644 13640 1708 13704
rect 1725 13640 1789 13704
rect 1806 13640 1870 13704
rect 1887 13640 1951 13704
rect 1968 13640 2032 13704
rect 2049 13640 2113 13704
rect 2130 13640 2194 13704
rect 2211 13640 2275 13704
rect 2292 13640 2356 13704
rect 2373 13640 2437 13704
rect 2454 13640 2518 13704
rect 2535 13640 2599 13704
rect 2616 13640 2680 13704
rect 2697 13640 2761 13704
rect 2778 13640 2842 13704
rect 2859 13640 2923 13704
rect 2940 13640 3004 13704
rect 3021 13640 3085 13704
rect 3102 13640 3166 13704
rect 3183 13640 3247 13704
rect 3264 13640 3328 13704
rect 3345 13640 3409 13704
rect 3426 13640 3490 13704
rect 3507 13640 3571 13704
rect 3588 13640 3652 13704
rect 3669 13640 3733 13704
rect 3750 13640 3814 13704
rect 3831 13640 3895 13704
rect 3912 13640 3976 13704
rect 3993 13640 4057 13704
rect 4074 13640 4138 13704
rect 4155 13640 4219 13704
rect 4236 13640 4300 13704
rect 4317 13640 4381 13704
rect 4399 13640 4463 13704
rect 4481 13640 4545 13704
rect 4563 13640 4627 13704
rect 4645 13640 4709 13704
rect 4727 13640 4791 13704
rect 4809 13640 4873 13704
rect 105 13558 169 13622
rect 186 13558 250 13622
rect 267 13558 331 13622
rect 348 13558 412 13622
rect 429 13558 493 13622
rect 510 13558 574 13622
rect 591 13558 655 13622
rect 672 13558 736 13622
rect 753 13558 817 13622
rect 834 13558 898 13622
rect 915 13558 979 13622
rect 996 13558 1060 13622
rect 1077 13558 1141 13622
rect 1158 13558 1222 13622
rect 1239 13558 1303 13622
rect 1320 13558 1384 13622
rect 1401 13558 1465 13622
rect 1482 13558 1546 13622
rect 1563 13558 1627 13622
rect 1644 13558 1708 13622
rect 1725 13558 1789 13622
rect 1806 13558 1870 13622
rect 1887 13558 1951 13622
rect 1968 13558 2032 13622
rect 2049 13558 2113 13622
rect 2130 13558 2194 13622
rect 2211 13558 2275 13622
rect 2292 13558 2356 13622
rect 2373 13558 2437 13622
rect 2454 13558 2518 13622
rect 2535 13558 2599 13622
rect 2616 13558 2680 13622
rect 2697 13558 2761 13622
rect 2778 13558 2842 13622
rect 2859 13558 2923 13622
rect 2940 13558 3004 13622
rect 3021 13558 3085 13622
rect 3102 13558 3166 13622
rect 3183 13558 3247 13622
rect 3264 13558 3328 13622
rect 3345 13558 3409 13622
rect 3426 13558 3490 13622
rect 3507 13558 3571 13622
rect 3588 13558 3652 13622
rect 3669 13558 3733 13622
rect 3750 13558 3814 13622
rect 3831 13558 3895 13622
rect 3912 13558 3976 13622
rect 3993 13558 4057 13622
rect 4074 13558 4138 13622
rect 4155 13558 4219 13622
rect 4236 13558 4300 13622
rect 4317 13558 4381 13622
rect 4399 13558 4463 13622
rect 4481 13558 4545 13622
rect 4563 13558 4627 13622
rect 4645 13558 4709 13622
rect 4727 13558 4791 13622
rect 4809 13558 4873 13622
rect 105 13476 169 13540
rect 186 13476 250 13540
rect 267 13476 331 13540
rect 348 13476 412 13540
rect 429 13476 493 13540
rect 510 13476 574 13540
rect 591 13476 655 13540
rect 672 13476 736 13540
rect 753 13476 817 13540
rect 834 13476 898 13540
rect 915 13476 979 13540
rect 996 13476 1060 13540
rect 1077 13476 1141 13540
rect 1158 13476 1222 13540
rect 1239 13476 1303 13540
rect 1320 13476 1384 13540
rect 1401 13476 1465 13540
rect 1482 13476 1546 13540
rect 1563 13476 1627 13540
rect 1644 13476 1708 13540
rect 1725 13476 1789 13540
rect 1806 13476 1870 13540
rect 1887 13476 1951 13540
rect 1968 13476 2032 13540
rect 2049 13476 2113 13540
rect 2130 13476 2194 13540
rect 2211 13476 2275 13540
rect 2292 13476 2356 13540
rect 2373 13476 2437 13540
rect 2454 13476 2518 13540
rect 2535 13476 2599 13540
rect 2616 13476 2680 13540
rect 2697 13476 2761 13540
rect 2778 13476 2842 13540
rect 2859 13476 2923 13540
rect 2940 13476 3004 13540
rect 3021 13476 3085 13540
rect 3102 13476 3166 13540
rect 3183 13476 3247 13540
rect 3264 13476 3328 13540
rect 3345 13476 3409 13540
rect 3426 13476 3490 13540
rect 3507 13476 3571 13540
rect 3588 13476 3652 13540
rect 3669 13476 3733 13540
rect 3750 13476 3814 13540
rect 3831 13476 3895 13540
rect 3912 13476 3976 13540
rect 3993 13476 4057 13540
rect 4074 13476 4138 13540
rect 4155 13476 4219 13540
rect 4236 13476 4300 13540
rect 4317 13476 4381 13540
rect 4399 13476 4463 13540
rect 4481 13476 4545 13540
rect 4563 13476 4627 13540
rect 4645 13476 4709 13540
rect 4727 13476 4791 13540
rect 4809 13476 4873 13540
rect 105 13394 169 13458
rect 186 13394 250 13458
rect 267 13394 331 13458
rect 348 13394 412 13458
rect 429 13394 493 13458
rect 510 13394 574 13458
rect 591 13394 655 13458
rect 672 13394 736 13458
rect 753 13394 817 13458
rect 834 13394 898 13458
rect 915 13394 979 13458
rect 996 13394 1060 13458
rect 1077 13394 1141 13458
rect 1158 13394 1222 13458
rect 1239 13394 1303 13458
rect 1320 13394 1384 13458
rect 1401 13394 1465 13458
rect 1482 13394 1546 13458
rect 1563 13394 1627 13458
rect 1644 13394 1708 13458
rect 1725 13394 1789 13458
rect 1806 13394 1870 13458
rect 1887 13394 1951 13458
rect 1968 13394 2032 13458
rect 2049 13394 2113 13458
rect 2130 13394 2194 13458
rect 2211 13394 2275 13458
rect 2292 13394 2356 13458
rect 2373 13394 2437 13458
rect 2454 13394 2518 13458
rect 2535 13394 2599 13458
rect 2616 13394 2680 13458
rect 2697 13394 2761 13458
rect 2778 13394 2842 13458
rect 2859 13394 2923 13458
rect 2940 13394 3004 13458
rect 3021 13394 3085 13458
rect 3102 13394 3166 13458
rect 3183 13394 3247 13458
rect 3264 13394 3328 13458
rect 3345 13394 3409 13458
rect 3426 13394 3490 13458
rect 3507 13394 3571 13458
rect 3588 13394 3652 13458
rect 3669 13394 3733 13458
rect 3750 13394 3814 13458
rect 3831 13394 3895 13458
rect 3912 13394 3976 13458
rect 3993 13394 4057 13458
rect 4074 13394 4138 13458
rect 4155 13394 4219 13458
rect 4236 13394 4300 13458
rect 4317 13394 4381 13458
rect 4399 13394 4463 13458
rect 4481 13394 4545 13458
rect 4563 13394 4627 13458
rect 4645 13394 4709 13458
rect 4727 13394 4791 13458
rect 4809 13394 4873 13458
rect 105 13312 169 13376
rect 186 13312 250 13376
rect 267 13312 331 13376
rect 348 13312 412 13376
rect 429 13312 493 13376
rect 510 13312 574 13376
rect 591 13312 655 13376
rect 672 13312 736 13376
rect 753 13312 817 13376
rect 834 13312 898 13376
rect 915 13312 979 13376
rect 996 13312 1060 13376
rect 1077 13312 1141 13376
rect 1158 13312 1222 13376
rect 1239 13312 1303 13376
rect 1320 13312 1384 13376
rect 1401 13312 1465 13376
rect 1482 13312 1546 13376
rect 1563 13312 1627 13376
rect 1644 13312 1708 13376
rect 1725 13312 1789 13376
rect 1806 13312 1870 13376
rect 1887 13312 1951 13376
rect 1968 13312 2032 13376
rect 2049 13312 2113 13376
rect 2130 13312 2194 13376
rect 2211 13312 2275 13376
rect 2292 13312 2356 13376
rect 2373 13312 2437 13376
rect 2454 13312 2518 13376
rect 2535 13312 2599 13376
rect 2616 13312 2680 13376
rect 2697 13312 2761 13376
rect 2778 13312 2842 13376
rect 2859 13312 2923 13376
rect 2940 13312 3004 13376
rect 3021 13312 3085 13376
rect 3102 13312 3166 13376
rect 3183 13312 3247 13376
rect 3264 13312 3328 13376
rect 3345 13312 3409 13376
rect 3426 13312 3490 13376
rect 3507 13312 3571 13376
rect 3588 13312 3652 13376
rect 3669 13312 3733 13376
rect 3750 13312 3814 13376
rect 3831 13312 3895 13376
rect 3912 13312 3976 13376
rect 3993 13312 4057 13376
rect 4074 13312 4138 13376
rect 4155 13312 4219 13376
rect 4236 13312 4300 13376
rect 4317 13312 4381 13376
rect 4399 13312 4463 13376
rect 4481 13312 4545 13376
rect 4563 13312 4627 13376
rect 4645 13312 4709 13376
rect 4727 13312 4791 13376
rect 4809 13312 4873 13376
rect 105 13230 169 13294
rect 186 13230 250 13294
rect 267 13230 331 13294
rect 348 13230 412 13294
rect 429 13230 493 13294
rect 510 13230 574 13294
rect 591 13230 655 13294
rect 672 13230 736 13294
rect 753 13230 817 13294
rect 834 13230 898 13294
rect 915 13230 979 13294
rect 996 13230 1060 13294
rect 1077 13230 1141 13294
rect 1158 13230 1222 13294
rect 1239 13230 1303 13294
rect 1320 13230 1384 13294
rect 1401 13230 1465 13294
rect 1482 13230 1546 13294
rect 1563 13230 1627 13294
rect 1644 13230 1708 13294
rect 1725 13230 1789 13294
rect 1806 13230 1870 13294
rect 1887 13230 1951 13294
rect 1968 13230 2032 13294
rect 2049 13230 2113 13294
rect 2130 13230 2194 13294
rect 2211 13230 2275 13294
rect 2292 13230 2356 13294
rect 2373 13230 2437 13294
rect 2454 13230 2518 13294
rect 2535 13230 2599 13294
rect 2616 13230 2680 13294
rect 2697 13230 2761 13294
rect 2778 13230 2842 13294
rect 2859 13230 2923 13294
rect 2940 13230 3004 13294
rect 3021 13230 3085 13294
rect 3102 13230 3166 13294
rect 3183 13230 3247 13294
rect 3264 13230 3328 13294
rect 3345 13230 3409 13294
rect 3426 13230 3490 13294
rect 3507 13230 3571 13294
rect 3588 13230 3652 13294
rect 3669 13230 3733 13294
rect 3750 13230 3814 13294
rect 3831 13230 3895 13294
rect 3912 13230 3976 13294
rect 3993 13230 4057 13294
rect 4074 13230 4138 13294
rect 4155 13230 4219 13294
rect 4236 13230 4300 13294
rect 4317 13230 4381 13294
rect 4399 13230 4463 13294
rect 4481 13230 4545 13294
rect 4563 13230 4627 13294
rect 4645 13230 4709 13294
rect 4727 13230 4791 13294
rect 4809 13230 4873 13294
rect 105 13148 169 13212
rect 186 13148 250 13212
rect 267 13148 331 13212
rect 348 13148 412 13212
rect 429 13148 493 13212
rect 510 13148 574 13212
rect 591 13148 655 13212
rect 672 13148 736 13212
rect 753 13148 817 13212
rect 834 13148 898 13212
rect 915 13148 979 13212
rect 996 13148 1060 13212
rect 1077 13148 1141 13212
rect 1158 13148 1222 13212
rect 1239 13148 1303 13212
rect 1320 13148 1384 13212
rect 1401 13148 1465 13212
rect 1482 13148 1546 13212
rect 1563 13148 1627 13212
rect 1644 13148 1708 13212
rect 1725 13148 1789 13212
rect 1806 13148 1870 13212
rect 1887 13148 1951 13212
rect 1968 13148 2032 13212
rect 2049 13148 2113 13212
rect 2130 13148 2194 13212
rect 2211 13148 2275 13212
rect 2292 13148 2356 13212
rect 2373 13148 2437 13212
rect 2454 13148 2518 13212
rect 2535 13148 2599 13212
rect 2616 13148 2680 13212
rect 2697 13148 2761 13212
rect 2778 13148 2842 13212
rect 2859 13148 2923 13212
rect 2940 13148 3004 13212
rect 3021 13148 3085 13212
rect 3102 13148 3166 13212
rect 3183 13148 3247 13212
rect 3264 13148 3328 13212
rect 3345 13148 3409 13212
rect 3426 13148 3490 13212
rect 3507 13148 3571 13212
rect 3588 13148 3652 13212
rect 3669 13148 3733 13212
rect 3750 13148 3814 13212
rect 3831 13148 3895 13212
rect 3912 13148 3976 13212
rect 3993 13148 4057 13212
rect 4074 13148 4138 13212
rect 4155 13148 4219 13212
rect 4236 13148 4300 13212
rect 4317 13148 4381 13212
rect 4399 13148 4463 13212
rect 4481 13148 4545 13212
rect 4563 13148 4627 13212
rect 4645 13148 4709 13212
rect 4727 13148 4791 13212
rect 4809 13148 4873 13212
rect 105 13066 169 13130
rect 186 13066 250 13130
rect 267 13066 331 13130
rect 348 13066 412 13130
rect 429 13066 493 13130
rect 510 13066 574 13130
rect 591 13066 655 13130
rect 672 13066 736 13130
rect 753 13066 817 13130
rect 834 13066 898 13130
rect 915 13066 979 13130
rect 996 13066 1060 13130
rect 1077 13066 1141 13130
rect 1158 13066 1222 13130
rect 1239 13066 1303 13130
rect 1320 13066 1384 13130
rect 1401 13066 1465 13130
rect 1482 13066 1546 13130
rect 1563 13066 1627 13130
rect 1644 13066 1708 13130
rect 1725 13066 1789 13130
rect 1806 13066 1870 13130
rect 1887 13066 1951 13130
rect 1968 13066 2032 13130
rect 2049 13066 2113 13130
rect 2130 13066 2194 13130
rect 2211 13066 2275 13130
rect 2292 13066 2356 13130
rect 2373 13066 2437 13130
rect 2454 13066 2518 13130
rect 2535 13066 2599 13130
rect 2616 13066 2680 13130
rect 2697 13066 2761 13130
rect 2778 13066 2842 13130
rect 2859 13066 2923 13130
rect 2940 13066 3004 13130
rect 3021 13066 3085 13130
rect 3102 13066 3166 13130
rect 3183 13066 3247 13130
rect 3264 13066 3328 13130
rect 3345 13066 3409 13130
rect 3426 13066 3490 13130
rect 3507 13066 3571 13130
rect 3588 13066 3652 13130
rect 3669 13066 3733 13130
rect 3750 13066 3814 13130
rect 3831 13066 3895 13130
rect 3912 13066 3976 13130
rect 3993 13066 4057 13130
rect 4074 13066 4138 13130
rect 4155 13066 4219 13130
rect 4236 13066 4300 13130
rect 4317 13066 4381 13130
rect 4399 13066 4463 13130
rect 4481 13066 4545 13130
rect 4563 13066 4627 13130
rect 4645 13066 4709 13130
rect 4727 13066 4791 13130
rect 4809 13066 4873 13130
rect 105 12984 169 13048
rect 186 12984 250 13048
rect 267 12984 331 13048
rect 348 12984 412 13048
rect 429 12984 493 13048
rect 510 12984 574 13048
rect 591 12984 655 13048
rect 672 12984 736 13048
rect 753 12984 817 13048
rect 834 12984 898 13048
rect 915 12984 979 13048
rect 996 12984 1060 13048
rect 1077 12984 1141 13048
rect 1158 12984 1222 13048
rect 1239 12984 1303 13048
rect 1320 12984 1384 13048
rect 1401 12984 1465 13048
rect 1482 12984 1546 13048
rect 1563 12984 1627 13048
rect 1644 12984 1708 13048
rect 1725 12984 1789 13048
rect 1806 12984 1870 13048
rect 1887 12984 1951 13048
rect 1968 12984 2032 13048
rect 2049 12984 2113 13048
rect 2130 12984 2194 13048
rect 2211 12984 2275 13048
rect 2292 12984 2356 13048
rect 2373 12984 2437 13048
rect 2454 12984 2518 13048
rect 2535 12984 2599 13048
rect 2616 12984 2680 13048
rect 2697 12984 2761 13048
rect 2778 12984 2842 13048
rect 2859 12984 2923 13048
rect 2940 12984 3004 13048
rect 3021 12984 3085 13048
rect 3102 12984 3166 13048
rect 3183 12984 3247 13048
rect 3264 12984 3328 13048
rect 3345 12984 3409 13048
rect 3426 12984 3490 13048
rect 3507 12984 3571 13048
rect 3588 12984 3652 13048
rect 3669 12984 3733 13048
rect 3750 12984 3814 13048
rect 3831 12984 3895 13048
rect 3912 12984 3976 13048
rect 3993 12984 4057 13048
rect 4074 12984 4138 13048
rect 4155 12984 4219 13048
rect 4236 12984 4300 13048
rect 4317 12984 4381 13048
rect 4399 12984 4463 13048
rect 4481 12984 4545 13048
rect 4563 12984 4627 13048
rect 4645 12984 4709 13048
rect 4727 12984 4791 13048
rect 4809 12984 4873 13048
rect 105 12902 169 12966
rect 186 12902 250 12966
rect 267 12902 331 12966
rect 348 12902 412 12966
rect 429 12902 493 12966
rect 510 12902 574 12966
rect 591 12902 655 12966
rect 672 12902 736 12966
rect 753 12902 817 12966
rect 834 12902 898 12966
rect 915 12902 979 12966
rect 996 12902 1060 12966
rect 1077 12902 1141 12966
rect 1158 12902 1222 12966
rect 1239 12902 1303 12966
rect 1320 12902 1384 12966
rect 1401 12902 1465 12966
rect 1482 12902 1546 12966
rect 1563 12902 1627 12966
rect 1644 12902 1708 12966
rect 1725 12902 1789 12966
rect 1806 12902 1870 12966
rect 1887 12902 1951 12966
rect 1968 12902 2032 12966
rect 2049 12902 2113 12966
rect 2130 12902 2194 12966
rect 2211 12902 2275 12966
rect 2292 12902 2356 12966
rect 2373 12902 2437 12966
rect 2454 12902 2518 12966
rect 2535 12902 2599 12966
rect 2616 12902 2680 12966
rect 2697 12902 2761 12966
rect 2778 12902 2842 12966
rect 2859 12902 2923 12966
rect 2940 12902 3004 12966
rect 3021 12902 3085 12966
rect 3102 12902 3166 12966
rect 3183 12902 3247 12966
rect 3264 12902 3328 12966
rect 3345 12902 3409 12966
rect 3426 12902 3490 12966
rect 3507 12902 3571 12966
rect 3588 12902 3652 12966
rect 3669 12902 3733 12966
rect 3750 12902 3814 12966
rect 3831 12902 3895 12966
rect 3912 12902 3976 12966
rect 3993 12902 4057 12966
rect 4074 12902 4138 12966
rect 4155 12902 4219 12966
rect 4236 12902 4300 12966
rect 4317 12902 4381 12966
rect 4399 12902 4463 12966
rect 4481 12902 4545 12966
rect 4563 12902 4627 12966
rect 4645 12902 4709 12966
rect 4727 12902 4791 12966
rect 4809 12902 4873 12966
rect 105 12820 169 12884
rect 186 12820 250 12884
rect 267 12820 331 12884
rect 348 12820 412 12884
rect 429 12820 493 12884
rect 510 12820 574 12884
rect 591 12820 655 12884
rect 672 12820 736 12884
rect 753 12820 817 12884
rect 834 12820 898 12884
rect 915 12820 979 12884
rect 996 12820 1060 12884
rect 1077 12820 1141 12884
rect 1158 12820 1222 12884
rect 1239 12820 1303 12884
rect 1320 12820 1384 12884
rect 1401 12820 1465 12884
rect 1482 12820 1546 12884
rect 1563 12820 1627 12884
rect 1644 12820 1708 12884
rect 1725 12820 1789 12884
rect 1806 12820 1870 12884
rect 1887 12820 1951 12884
rect 1968 12820 2032 12884
rect 2049 12820 2113 12884
rect 2130 12820 2194 12884
rect 2211 12820 2275 12884
rect 2292 12820 2356 12884
rect 2373 12820 2437 12884
rect 2454 12820 2518 12884
rect 2535 12820 2599 12884
rect 2616 12820 2680 12884
rect 2697 12820 2761 12884
rect 2778 12820 2842 12884
rect 2859 12820 2923 12884
rect 2940 12820 3004 12884
rect 3021 12820 3085 12884
rect 3102 12820 3166 12884
rect 3183 12820 3247 12884
rect 3264 12820 3328 12884
rect 3345 12820 3409 12884
rect 3426 12820 3490 12884
rect 3507 12820 3571 12884
rect 3588 12820 3652 12884
rect 3669 12820 3733 12884
rect 3750 12820 3814 12884
rect 3831 12820 3895 12884
rect 3912 12820 3976 12884
rect 3993 12820 4057 12884
rect 4074 12820 4138 12884
rect 4155 12820 4219 12884
rect 4236 12820 4300 12884
rect 4317 12820 4381 12884
rect 4399 12820 4463 12884
rect 4481 12820 4545 12884
rect 4563 12820 4627 12884
rect 4645 12820 4709 12884
rect 4727 12820 4791 12884
rect 4809 12820 4873 12884
rect 10084 13640 10148 13704
rect 10165 13640 10229 13704
rect 10246 13640 10310 13704
rect 10327 13640 10391 13704
rect 10408 13640 10472 13704
rect 10489 13640 10553 13704
rect 10570 13640 10634 13704
rect 10651 13640 10715 13704
rect 10732 13640 10796 13704
rect 10813 13640 10877 13704
rect 10894 13640 10958 13704
rect 10975 13640 11039 13704
rect 11056 13640 11120 13704
rect 11137 13640 11201 13704
rect 11218 13640 11282 13704
rect 11299 13640 11363 13704
rect 11380 13640 11444 13704
rect 11461 13640 11525 13704
rect 11542 13640 11606 13704
rect 11623 13640 11687 13704
rect 11704 13640 11768 13704
rect 11785 13640 11849 13704
rect 11866 13640 11930 13704
rect 11947 13640 12011 13704
rect 12028 13640 12092 13704
rect 12109 13640 12173 13704
rect 12190 13640 12254 13704
rect 12271 13640 12335 13704
rect 12352 13640 12416 13704
rect 12433 13640 12497 13704
rect 12514 13640 12578 13704
rect 12595 13640 12659 13704
rect 12676 13640 12740 13704
rect 12757 13640 12821 13704
rect 12838 13640 12902 13704
rect 12919 13640 12983 13704
rect 13000 13640 13064 13704
rect 13081 13640 13145 13704
rect 13162 13640 13226 13704
rect 13243 13640 13307 13704
rect 13324 13640 13388 13704
rect 13405 13640 13469 13704
rect 13486 13640 13550 13704
rect 13567 13640 13631 13704
rect 13648 13640 13712 13704
rect 13729 13640 13793 13704
rect 13810 13640 13874 13704
rect 13891 13640 13955 13704
rect 13972 13640 14036 13704
rect 14053 13640 14117 13704
rect 14134 13640 14198 13704
rect 14215 13640 14279 13704
rect 14296 13640 14360 13704
rect 14378 13640 14442 13704
rect 14460 13640 14524 13704
rect 14542 13640 14606 13704
rect 14624 13640 14688 13704
rect 14706 13640 14770 13704
rect 14788 13640 14852 13704
rect 10084 13558 10148 13622
rect 10165 13558 10229 13622
rect 10246 13558 10310 13622
rect 10327 13558 10391 13622
rect 10408 13558 10472 13622
rect 10489 13558 10553 13622
rect 10570 13558 10634 13622
rect 10651 13558 10715 13622
rect 10732 13558 10796 13622
rect 10813 13558 10877 13622
rect 10894 13558 10958 13622
rect 10975 13558 11039 13622
rect 11056 13558 11120 13622
rect 11137 13558 11201 13622
rect 11218 13558 11282 13622
rect 11299 13558 11363 13622
rect 11380 13558 11444 13622
rect 11461 13558 11525 13622
rect 11542 13558 11606 13622
rect 11623 13558 11687 13622
rect 11704 13558 11768 13622
rect 11785 13558 11849 13622
rect 11866 13558 11930 13622
rect 11947 13558 12011 13622
rect 12028 13558 12092 13622
rect 12109 13558 12173 13622
rect 12190 13558 12254 13622
rect 12271 13558 12335 13622
rect 12352 13558 12416 13622
rect 12433 13558 12497 13622
rect 12514 13558 12578 13622
rect 12595 13558 12659 13622
rect 12676 13558 12740 13622
rect 12757 13558 12821 13622
rect 12838 13558 12902 13622
rect 12919 13558 12983 13622
rect 13000 13558 13064 13622
rect 13081 13558 13145 13622
rect 13162 13558 13226 13622
rect 13243 13558 13307 13622
rect 13324 13558 13388 13622
rect 13405 13558 13469 13622
rect 13486 13558 13550 13622
rect 13567 13558 13631 13622
rect 13648 13558 13712 13622
rect 13729 13558 13793 13622
rect 13810 13558 13874 13622
rect 13891 13558 13955 13622
rect 13972 13558 14036 13622
rect 14053 13558 14117 13622
rect 14134 13558 14198 13622
rect 14215 13558 14279 13622
rect 14296 13558 14360 13622
rect 14378 13558 14442 13622
rect 14460 13558 14524 13622
rect 14542 13558 14606 13622
rect 14624 13558 14688 13622
rect 14706 13558 14770 13622
rect 14788 13558 14852 13622
rect 10084 13476 10148 13540
rect 10165 13476 10229 13540
rect 10246 13476 10310 13540
rect 10327 13476 10391 13540
rect 10408 13476 10472 13540
rect 10489 13476 10553 13540
rect 10570 13476 10634 13540
rect 10651 13476 10715 13540
rect 10732 13476 10796 13540
rect 10813 13476 10877 13540
rect 10894 13476 10958 13540
rect 10975 13476 11039 13540
rect 11056 13476 11120 13540
rect 11137 13476 11201 13540
rect 11218 13476 11282 13540
rect 11299 13476 11363 13540
rect 11380 13476 11444 13540
rect 11461 13476 11525 13540
rect 11542 13476 11606 13540
rect 11623 13476 11687 13540
rect 11704 13476 11768 13540
rect 11785 13476 11849 13540
rect 11866 13476 11930 13540
rect 11947 13476 12011 13540
rect 12028 13476 12092 13540
rect 12109 13476 12173 13540
rect 12190 13476 12254 13540
rect 12271 13476 12335 13540
rect 12352 13476 12416 13540
rect 12433 13476 12497 13540
rect 12514 13476 12578 13540
rect 12595 13476 12659 13540
rect 12676 13476 12740 13540
rect 12757 13476 12821 13540
rect 12838 13476 12902 13540
rect 12919 13476 12983 13540
rect 13000 13476 13064 13540
rect 13081 13476 13145 13540
rect 13162 13476 13226 13540
rect 13243 13476 13307 13540
rect 13324 13476 13388 13540
rect 13405 13476 13469 13540
rect 13486 13476 13550 13540
rect 13567 13476 13631 13540
rect 13648 13476 13712 13540
rect 13729 13476 13793 13540
rect 13810 13476 13874 13540
rect 13891 13476 13955 13540
rect 13972 13476 14036 13540
rect 14053 13476 14117 13540
rect 14134 13476 14198 13540
rect 14215 13476 14279 13540
rect 14296 13476 14360 13540
rect 14378 13476 14442 13540
rect 14460 13476 14524 13540
rect 14542 13476 14606 13540
rect 14624 13476 14688 13540
rect 14706 13476 14770 13540
rect 14788 13476 14852 13540
rect 10084 13394 10148 13458
rect 10165 13394 10229 13458
rect 10246 13394 10310 13458
rect 10327 13394 10391 13458
rect 10408 13394 10472 13458
rect 10489 13394 10553 13458
rect 10570 13394 10634 13458
rect 10651 13394 10715 13458
rect 10732 13394 10796 13458
rect 10813 13394 10877 13458
rect 10894 13394 10958 13458
rect 10975 13394 11039 13458
rect 11056 13394 11120 13458
rect 11137 13394 11201 13458
rect 11218 13394 11282 13458
rect 11299 13394 11363 13458
rect 11380 13394 11444 13458
rect 11461 13394 11525 13458
rect 11542 13394 11606 13458
rect 11623 13394 11687 13458
rect 11704 13394 11768 13458
rect 11785 13394 11849 13458
rect 11866 13394 11930 13458
rect 11947 13394 12011 13458
rect 12028 13394 12092 13458
rect 12109 13394 12173 13458
rect 12190 13394 12254 13458
rect 12271 13394 12335 13458
rect 12352 13394 12416 13458
rect 12433 13394 12497 13458
rect 12514 13394 12578 13458
rect 12595 13394 12659 13458
rect 12676 13394 12740 13458
rect 12757 13394 12821 13458
rect 12838 13394 12902 13458
rect 12919 13394 12983 13458
rect 13000 13394 13064 13458
rect 13081 13394 13145 13458
rect 13162 13394 13226 13458
rect 13243 13394 13307 13458
rect 13324 13394 13388 13458
rect 13405 13394 13469 13458
rect 13486 13394 13550 13458
rect 13567 13394 13631 13458
rect 13648 13394 13712 13458
rect 13729 13394 13793 13458
rect 13810 13394 13874 13458
rect 13891 13394 13955 13458
rect 13972 13394 14036 13458
rect 14053 13394 14117 13458
rect 14134 13394 14198 13458
rect 14215 13394 14279 13458
rect 14296 13394 14360 13458
rect 14378 13394 14442 13458
rect 14460 13394 14524 13458
rect 14542 13394 14606 13458
rect 14624 13394 14688 13458
rect 14706 13394 14770 13458
rect 14788 13394 14852 13458
rect 10084 13312 10148 13376
rect 10165 13312 10229 13376
rect 10246 13312 10310 13376
rect 10327 13312 10391 13376
rect 10408 13312 10472 13376
rect 10489 13312 10553 13376
rect 10570 13312 10634 13376
rect 10651 13312 10715 13376
rect 10732 13312 10796 13376
rect 10813 13312 10877 13376
rect 10894 13312 10958 13376
rect 10975 13312 11039 13376
rect 11056 13312 11120 13376
rect 11137 13312 11201 13376
rect 11218 13312 11282 13376
rect 11299 13312 11363 13376
rect 11380 13312 11444 13376
rect 11461 13312 11525 13376
rect 11542 13312 11606 13376
rect 11623 13312 11687 13376
rect 11704 13312 11768 13376
rect 11785 13312 11849 13376
rect 11866 13312 11930 13376
rect 11947 13312 12011 13376
rect 12028 13312 12092 13376
rect 12109 13312 12173 13376
rect 12190 13312 12254 13376
rect 12271 13312 12335 13376
rect 12352 13312 12416 13376
rect 12433 13312 12497 13376
rect 12514 13312 12578 13376
rect 12595 13312 12659 13376
rect 12676 13312 12740 13376
rect 12757 13312 12821 13376
rect 12838 13312 12902 13376
rect 12919 13312 12983 13376
rect 13000 13312 13064 13376
rect 13081 13312 13145 13376
rect 13162 13312 13226 13376
rect 13243 13312 13307 13376
rect 13324 13312 13388 13376
rect 13405 13312 13469 13376
rect 13486 13312 13550 13376
rect 13567 13312 13631 13376
rect 13648 13312 13712 13376
rect 13729 13312 13793 13376
rect 13810 13312 13874 13376
rect 13891 13312 13955 13376
rect 13972 13312 14036 13376
rect 14053 13312 14117 13376
rect 14134 13312 14198 13376
rect 14215 13312 14279 13376
rect 14296 13312 14360 13376
rect 14378 13312 14442 13376
rect 14460 13312 14524 13376
rect 14542 13312 14606 13376
rect 14624 13312 14688 13376
rect 14706 13312 14770 13376
rect 14788 13312 14852 13376
rect 10084 13230 10148 13294
rect 10165 13230 10229 13294
rect 10246 13230 10310 13294
rect 10327 13230 10391 13294
rect 10408 13230 10472 13294
rect 10489 13230 10553 13294
rect 10570 13230 10634 13294
rect 10651 13230 10715 13294
rect 10732 13230 10796 13294
rect 10813 13230 10877 13294
rect 10894 13230 10958 13294
rect 10975 13230 11039 13294
rect 11056 13230 11120 13294
rect 11137 13230 11201 13294
rect 11218 13230 11282 13294
rect 11299 13230 11363 13294
rect 11380 13230 11444 13294
rect 11461 13230 11525 13294
rect 11542 13230 11606 13294
rect 11623 13230 11687 13294
rect 11704 13230 11768 13294
rect 11785 13230 11849 13294
rect 11866 13230 11930 13294
rect 11947 13230 12011 13294
rect 12028 13230 12092 13294
rect 12109 13230 12173 13294
rect 12190 13230 12254 13294
rect 12271 13230 12335 13294
rect 12352 13230 12416 13294
rect 12433 13230 12497 13294
rect 12514 13230 12578 13294
rect 12595 13230 12659 13294
rect 12676 13230 12740 13294
rect 12757 13230 12821 13294
rect 12838 13230 12902 13294
rect 12919 13230 12983 13294
rect 13000 13230 13064 13294
rect 13081 13230 13145 13294
rect 13162 13230 13226 13294
rect 13243 13230 13307 13294
rect 13324 13230 13388 13294
rect 13405 13230 13469 13294
rect 13486 13230 13550 13294
rect 13567 13230 13631 13294
rect 13648 13230 13712 13294
rect 13729 13230 13793 13294
rect 13810 13230 13874 13294
rect 13891 13230 13955 13294
rect 13972 13230 14036 13294
rect 14053 13230 14117 13294
rect 14134 13230 14198 13294
rect 14215 13230 14279 13294
rect 14296 13230 14360 13294
rect 14378 13230 14442 13294
rect 14460 13230 14524 13294
rect 14542 13230 14606 13294
rect 14624 13230 14688 13294
rect 14706 13230 14770 13294
rect 14788 13230 14852 13294
rect 10084 13148 10148 13212
rect 10165 13148 10229 13212
rect 10246 13148 10310 13212
rect 10327 13148 10391 13212
rect 10408 13148 10472 13212
rect 10489 13148 10553 13212
rect 10570 13148 10634 13212
rect 10651 13148 10715 13212
rect 10732 13148 10796 13212
rect 10813 13148 10877 13212
rect 10894 13148 10958 13212
rect 10975 13148 11039 13212
rect 11056 13148 11120 13212
rect 11137 13148 11201 13212
rect 11218 13148 11282 13212
rect 11299 13148 11363 13212
rect 11380 13148 11444 13212
rect 11461 13148 11525 13212
rect 11542 13148 11606 13212
rect 11623 13148 11687 13212
rect 11704 13148 11768 13212
rect 11785 13148 11849 13212
rect 11866 13148 11930 13212
rect 11947 13148 12011 13212
rect 12028 13148 12092 13212
rect 12109 13148 12173 13212
rect 12190 13148 12254 13212
rect 12271 13148 12335 13212
rect 12352 13148 12416 13212
rect 12433 13148 12497 13212
rect 12514 13148 12578 13212
rect 12595 13148 12659 13212
rect 12676 13148 12740 13212
rect 12757 13148 12821 13212
rect 12838 13148 12902 13212
rect 12919 13148 12983 13212
rect 13000 13148 13064 13212
rect 13081 13148 13145 13212
rect 13162 13148 13226 13212
rect 13243 13148 13307 13212
rect 13324 13148 13388 13212
rect 13405 13148 13469 13212
rect 13486 13148 13550 13212
rect 13567 13148 13631 13212
rect 13648 13148 13712 13212
rect 13729 13148 13793 13212
rect 13810 13148 13874 13212
rect 13891 13148 13955 13212
rect 13972 13148 14036 13212
rect 14053 13148 14117 13212
rect 14134 13148 14198 13212
rect 14215 13148 14279 13212
rect 14296 13148 14360 13212
rect 14378 13148 14442 13212
rect 14460 13148 14524 13212
rect 14542 13148 14606 13212
rect 14624 13148 14688 13212
rect 14706 13148 14770 13212
rect 14788 13148 14852 13212
rect 10084 13066 10148 13130
rect 10165 13066 10229 13130
rect 10246 13066 10310 13130
rect 10327 13066 10391 13130
rect 10408 13066 10472 13130
rect 10489 13066 10553 13130
rect 10570 13066 10634 13130
rect 10651 13066 10715 13130
rect 10732 13066 10796 13130
rect 10813 13066 10877 13130
rect 10894 13066 10958 13130
rect 10975 13066 11039 13130
rect 11056 13066 11120 13130
rect 11137 13066 11201 13130
rect 11218 13066 11282 13130
rect 11299 13066 11363 13130
rect 11380 13066 11444 13130
rect 11461 13066 11525 13130
rect 11542 13066 11606 13130
rect 11623 13066 11687 13130
rect 11704 13066 11768 13130
rect 11785 13066 11849 13130
rect 11866 13066 11930 13130
rect 11947 13066 12011 13130
rect 12028 13066 12092 13130
rect 12109 13066 12173 13130
rect 12190 13066 12254 13130
rect 12271 13066 12335 13130
rect 12352 13066 12416 13130
rect 12433 13066 12497 13130
rect 12514 13066 12578 13130
rect 12595 13066 12659 13130
rect 12676 13066 12740 13130
rect 12757 13066 12821 13130
rect 12838 13066 12902 13130
rect 12919 13066 12983 13130
rect 13000 13066 13064 13130
rect 13081 13066 13145 13130
rect 13162 13066 13226 13130
rect 13243 13066 13307 13130
rect 13324 13066 13388 13130
rect 13405 13066 13469 13130
rect 13486 13066 13550 13130
rect 13567 13066 13631 13130
rect 13648 13066 13712 13130
rect 13729 13066 13793 13130
rect 13810 13066 13874 13130
rect 13891 13066 13955 13130
rect 13972 13066 14036 13130
rect 14053 13066 14117 13130
rect 14134 13066 14198 13130
rect 14215 13066 14279 13130
rect 14296 13066 14360 13130
rect 14378 13066 14442 13130
rect 14460 13066 14524 13130
rect 14542 13066 14606 13130
rect 14624 13066 14688 13130
rect 14706 13066 14770 13130
rect 14788 13066 14852 13130
rect 10084 12984 10148 13048
rect 10165 12984 10229 13048
rect 10246 12984 10310 13048
rect 10327 12984 10391 13048
rect 10408 12984 10472 13048
rect 10489 12984 10553 13048
rect 10570 12984 10634 13048
rect 10651 12984 10715 13048
rect 10732 12984 10796 13048
rect 10813 12984 10877 13048
rect 10894 12984 10958 13048
rect 10975 12984 11039 13048
rect 11056 12984 11120 13048
rect 11137 12984 11201 13048
rect 11218 12984 11282 13048
rect 11299 12984 11363 13048
rect 11380 12984 11444 13048
rect 11461 12984 11525 13048
rect 11542 12984 11606 13048
rect 11623 12984 11687 13048
rect 11704 12984 11768 13048
rect 11785 12984 11849 13048
rect 11866 12984 11930 13048
rect 11947 12984 12011 13048
rect 12028 12984 12092 13048
rect 12109 12984 12173 13048
rect 12190 12984 12254 13048
rect 12271 12984 12335 13048
rect 12352 12984 12416 13048
rect 12433 12984 12497 13048
rect 12514 12984 12578 13048
rect 12595 12984 12659 13048
rect 12676 12984 12740 13048
rect 12757 12984 12821 13048
rect 12838 12984 12902 13048
rect 12919 12984 12983 13048
rect 13000 12984 13064 13048
rect 13081 12984 13145 13048
rect 13162 12984 13226 13048
rect 13243 12984 13307 13048
rect 13324 12984 13388 13048
rect 13405 12984 13469 13048
rect 13486 12984 13550 13048
rect 13567 12984 13631 13048
rect 13648 12984 13712 13048
rect 13729 12984 13793 13048
rect 13810 12984 13874 13048
rect 13891 12984 13955 13048
rect 13972 12984 14036 13048
rect 14053 12984 14117 13048
rect 14134 12984 14198 13048
rect 14215 12984 14279 13048
rect 14296 12984 14360 13048
rect 14378 12984 14442 13048
rect 14460 12984 14524 13048
rect 14542 12984 14606 13048
rect 14624 12984 14688 13048
rect 14706 12984 14770 13048
rect 14788 12984 14852 13048
rect 10084 12902 10148 12966
rect 10165 12902 10229 12966
rect 10246 12902 10310 12966
rect 10327 12902 10391 12966
rect 10408 12902 10472 12966
rect 10489 12902 10553 12966
rect 10570 12902 10634 12966
rect 10651 12902 10715 12966
rect 10732 12902 10796 12966
rect 10813 12902 10877 12966
rect 10894 12902 10958 12966
rect 10975 12902 11039 12966
rect 11056 12902 11120 12966
rect 11137 12902 11201 12966
rect 11218 12902 11282 12966
rect 11299 12902 11363 12966
rect 11380 12902 11444 12966
rect 11461 12902 11525 12966
rect 11542 12902 11606 12966
rect 11623 12902 11687 12966
rect 11704 12902 11768 12966
rect 11785 12902 11849 12966
rect 11866 12902 11930 12966
rect 11947 12902 12011 12966
rect 12028 12902 12092 12966
rect 12109 12902 12173 12966
rect 12190 12902 12254 12966
rect 12271 12902 12335 12966
rect 12352 12902 12416 12966
rect 12433 12902 12497 12966
rect 12514 12902 12578 12966
rect 12595 12902 12659 12966
rect 12676 12902 12740 12966
rect 12757 12902 12821 12966
rect 12838 12902 12902 12966
rect 12919 12902 12983 12966
rect 13000 12902 13064 12966
rect 13081 12902 13145 12966
rect 13162 12902 13226 12966
rect 13243 12902 13307 12966
rect 13324 12902 13388 12966
rect 13405 12902 13469 12966
rect 13486 12902 13550 12966
rect 13567 12902 13631 12966
rect 13648 12902 13712 12966
rect 13729 12902 13793 12966
rect 13810 12902 13874 12966
rect 13891 12902 13955 12966
rect 13972 12902 14036 12966
rect 14053 12902 14117 12966
rect 14134 12902 14198 12966
rect 14215 12902 14279 12966
rect 14296 12902 14360 12966
rect 14378 12902 14442 12966
rect 14460 12902 14524 12966
rect 14542 12902 14606 12966
rect 14624 12902 14688 12966
rect 14706 12902 14770 12966
rect 14788 12902 14852 12966
rect 10084 12820 10148 12884
rect 10165 12820 10229 12884
rect 10246 12820 10310 12884
rect 10327 12820 10391 12884
rect 10408 12820 10472 12884
rect 10489 12820 10553 12884
rect 10570 12820 10634 12884
rect 10651 12820 10715 12884
rect 10732 12820 10796 12884
rect 10813 12820 10877 12884
rect 10894 12820 10958 12884
rect 10975 12820 11039 12884
rect 11056 12820 11120 12884
rect 11137 12820 11201 12884
rect 11218 12820 11282 12884
rect 11299 12820 11363 12884
rect 11380 12820 11444 12884
rect 11461 12820 11525 12884
rect 11542 12820 11606 12884
rect 11623 12820 11687 12884
rect 11704 12820 11768 12884
rect 11785 12820 11849 12884
rect 11866 12820 11930 12884
rect 11947 12820 12011 12884
rect 12028 12820 12092 12884
rect 12109 12820 12173 12884
rect 12190 12820 12254 12884
rect 12271 12820 12335 12884
rect 12352 12820 12416 12884
rect 12433 12820 12497 12884
rect 12514 12820 12578 12884
rect 12595 12820 12659 12884
rect 12676 12820 12740 12884
rect 12757 12820 12821 12884
rect 12838 12820 12902 12884
rect 12919 12820 12983 12884
rect 13000 12820 13064 12884
rect 13081 12820 13145 12884
rect 13162 12820 13226 12884
rect 13243 12820 13307 12884
rect 13324 12820 13388 12884
rect 13405 12820 13469 12884
rect 13486 12820 13550 12884
rect 13567 12820 13631 12884
rect 13648 12820 13712 12884
rect 13729 12820 13793 12884
rect 13810 12820 13874 12884
rect 13891 12820 13955 12884
rect 13972 12820 14036 12884
rect 14053 12820 14117 12884
rect 14134 12820 14198 12884
rect 14215 12820 14279 12884
rect 14296 12820 14360 12884
rect 14378 12820 14442 12884
rect 14460 12820 14524 12884
rect 14542 12820 14606 12884
rect 14624 12820 14688 12884
rect 14706 12820 14770 12884
rect 14788 12820 14852 12884
rect 105 4820 169 4884
rect 186 4820 250 4884
rect 267 4820 331 4884
rect 348 4820 412 4884
rect 429 4820 493 4884
rect 510 4820 574 4884
rect 591 4820 655 4884
rect 672 4820 736 4884
rect 753 4820 817 4884
rect 834 4820 898 4884
rect 915 4820 979 4884
rect 996 4820 1060 4884
rect 1077 4820 1141 4884
rect 1158 4820 1222 4884
rect 1239 4820 1303 4884
rect 1320 4820 1384 4884
rect 1401 4820 1465 4884
rect 1482 4820 1546 4884
rect 1563 4820 1627 4884
rect 1644 4820 1708 4884
rect 1725 4820 1789 4884
rect 1806 4820 1870 4884
rect 1887 4820 1951 4884
rect 1968 4820 2032 4884
rect 2049 4820 2113 4884
rect 2130 4820 2194 4884
rect 2211 4820 2275 4884
rect 2292 4820 2356 4884
rect 2373 4820 2437 4884
rect 2454 4820 2518 4884
rect 2535 4820 2599 4884
rect 2616 4820 2680 4884
rect 2697 4820 2761 4884
rect 2778 4820 2842 4884
rect 2859 4820 2923 4884
rect 2940 4820 3004 4884
rect 3021 4820 3085 4884
rect 3102 4820 3166 4884
rect 3183 4820 3247 4884
rect 3264 4820 3328 4884
rect 3345 4820 3409 4884
rect 3426 4820 3490 4884
rect 3507 4820 3571 4884
rect 3588 4820 3652 4884
rect 3669 4820 3733 4884
rect 3750 4820 3814 4884
rect 3831 4820 3895 4884
rect 3912 4820 3976 4884
rect 3993 4820 4057 4884
rect 4074 4820 4138 4884
rect 4155 4820 4219 4884
rect 4236 4820 4300 4884
rect 4317 4820 4381 4884
rect 4399 4820 4463 4884
rect 4481 4820 4545 4884
rect 4563 4820 4627 4884
rect 4645 4820 4709 4884
rect 4727 4820 4791 4884
rect 4809 4820 4873 4884
rect 105 4734 169 4798
rect 186 4734 250 4798
rect 267 4734 331 4798
rect 348 4734 412 4798
rect 429 4734 493 4798
rect 510 4734 574 4798
rect 591 4734 655 4798
rect 672 4734 736 4798
rect 753 4734 817 4798
rect 834 4734 898 4798
rect 915 4734 979 4798
rect 996 4734 1060 4798
rect 1077 4734 1141 4798
rect 1158 4734 1222 4798
rect 1239 4734 1303 4798
rect 1320 4734 1384 4798
rect 1401 4734 1465 4798
rect 1482 4734 1546 4798
rect 1563 4734 1627 4798
rect 1644 4734 1708 4798
rect 1725 4734 1789 4798
rect 1806 4734 1870 4798
rect 1887 4734 1951 4798
rect 1968 4734 2032 4798
rect 2049 4734 2113 4798
rect 2130 4734 2194 4798
rect 2211 4734 2275 4798
rect 2292 4734 2356 4798
rect 2373 4734 2437 4798
rect 2454 4734 2518 4798
rect 2535 4734 2599 4798
rect 2616 4734 2680 4798
rect 2697 4734 2761 4798
rect 2778 4734 2842 4798
rect 2859 4734 2923 4798
rect 2940 4734 3004 4798
rect 3021 4734 3085 4798
rect 3102 4734 3166 4798
rect 3183 4734 3247 4798
rect 3264 4734 3328 4798
rect 3345 4734 3409 4798
rect 3426 4734 3490 4798
rect 3507 4734 3571 4798
rect 3588 4734 3652 4798
rect 3669 4734 3733 4798
rect 3750 4734 3814 4798
rect 3831 4734 3895 4798
rect 3912 4734 3976 4798
rect 3993 4734 4057 4798
rect 4074 4734 4138 4798
rect 4155 4734 4219 4798
rect 4236 4734 4300 4798
rect 4317 4734 4381 4798
rect 4399 4734 4463 4798
rect 4481 4734 4545 4798
rect 4563 4734 4627 4798
rect 4645 4734 4709 4798
rect 4727 4734 4791 4798
rect 4809 4734 4873 4798
rect 105 4648 169 4712
rect 186 4648 250 4712
rect 267 4648 331 4712
rect 348 4648 412 4712
rect 429 4648 493 4712
rect 510 4648 574 4712
rect 591 4648 655 4712
rect 672 4648 736 4712
rect 753 4648 817 4712
rect 834 4648 898 4712
rect 915 4648 979 4712
rect 996 4648 1060 4712
rect 1077 4648 1141 4712
rect 1158 4648 1222 4712
rect 1239 4648 1303 4712
rect 1320 4648 1384 4712
rect 1401 4648 1465 4712
rect 1482 4648 1546 4712
rect 1563 4648 1627 4712
rect 1644 4648 1708 4712
rect 1725 4648 1789 4712
rect 1806 4648 1870 4712
rect 1887 4648 1951 4712
rect 1968 4648 2032 4712
rect 2049 4648 2113 4712
rect 2130 4648 2194 4712
rect 2211 4648 2275 4712
rect 2292 4648 2356 4712
rect 2373 4648 2437 4712
rect 2454 4648 2518 4712
rect 2535 4648 2599 4712
rect 2616 4648 2680 4712
rect 2697 4648 2761 4712
rect 2778 4648 2842 4712
rect 2859 4648 2923 4712
rect 2940 4648 3004 4712
rect 3021 4648 3085 4712
rect 3102 4648 3166 4712
rect 3183 4648 3247 4712
rect 3264 4648 3328 4712
rect 3345 4648 3409 4712
rect 3426 4648 3490 4712
rect 3507 4648 3571 4712
rect 3588 4648 3652 4712
rect 3669 4648 3733 4712
rect 3750 4648 3814 4712
rect 3831 4648 3895 4712
rect 3912 4648 3976 4712
rect 3993 4648 4057 4712
rect 4074 4648 4138 4712
rect 4155 4648 4219 4712
rect 4236 4648 4300 4712
rect 4317 4648 4381 4712
rect 4399 4648 4463 4712
rect 4481 4648 4545 4712
rect 4563 4648 4627 4712
rect 4645 4648 4709 4712
rect 4727 4648 4791 4712
rect 4809 4648 4873 4712
rect 105 4562 169 4626
rect 186 4562 250 4626
rect 267 4562 331 4626
rect 348 4562 412 4626
rect 429 4562 493 4626
rect 510 4562 574 4626
rect 591 4562 655 4626
rect 672 4562 736 4626
rect 753 4562 817 4626
rect 834 4562 898 4626
rect 915 4562 979 4626
rect 996 4562 1060 4626
rect 1077 4562 1141 4626
rect 1158 4562 1222 4626
rect 1239 4562 1303 4626
rect 1320 4562 1384 4626
rect 1401 4562 1465 4626
rect 1482 4562 1546 4626
rect 1563 4562 1627 4626
rect 1644 4562 1708 4626
rect 1725 4562 1789 4626
rect 1806 4562 1870 4626
rect 1887 4562 1951 4626
rect 1968 4562 2032 4626
rect 2049 4562 2113 4626
rect 2130 4562 2194 4626
rect 2211 4562 2275 4626
rect 2292 4562 2356 4626
rect 2373 4562 2437 4626
rect 2454 4562 2518 4626
rect 2535 4562 2599 4626
rect 2616 4562 2680 4626
rect 2697 4562 2761 4626
rect 2778 4562 2842 4626
rect 2859 4562 2923 4626
rect 2940 4562 3004 4626
rect 3021 4562 3085 4626
rect 3102 4562 3166 4626
rect 3183 4562 3247 4626
rect 3264 4562 3328 4626
rect 3345 4562 3409 4626
rect 3426 4562 3490 4626
rect 3507 4562 3571 4626
rect 3588 4562 3652 4626
rect 3669 4562 3733 4626
rect 3750 4562 3814 4626
rect 3831 4562 3895 4626
rect 3912 4562 3976 4626
rect 3993 4562 4057 4626
rect 4074 4562 4138 4626
rect 4155 4562 4219 4626
rect 4236 4562 4300 4626
rect 4317 4562 4381 4626
rect 4399 4562 4463 4626
rect 4481 4562 4545 4626
rect 4563 4562 4627 4626
rect 4645 4562 4709 4626
rect 4727 4562 4791 4626
rect 4809 4562 4873 4626
rect 105 4476 169 4540
rect 186 4476 250 4540
rect 267 4476 331 4540
rect 348 4476 412 4540
rect 429 4476 493 4540
rect 510 4476 574 4540
rect 591 4476 655 4540
rect 672 4476 736 4540
rect 753 4476 817 4540
rect 834 4476 898 4540
rect 915 4476 979 4540
rect 996 4476 1060 4540
rect 1077 4476 1141 4540
rect 1158 4476 1222 4540
rect 1239 4476 1303 4540
rect 1320 4476 1384 4540
rect 1401 4476 1465 4540
rect 1482 4476 1546 4540
rect 1563 4476 1627 4540
rect 1644 4476 1708 4540
rect 1725 4476 1789 4540
rect 1806 4476 1870 4540
rect 1887 4476 1951 4540
rect 1968 4476 2032 4540
rect 2049 4476 2113 4540
rect 2130 4476 2194 4540
rect 2211 4476 2275 4540
rect 2292 4476 2356 4540
rect 2373 4476 2437 4540
rect 2454 4476 2518 4540
rect 2535 4476 2599 4540
rect 2616 4476 2680 4540
rect 2697 4476 2761 4540
rect 2778 4476 2842 4540
rect 2859 4476 2923 4540
rect 2940 4476 3004 4540
rect 3021 4476 3085 4540
rect 3102 4476 3166 4540
rect 3183 4476 3247 4540
rect 3264 4476 3328 4540
rect 3345 4476 3409 4540
rect 3426 4476 3490 4540
rect 3507 4476 3571 4540
rect 3588 4476 3652 4540
rect 3669 4476 3733 4540
rect 3750 4476 3814 4540
rect 3831 4476 3895 4540
rect 3912 4476 3976 4540
rect 3993 4476 4057 4540
rect 4074 4476 4138 4540
rect 4155 4476 4219 4540
rect 4236 4476 4300 4540
rect 4317 4476 4381 4540
rect 4399 4476 4463 4540
rect 4481 4476 4545 4540
rect 4563 4476 4627 4540
rect 4645 4476 4709 4540
rect 4727 4476 4791 4540
rect 4809 4476 4873 4540
rect 105 4390 169 4454
rect 186 4390 250 4454
rect 267 4390 331 4454
rect 348 4390 412 4454
rect 429 4390 493 4454
rect 510 4390 574 4454
rect 591 4390 655 4454
rect 672 4390 736 4454
rect 753 4390 817 4454
rect 834 4390 898 4454
rect 915 4390 979 4454
rect 996 4390 1060 4454
rect 1077 4390 1141 4454
rect 1158 4390 1222 4454
rect 1239 4390 1303 4454
rect 1320 4390 1384 4454
rect 1401 4390 1465 4454
rect 1482 4390 1546 4454
rect 1563 4390 1627 4454
rect 1644 4390 1708 4454
rect 1725 4390 1789 4454
rect 1806 4390 1870 4454
rect 1887 4390 1951 4454
rect 1968 4390 2032 4454
rect 2049 4390 2113 4454
rect 2130 4390 2194 4454
rect 2211 4390 2275 4454
rect 2292 4390 2356 4454
rect 2373 4390 2437 4454
rect 2454 4390 2518 4454
rect 2535 4390 2599 4454
rect 2616 4390 2680 4454
rect 2697 4390 2761 4454
rect 2778 4390 2842 4454
rect 2859 4390 2923 4454
rect 2940 4390 3004 4454
rect 3021 4390 3085 4454
rect 3102 4390 3166 4454
rect 3183 4390 3247 4454
rect 3264 4390 3328 4454
rect 3345 4390 3409 4454
rect 3426 4390 3490 4454
rect 3507 4390 3571 4454
rect 3588 4390 3652 4454
rect 3669 4390 3733 4454
rect 3750 4390 3814 4454
rect 3831 4390 3895 4454
rect 3912 4390 3976 4454
rect 3993 4390 4057 4454
rect 4074 4390 4138 4454
rect 4155 4390 4219 4454
rect 4236 4390 4300 4454
rect 4317 4390 4381 4454
rect 4399 4390 4463 4454
rect 4481 4390 4545 4454
rect 4563 4390 4627 4454
rect 4645 4390 4709 4454
rect 4727 4390 4791 4454
rect 4809 4390 4873 4454
rect 105 4304 169 4368
rect 186 4304 250 4368
rect 267 4304 331 4368
rect 348 4304 412 4368
rect 429 4304 493 4368
rect 510 4304 574 4368
rect 591 4304 655 4368
rect 672 4304 736 4368
rect 753 4304 817 4368
rect 834 4304 898 4368
rect 915 4304 979 4368
rect 996 4304 1060 4368
rect 1077 4304 1141 4368
rect 1158 4304 1222 4368
rect 1239 4304 1303 4368
rect 1320 4304 1384 4368
rect 1401 4304 1465 4368
rect 1482 4304 1546 4368
rect 1563 4304 1627 4368
rect 1644 4304 1708 4368
rect 1725 4304 1789 4368
rect 1806 4304 1870 4368
rect 1887 4304 1951 4368
rect 1968 4304 2032 4368
rect 2049 4304 2113 4368
rect 2130 4304 2194 4368
rect 2211 4304 2275 4368
rect 2292 4304 2356 4368
rect 2373 4304 2437 4368
rect 2454 4304 2518 4368
rect 2535 4304 2599 4368
rect 2616 4304 2680 4368
rect 2697 4304 2761 4368
rect 2778 4304 2842 4368
rect 2859 4304 2923 4368
rect 2940 4304 3004 4368
rect 3021 4304 3085 4368
rect 3102 4304 3166 4368
rect 3183 4304 3247 4368
rect 3264 4304 3328 4368
rect 3345 4304 3409 4368
rect 3426 4304 3490 4368
rect 3507 4304 3571 4368
rect 3588 4304 3652 4368
rect 3669 4304 3733 4368
rect 3750 4304 3814 4368
rect 3831 4304 3895 4368
rect 3912 4304 3976 4368
rect 3993 4304 4057 4368
rect 4074 4304 4138 4368
rect 4155 4304 4219 4368
rect 4236 4304 4300 4368
rect 4317 4304 4381 4368
rect 4399 4304 4463 4368
rect 4481 4304 4545 4368
rect 4563 4304 4627 4368
rect 4645 4304 4709 4368
rect 4727 4304 4791 4368
rect 4809 4304 4873 4368
rect 105 4218 169 4282
rect 186 4218 250 4282
rect 267 4218 331 4282
rect 348 4218 412 4282
rect 429 4218 493 4282
rect 510 4218 574 4282
rect 591 4218 655 4282
rect 672 4218 736 4282
rect 753 4218 817 4282
rect 834 4218 898 4282
rect 915 4218 979 4282
rect 996 4218 1060 4282
rect 1077 4218 1141 4282
rect 1158 4218 1222 4282
rect 1239 4218 1303 4282
rect 1320 4218 1384 4282
rect 1401 4218 1465 4282
rect 1482 4218 1546 4282
rect 1563 4218 1627 4282
rect 1644 4218 1708 4282
rect 1725 4218 1789 4282
rect 1806 4218 1870 4282
rect 1887 4218 1951 4282
rect 1968 4218 2032 4282
rect 2049 4218 2113 4282
rect 2130 4218 2194 4282
rect 2211 4218 2275 4282
rect 2292 4218 2356 4282
rect 2373 4218 2437 4282
rect 2454 4218 2518 4282
rect 2535 4218 2599 4282
rect 2616 4218 2680 4282
rect 2697 4218 2761 4282
rect 2778 4218 2842 4282
rect 2859 4218 2923 4282
rect 2940 4218 3004 4282
rect 3021 4218 3085 4282
rect 3102 4218 3166 4282
rect 3183 4218 3247 4282
rect 3264 4218 3328 4282
rect 3345 4218 3409 4282
rect 3426 4218 3490 4282
rect 3507 4218 3571 4282
rect 3588 4218 3652 4282
rect 3669 4218 3733 4282
rect 3750 4218 3814 4282
rect 3831 4218 3895 4282
rect 3912 4218 3976 4282
rect 3993 4218 4057 4282
rect 4074 4218 4138 4282
rect 4155 4218 4219 4282
rect 4236 4218 4300 4282
rect 4317 4218 4381 4282
rect 4399 4218 4463 4282
rect 4481 4218 4545 4282
rect 4563 4218 4627 4282
rect 4645 4218 4709 4282
rect 4727 4218 4791 4282
rect 4809 4218 4873 4282
rect 105 4132 169 4196
rect 186 4132 250 4196
rect 267 4132 331 4196
rect 348 4132 412 4196
rect 429 4132 493 4196
rect 510 4132 574 4196
rect 591 4132 655 4196
rect 672 4132 736 4196
rect 753 4132 817 4196
rect 834 4132 898 4196
rect 915 4132 979 4196
rect 996 4132 1060 4196
rect 1077 4132 1141 4196
rect 1158 4132 1222 4196
rect 1239 4132 1303 4196
rect 1320 4132 1384 4196
rect 1401 4132 1465 4196
rect 1482 4132 1546 4196
rect 1563 4132 1627 4196
rect 1644 4132 1708 4196
rect 1725 4132 1789 4196
rect 1806 4132 1870 4196
rect 1887 4132 1951 4196
rect 1968 4132 2032 4196
rect 2049 4132 2113 4196
rect 2130 4132 2194 4196
rect 2211 4132 2275 4196
rect 2292 4132 2356 4196
rect 2373 4132 2437 4196
rect 2454 4132 2518 4196
rect 2535 4132 2599 4196
rect 2616 4132 2680 4196
rect 2697 4132 2761 4196
rect 2778 4132 2842 4196
rect 2859 4132 2923 4196
rect 2940 4132 3004 4196
rect 3021 4132 3085 4196
rect 3102 4132 3166 4196
rect 3183 4132 3247 4196
rect 3264 4132 3328 4196
rect 3345 4132 3409 4196
rect 3426 4132 3490 4196
rect 3507 4132 3571 4196
rect 3588 4132 3652 4196
rect 3669 4132 3733 4196
rect 3750 4132 3814 4196
rect 3831 4132 3895 4196
rect 3912 4132 3976 4196
rect 3993 4132 4057 4196
rect 4074 4132 4138 4196
rect 4155 4132 4219 4196
rect 4236 4132 4300 4196
rect 4317 4132 4381 4196
rect 4399 4132 4463 4196
rect 4481 4132 4545 4196
rect 4563 4132 4627 4196
rect 4645 4132 4709 4196
rect 4727 4132 4791 4196
rect 4809 4132 4873 4196
rect 105 4046 169 4110
rect 186 4046 250 4110
rect 267 4046 331 4110
rect 348 4046 412 4110
rect 429 4046 493 4110
rect 510 4046 574 4110
rect 591 4046 655 4110
rect 672 4046 736 4110
rect 753 4046 817 4110
rect 834 4046 898 4110
rect 915 4046 979 4110
rect 996 4046 1060 4110
rect 1077 4046 1141 4110
rect 1158 4046 1222 4110
rect 1239 4046 1303 4110
rect 1320 4046 1384 4110
rect 1401 4046 1465 4110
rect 1482 4046 1546 4110
rect 1563 4046 1627 4110
rect 1644 4046 1708 4110
rect 1725 4046 1789 4110
rect 1806 4046 1870 4110
rect 1887 4046 1951 4110
rect 1968 4046 2032 4110
rect 2049 4046 2113 4110
rect 2130 4046 2194 4110
rect 2211 4046 2275 4110
rect 2292 4046 2356 4110
rect 2373 4046 2437 4110
rect 2454 4046 2518 4110
rect 2535 4046 2599 4110
rect 2616 4046 2680 4110
rect 2697 4046 2761 4110
rect 2778 4046 2842 4110
rect 2859 4046 2923 4110
rect 2940 4046 3004 4110
rect 3021 4046 3085 4110
rect 3102 4046 3166 4110
rect 3183 4046 3247 4110
rect 3264 4046 3328 4110
rect 3345 4046 3409 4110
rect 3426 4046 3490 4110
rect 3507 4046 3571 4110
rect 3588 4046 3652 4110
rect 3669 4046 3733 4110
rect 3750 4046 3814 4110
rect 3831 4046 3895 4110
rect 3912 4046 3976 4110
rect 3993 4046 4057 4110
rect 4074 4046 4138 4110
rect 4155 4046 4219 4110
rect 4236 4046 4300 4110
rect 4317 4046 4381 4110
rect 4399 4046 4463 4110
rect 4481 4046 4545 4110
rect 4563 4046 4627 4110
rect 4645 4046 4709 4110
rect 4727 4046 4791 4110
rect 4809 4046 4873 4110
rect 105 3960 169 4024
rect 186 3960 250 4024
rect 267 3960 331 4024
rect 348 3960 412 4024
rect 429 3960 493 4024
rect 510 3960 574 4024
rect 591 3960 655 4024
rect 672 3960 736 4024
rect 753 3960 817 4024
rect 834 3960 898 4024
rect 915 3960 979 4024
rect 996 3960 1060 4024
rect 1077 3960 1141 4024
rect 1158 3960 1222 4024
rect 1239 3960 1303 4024
rect 1320 3960 1384 4024
rect 1401 3960 1465 4024
rect 1482 3960 1546 4024
rect 1563 3960 1627 4024
rect 1644 3960 1708 4024
rect 1725 3960 1789 4024
rect 1806 3960 1870 4024
rect 1887 3960 1951 4024
rect 1968 3960 2032 4024
rect 2049 3960 2113 4024
rect 2130 3960 2194 4024
rect 2211 3960 2275 4024
rect 2292 3960 2356 4024
rect 2373 3960 2437 4024
rect 2454 3960 2518 4024
rect 2535 3960 2599 4024
rect 2616 3960 2680 4024
rect 2697 3960 2761 4024
rect 2778 3960 2842 4024
rect 2859 3960 2923 4024
rect 2940 3960 3004 4024
rect 3021 3960 3085 4024
rect 3102 3960 3166 4024
rect 3183 3960 3247 4024
rect 3264 3960 3328 4024
rect 3345 3960 3409 4024
rect 3426 3960 3490 4024
rect 3507 3960 3571 4024
rect 3588 3960 3652 4024
rect 3669 3960 3733 4024
rect 3750 3960 3814 4024
rect 3831 3960 3895 4024
rect 3912 3960 3976 4024
rect 3993 3960 4057 4024
rect 4074 3960 4138 4024
rect 4155 3960 4219 4024
rect 4236 3960 4300 4024
rect 4317 3960 4381 4024
rect 4399 3960 4463 4024
rect 4481 3960 4545 4024
rect 4563 3960 4627 4024
rect 4645 3960 4709 4024
rect 4727 3960 4791 4024
rect 4809 3960 4873 4024
rect 10084 4820 10148 4884
rect 10165 4820 10229 4884
rect 10246 4820 10310 4884
rect 10327 4820 10391 4884
rect 10408 4820 10472 4884
rect 10489 4820 10553 4884
rect 10570 4820 10634 4884
rect 10651 4820 10715 4884
rect 10732 4820 10796 4884
rect 10813 4820 10877 4884
rect 10894 4820 10958 4884
rect 10975 4820 11039 4884
rect 11056 4820 11120 4884
rect 11137 4820 11201 4884
rect 11218 4820 11282 4884
rect 11299 4820 11363 4884
rect 11380 4820 11444 4884
rect 11461 4820 11525 4884
rect 11542 4820 11606 4884
rect 11623 4820 11687 4884
rect 11704 4820 11768 4884
rect 11785 4820 11849 4884
rect 11866 4820 11930 4884
rect 11947 4820 12011 4884
rect 12028 4820 12092 4884
rect 12109 4820 12173 4884
rect 12190 4820 12254 4884
rect 12271 4820 12335 4884
rect 12352 4820 12416 4884
rect 12433 4820 12497 4884
rect 12514 4820 12578 4884
rect 12595 4820 12659 4884
rect 12676 4820 12740 4884
rect 12757 4820 12821 4884
rect 12838 4820 12902 4884
rect 12919 4820 12983 4884
rect 13000 4820 13064 4884
rect 13081 4820 13145 4884
rect 13162 4820 13226 4884
rect 13243 4820 13307 4884
rect 13324 4820 13388 4884
rect 13405 4820 13469 4884
rect 13486 4820 13550 4884
rect 13567 4820 13631 4884
rect 13648 4820 13712 4884
rect 13729 4820 13793 4884
rect 13810 4820 13874 4884
rect 13891 4820 13955 4884
rect 13972 4820 14036 4884
rect 14053 4820 14117 4884
rect 14134 4820 14198 4884
rect 14215 4820 14279 4884
rect 14296 4820 14360 4884
rect 14378 4820 14442 4884
rect 14460 4820 14524 4884
rect 14542 4820 14606 4884
rect 14624 4820 14688 4884
rect 14706 4820 14770 4884
rect 14788 4820 14852 4884
rect 10084 4734 10148 4798
rect 10165 4734 10229 4798
rect 10246 4734 10310 4798
rect 10327 4734 10391 4798
rect 10408 4734 10472 4798
rect 10489 4734 10553 4798
rect 10570 4734 10634 4798
rect 10651 4734 10715 4798
rect 10732 4734 10796 4798
rect 10813 4734 10877 4798
rect 10894 4734 10958 4798
rect 10975 4734 11039 4798
rect 11056 4734 11120 4798
rect 11137 4734 11201 4798
rect 11218 4734 11282 4798
rect 11299 4734 11363 4798
rect 11380 4734 11444 4798
rect 11461 4734 11525 4798
rect 11542 4734 11606 4798
rect 11623 4734 11687 4798
rect 11704 4734 11768 4798
rect 11785 4734 11849 4798
rect 11866 4734 11930 4798
rect 11947 4734 12011 4798
rect 12028 4734 12092 4798
rect 12109 4734 12173 4798
rect 12190 4734 12254 4798
rect 12271 4734 12335 4798
rect 12352 4734 12416 4798
rect 12433 4734 12497 4798
rect 12514 4734 12578 4798
rect 12595 4734 12659 4798
rect 12676 4734 12740 4798
rect 12757 4734 12821 4798
rect 12838 4734 12902 4798
rect 12919 4734 12983 4798
rect 13000 4734 13064 4798
rect 13081 4734 13145 4798
rect 13162 4734 13226 4798
rect 13243 4734 13307 4798
rect 13324 4734 13388 4798
rect 13405 4734 13469 4798
rect 13486 4734 13550 4798
rect 13567 4734 13631 4798
rect 13648 4734 13712 4798
rect 13729 4734 13793 4798
rect 13810 4734 13874 4798
rect 13891 4734 13955 4798
rect 13972 4734 14036 4798
rect 14053 4734 14117 4798
rect 14134 4734 14198 4798
rect 14215 4734 14279 4798
rect 14296 4734 14360 4798
rect 14378 4734 14442 4798
rect 14460 4734 14524 4798
rect 14542 4734 14606 4798
rect 14624 4734 14688 4798
rect 14706 4734 14770 4798
rect 14788 4734 14852 4798
rect 10084 4648 10148 4712
rect 10165 4648 10229 4712
rect 10246 4648 10310 4712
rect 10327 4648 10391 4712
rect 10408 4648 10472 4712
rect 10489 4648 10553 4712
rect 10570 4648 10634 4712
rect 10651 4648 10715 4712
rect 10732 4648 10796 4712
rect 10813 4648 10877 4712
rect 10894 4648 10958 4712
rect 10975 4648 11039 4712
rect 11056 4648 11120 4712
rect 11137 4648 11201 4712
rect 11218 4648 11282 4712
rect 11299 4648 11363 4712
rect 11380 4648 11444 4712
rect 11461 4648 11525 4712
rect 11542 4648 11606 4712
rect 11623 4648 11687 4712
rect 11704 4648 11768 4712
rect 11785 4648 11849 4712
rect 11866 4648 11930 4712
rect 11947 4648 12011 4712
rect 12028 4648 12092 4712
rect 12109 4648 12173 4712
rect 12190 4648 12254 4712
rect 12271 4648 12335 4712
rect 12352 4648 12416 4712
rect 12433 4648 12497 4712
rect 12514 4648 12578 4712
rect 12595 4648 12659 4712
rect 12676 4648 12740 4712
rect 12757 4648 12821 4712
rect 12838 4648 12902 4712
rect 12919 4648 12983 4712
rect 13000 4648 13064 4712
rect 13081 4648 13145 4712
rect 13162 4648 13226 4712
rect 13243 4648 13307 4712
rect 13324 4648 13388 4712
rect 13405 4648 13469 4712
rect 13486 4648 13550 4712
rect 13567 4648 13631 4712
rect 13648 4648 13712 4712
rect 13729 4648 13793 4712
rect 13810 4648 13874 4712
rect 13891 4648 13955 4712
rect 13972 4648 14036 4712
rect 14053 4648 14117 4712
rect 14134 4648 14198 4712
rect 14215 4648 14279 4712
rect 14296 4648 14360 4712
rect 14378 4648 14442 4712
rect 14460 4648 14524 4712
rect 14542 4648 14606 4712
rect 14624 4648 14688 4712
rect 14706 4648 14770 4712
rect 14788 4648 14852 4712
rect 10084 4562 10148 4626
rect 10165 4562 10229 4626
rect 10246 4562 10310 4626
rect 10327 4562 10391 4626
rect 10408 4562 10472 4626
rect 10489 4562 10553 4626
rect 10570 4562 10634 4626
rect 10651 4562 10715 4626
rect 10732 4562 10796 4626
rect 10813 4562 10877 4626
rect 10894 4562 10958 4626
rect 10975 4562 11039 4626
rect 11056 4562 11120 4626
rect 11137 4562 11201 4626
rect 11218 4562 11282 4626
rect 11299 4562 11363 4626
rect 11380 4562 11444 4626
rect 11461 4562 11525 4626
rect 11542 4562 11606 4626
rect 11623 4562 11687 4626
rect 11704 4562 11768 4626
rect 11785 4562 11849 4626
rect 11866 4562 11930 4626
rect 11947 4562 12011 4626
rect 12028 4562 12092 4626
rect 12109 4562 12173 4626
rect 12190 4562 12254 4626
rect 12271 4562 12335 4626
rect 12352 4562 12416 4626
rect 12433 4562 12497 4626
rect 12514 4562 12578 4626
rect 12595 4562 12659 4626
rect 12676 4562 12740 4626
rect 12757 4562 12821 4626
rect 12838 4562 12902 4626
rect 12919 4562 12983 4626
rect 13000 4562 13064 4626
rect 13081 4562 13145 4626
rect 13162 4562 13226 4626
rect 13243 4562 13307 4626
rect 13324 4562 13388 4626
rect 13405 4562 13469 4626
rect 13486 4562 13550 4626
rect 13567 4562 13631 4626
rect 13648 4562 13712 4626
rect 13729 4562 13793 4626
rect 13810 4562 13874 4626
rect 13891 4562 13955 4626
rect 13972 4562 14036 4626
rect 14053 4562 14117 4626
rect 14134 4562 14198 4626
rect 14215 4562 14279 4626
rect 14296 4562 14360 4626
rect 14378 4562 14442 4626
rect 14460 4562 14524 4626
rect 14542 4562 14606 4626
rect 14624 4562 14688 4626
rect 14706 4562 14770 4626
rect 14788 4562 14852 4626
rect 10084 4476 10148 4540
rect 10165 4476 10229 4540
rect 10246 4476 10310 4540
rect 10327 4476 10391 4540
rect 10408 4476 10472 4540
rect 10489 4476 10553 4540
rect 10570 4476 10634 4540
rect 10651 4476 10715 4540
rect 10732 4476 10796 4540
rect 10813 4476 10877 4540
rect 10894 4476 10958 4540
rect 10975 4476 11039 4540
rect 11056 4476 11120 4540
rect 11137 4476 11201 4540
rect 11218 4476 11282 4540
rect 11299 4476 11363 4540
rect 11380 4476 11444 4540
rect 11461 4476 11525 4540
rect 11542 4476 11606 4540
rect 11623 4476 11687 4540
rect 11704 4476 11768 4540
rect 11785 4476 11849 4540
rect 11866 4476 11930 4540
rect 11947 4476 12011 4540
rect 12028 4476 12092 4540
rect 12109 4476 12173 4540
rect 12190 4476 12254 4540
rect 12271 4476 12335 4540
rect 12352 4476 12416 4540
rect 12433 4476 12497 4540
rect 12514 4476 12578 4540
rect 12595 4476 12659 4540
rect 12676 4476 12740 4540
rect 12757 4476 12821 4540
rect 12838 4476 12902 4540
rect 12919 4476 12983 4540
rect 13000 4476 13064 4540
rect 13081 4476 13145 4540
rect 13162 4476 13226 4540
rect 13243 4476 13307 4540
rect 13324 4476 13388 4540
rect 13405 4476 13469 4540
rect 13486 4476 13550 4540
rect 13567 4476 13631 4540
rect 13648 4476 13712 4540
rect 13729 4476 13793 4540
rect 13810 4476 13874 4540
rect 13891 4476 13955 4540
rect 13972 4476 14036 4540
rect 14053 4476 14117 4540
rect 14134 4476 14198 4540
rect 14215 4476 14279 4540
rect 14296 4476 14360 4540
rect 14378 4476 14442 4540
rect 14460 4476 14524 4540
rect 14542 4476 14606 4540
rect 14624 4476 14688 4540
rect 14706 4476 14770 4540
rect 14788 4476 14852 4540
rect 10084 4390 10148 4454
rect 10165 4390 10229 4454
rect 10246 4390 10310 4454
rect 10327 4390 10391 4454
rect 10408 4390 10472 4454
rect 10489 4390 10553 4454
rect 10570 4390 10634 4454
rect 10651 4390 10715 4454
rect 10732 4390 10796 4454
rect 10813 4390 10877 4454
rect 10894 4390 10958 4454
rect 10975 4390 11039 4454
rect 11056 4390 11120 4454
rect 11137 4390 11201 4454
rect 11218 4390 11282 4454
rect 11299 4390 11363 4454
rect 11380 4390 11444 4454
rect 11461 4390 11525 4454
rect 11542 4390 11606 4454
rect 11623 4390 11687 4454
rect 11704 4390 11768 4454
rect 11785 4390 11849 4454
rect 11866 4390 11930 4454
rect 11947 4390 12011 4454
rect 12028 4390 12092 4454
rect 12109 4390 12173 4454
rect 12190 4390 12254 4454
rect 12271 4390 12335 4454
rect 12352 4390 12416 4454
rect 12433 4390 12497 4454
rect 12514 4390 12578 4454
rect 12595 4390 12659 4454
rect 12676 4390 12740 4454
rect 12757 4390 12821 4454
rect 12838 4390 12902 4454
rect 12919 4390 12983 4454
rect 13000 4390 13064 4454
rect 13081 4390 13145 4454
rect 13162 4390 13226 4454
rect 13243 4390 13307 4454
rect 13324 4390 13388 4454
rect 13405 4390 13469 4454
rect 13486 4390 13550 4454
rect 13567 4390 13631 4454
rect 13648 4390 13712 4454
rect 13729 4390 13793 4454
rect 13810 4390 13874 4454
rect 13891 4390 13955 4454
rect 13972 4390 14036 4454
rect 14053 4390 14117 4454
rect 14134 4390 14198 4454
rect 14215 4390 14279 4454
rect 14296 4390 14360 4454
rect 14378 4390 14442 4454
rect 14460 4390 14524 4454
rect 14542 4390 14606 4454
rect 14624 4390 14688 4454
rect 14706 4390 14770 4454
rect 14788 4390 14852 4454
rect 10084 4304 10148 4368
rect 10165 4304 10229 4368
rect 10246 4304 10310 4368
rect 10327 4304 10391 4368
rect 10408 4304 10472 4368
rect 10489 4304 10553 4368
rect 10570 4304 10634 4368
rect 10651 4304 10715 4368
rect 10732 4304 10796 4368
rect 10813 4304 10877 4368
rect 10894 4304 10958 4368
rect 10975 4304 11039 4368
rect 11056 4304 11120 4368
rect 11137 4304 11201 4368
rect 11218 4304 11282 4368
rect 11299 4304 11363 4368
rect 11380 4304 11444 4368
rect 11461 4304 11525 4368
rect 11542 4304 11606 4368
rect 11623 4304 11687 4368
rect 11704 4304 11768 4368
rect 11785 4304 11849 4368
rect 11866 4304 11930 4368
rect 11947 4304 12011 4368
rect 12028 4304 12092 4368
rect 12109 4304 12173 4368
rect 12190 4304 12254 4368
rect 12271 4304 12335 4368
rect 12352 4304 12416 4368
rect 12433 4304 12497 4368
rect 12514 4304 12578 4368
rect 12595 4304 12659 4368
rect 12676 4304 12740 4368
rect 12757 4304 12821 4368
rect 12838 4304 12902 4368
rect 12919 4304 12983 4368
rect 13000 4304 13064 4368
rect 13081 4304 13145 4368
rect 13162 4304 13226 4368
rect 13243 4304 13307 4368
rect 13324 4304 13388 4368
rect 13405 4304 13469 4368
rect 13486 4304 13550 4368
rect 13567 4304 13631 4368
rect 13648 4304 13712 4368
rect 13729 4304 13793 4368
rect 13810 4304 13874 4368
rect 13891 4304 13955 4368
rect 13972 4304 14036 4368
rect 14053 4304 14117 4368
rect 14134 4304 14198 4368
rect 14215 4304 14279 4368
rect 14296 4304 14360 4368
rect 14378 4304 14442 4368
rect 14460 4304 14524 4368
rect 14542 4304 14606 4368
rect 14624 4304 14688 4368
rect 14706 4304 14770 4368
rect 14788 4304 14852 4368
rect 10084 4218 10148 4282
rect 10165 4218 10229 4282
rect 10246 4218 10310 4282
rect 10327 4218 10391 4282
rect 10408 4218 10472 4282
rect 10489 4218 10553 4282
rect 10570 4218 10634 4282
rect 10651 4218 10715 4282
rect 10732 4218 10796 4282
rect 10813 4218 10877 4282
rect 10894 4218 10958 4282
rect 10975 4218 11039 4282
rect 11056 4218 11120 4282
rect 11137 4218 11201 4282
rect 11218 4218 11282 4282
rect 11299 4218 11363 4282
rect 11380 4218 11444 4282
rect 11461 4218 11525 4282
rect 11542 4218 11606 4282
rect 11623 4218 11687 4282
rect 11704 4218 11768 4282
rect 11785 4218 11849 4282
rect 11866 4218 11930 4282
rect 11947 4218 12011 4282
rect 12028 4218 12092 4282
rect 12109 4218 12173 4282
rect 12190 4218 12254 4282
rect 12271 4218 12335 4282
rect 12352 4218 12416 4282
rect 12433 4218 12497 4282
rect 12514 4218 12578 4282
rect 12595 4218 12659 4282
rect 12676 4218 12740 4282
rect 12757 4218 12821 4282
rect 12838 4218 12902 4282
rect 12919 4218 12983 4282
rect 13000 4218 13064 4282
rect 13081 4218 13145 4282
rect 13162 4218 13226 4282
rect 13243 4218 13307 4282
rect 13324 4218 13388 4282
rect 13405 4218 13469 4282
rect 13486 4218 13550 4282
rect 13567 4218 13631 4282
rect 13648 4218 13712 4282
rect 13729 4218 13793 4282
rect 13810 4218 13874 4282
rect 13891 4218 13955 4282
rect 13972 4218 14036 4282
rect 14053 4218 14117 4282
rect 14134 4218 14198 4282
rect 14215 4218 14279 4282
rect 14296 4218 14360 4282
rect 14378 4218 14442 4282
rect 14460 4218 14524 4282
rect 14542 4218 14606 4282
rect 14624 4218 14688 4282
rect 14706 4218 14770 4282
rect 14788 4218 14852 4282
rect 10084 4132 10148 4196
rect 10165 4132 10229 4196
rect 10246 4132 10310 4196
rect 10327 4132 10391 4196
rect 10408 4132 10472 4196
rect 10489 4132 10553 4196
rect 10570 4132 10634 4196
rect 10651 4132 10715 4196
rect 10732 4132 10796 4196
rect 10813 4132 10877 4196
rect 10894 4132 10958 4196
rect 10975 4132 11039 4196
rect 11056 4132 11120 4196
rect 11137 4132 11201 4196
rect 11218 4132 11282 4196
rect 11299 4132 11363 4196
rect 11380 4132 11444 4196
rect 11461 4132 11525 4196
rect 11542 4132 11606 4196
rect 11623 4132 11687 4196
rect 11704 4132 11768 4196
rect 11785 4132 11849 4196
rect 11866 4132 11930 4196
rect 11947 4132 12011 4196
rect 12028 4132 12092 4196
rect 12109 4132 12173 4196
rect 12190 4132 12254 4196
rect 12271 4132 12335 4196
rect 12352 4132 12416 4196
rect 12433 4132 12497 4196
rect 12514 4132 12578 4196
rect 12595 4132 12659 4196
rect 12676 4132 12740 4196
rect 12757 4132 12821 4196
rect 12838 4132 12902 4196
rect 12919 4132 12983 4196
rect 13000 4132 13064 4196
rect 13081 4132 13145 4196
rect 13162 4132 13226 4196
rect 13243 4132 13307 4196
rect 13324 4132 13388 4196
rect 13405 4132 13469 4196
rect 13486 4132 13550 4196
rect 13567 4132 13631 4196
rect 13648 4132 13712 4196
rect 13729 4132 13793 4196
rect 13810 4132 13874 4196
rect 13891 4132 13955 4196
rect 13972 4132 14036 4196
rect 14053 4132 14117 4196
rect 14134 4132 14198 4196
rect 14215 4132 14279 4196
rect 14296 4132 14360 4196
rect 14378 4132 14442 4196
rect 14460 4132 14524 4196
rect 14542 4132 14606 4196
rect 14624 4132 14688 4196
rect 14706 4132 14770 4196
rect 14788 4132 14852 4196
rect 10084 4046 10148 4110
rect 10165 4046 10229 4110
rect 10246 4046 10310 4110
rect 10327 4046 10391 4110
rect 10408 4046 10472 4110
rect 10489 4046 10553 4110
rect 10570 4046 10634 4110
rect 10651 4046 10715 4110
rect 10732 4046 10796 4110
rect 10813 4046 10877 4110
rect 10894 4046 10958 4110
rect 10975 4046 11039 4110
rect 11056 4046 11120 4110
rect 11137 4046 11201 4110
rect 11218 4046 11282 4110
rect 11299 4046 11363 4110
rect 11380 4046 11444 4110
rect 11461 4046 11525 4110
rect 11542 4046 11606 4110
rect 11623 4046 11687 4110
rect 11704 4046 11768 4110
rect 11785 4046 11849 4110
rect 11866 4046 11930 4110
rect 11947 4046 12011 4110
rect 12028 4046 12092 4110
rect 12109 4046 12173 4110
rect 12190 4046 12254 4110
rect 12271 4046 12335 4110
rect 12352 4046 12416 4110
rect 12433 4046 12497 4110
rect 12514 4046 12578 4110
rect 12595 4046 12659 4110
rect 12676 4046 12740 4110
rect 12757 4046 12821 4110
rect 12838 4046 12902 4110
rect 12919 4046 12983 4110
rect 13000 4046 13064 4110
rect 13081 4046 13145 4110
rect 13162 4046 13226 4110
rect 13243 4046 13307 4110
rect 13324 4046 13388 4110
rect 13405 4046 13469 4110
rect 13486 4046 13550 4110
rect 13567 4046 13631 4110
rect 13648 4046 13712 4110
rect 13729 4046 13793 4110
rect 13810 4046 13874 4110
rect 13891 4046 13955 4110
rect 13972 4046 14036 4110
rect 14053 4046 14117 4110
rect 14134 4046 14198 4110
rect 14215 4046 14279 4110
rect 14296 4046 14360 4110
rect 14378 4046 14442 4110
rect 14460 4046 14524 4110
rect 14542 4046 14606 4110
rect 14624 4046 14688 4110
rect 14706 4046 14770 4110
rect 14788 4046 14852 4110
rect 10084 3960 10148 4024
rect 10165 3960 10229 4024
rect 10246 3960 10310 4024
rect 10327 3960 10391 4024
rect 10408 3960 10472 4024
rect 10489 3960 10553 4024
rect 10570 3960 10634 4024
rect 10651 3960 10715 4024
rect 10732 3960 10796 4024
rect 10813 3960 10877 4024
rect 10894 3960 10958 4024
rect 10975 3960 11039 4024
rect 11056 3960 11120 4024
rect 11137 3960 11201 4024
rect 11218 3960 11282 4024
rect 11299 3960 11363 4024
rect 11380 3960 11444 4024
rect 11461 3960 11525 4024
rect 11542 3960 11606 4024
rect 11623 3960 11687 4024
rect 11704 3960 11768 4024
rect 11785 3960 11849 4024
rect 11866 3960 11930 4024
rect 11947 3960 12011 4024
rect 12028 3960 12092 4024
rect 12109 3960 12173 4024
rect 12190 3960 12254 4024
rect 12271 3960 12335 4024
rect 12352 3960 12416 4024
rect 12433 3960 12497 4024
rect 12514 3960 12578 4024
rect 12595 3960 12659 4024
rect 12676 3960 12740 4024
rect 12757 3960 12821 4024
rect 12838 3960 12902 4024
rect 12919 3960 12983 4024
rect 13000 3960 13064 4024
rect 13081 3960 13145 4024
rect 13162 3960 13226 4024
rect 13243 3960 13307 4024
rect 13324 3960 13388 4024
rect 13405 3960 13469 4024
rect 13486 3960 13550 4024
rect 13567 3960 13631 4024
rect 13648 3960 13712 4024
rect 13729 3960 13793 4024
rect 13810 3960 13874 4024
rect 13891 3960 13955 4024
rect 13972 3960 14036 4024
rect 14053 3960 14117 4024
rect 14134 3960 14198 4024
rect 14215 3960 14279 4024
rect 14296 3960 14360 4024
rect 14378 3960 14442 4024
rect 14460 3960 14524 4024
rect 14542 3960 14606 4024
rect 14624 3960 14688 4024
rect 14706 3960 14770 4024
rect 14788 3960 14852 4024
<< metal4 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 18954 254 19000
rect 14746 18954 15000 19000
rect 0 18950 3948 18954
rect 0 18886 162 18950
rect 226 18886 243 18950
rect 307 18886 324 18950
rect 388 18886 405 18950
rect 469 18886 486 18950
rect 550 18886 567 18950
rect 631 18886 648 18950
rect 712 18886 729 18950
rect 793 18886 810 18950
rect 874 18886 891 18950
rect 955 18886 972 18950
rect 1036 18886 1053 18950
rect 1117 18886 1134 18950
rect 1198 18886 1215 18950
rect 1279 18886 1296 18950
rect 1360 18886 1377 18950
rect 1441 18886 1458 18950
rect 1522 18886 1539 18950
rect 1603 18886 1620 18950
rect 1684 18886 1701 18950
rect 1765 18886 1782 18950
rect 1846 18886 1863 18950
rect 1927 18886 1944 18950
rect 2008 18886 2025 18950
rect 2089 18886 2106 18950
rect 2170 18886 2187 18950
rect 2251 18886 2268 18950
rect 2332 18886 2349 18950
rect 2413 18886 2430 18950
rect 2494 18886 2511 18950
rect 2575 18886 2592 18950
rect 2656 18886 2673 18950
rect 2737 18886 2754 18950
rect 2818 18886 2835 18950
rect 2899 18886 2916 18950
rect 2980 18886 2997 18950
rect 3061 18886 3078 18950
rect 3142 18886 3159 18950
rect 3223 18886 3240 18950
rect 3304 18886 3321 18950
rect 3385 18886 3402 18950
rect 3466 18886 3483 18950
rect 3547 18886 3563 18950
rect 3627 18886 3643 18950
rect 3707 18886 3723 18950
rect 3787 18886 3803 18950
rect 3867 18886 3883 18950
rect 3947 18886 3948 18950
rect 0 18866 3948 18886
rect 0 18802 162 18866
rect 226 18802 243 18866
rect 307 18802 324 18866
rect 388 18802 405 18866
rect 469 18802 486 18866
rect 550 18802 567 18866
rect 631 18802 648 18866
rect 712 18802 729 18866
rect 793 18802 810 18866
rect 874 18802 891 18866
rect 955 18802 972 18866
rect 1036 18802 1053 18866
rect 1117 18802 1134 18866
rect 1198 18802 1215 18866
rect 1279 18802 1296 18866
rect 1360 18802 1377 18866
rect 1441 18802 1458 18866
rect 1522 18802 1539 18866
rect 1603 18802 1620 18866
rect 1684 18802 1701 18866
rect 1765 18802 1782 18866
rect 1846 18802 1863 18866
rect 1927 18802 1944 18866
rect 2008 18802 2025 18866
rect 2089 18802 2106 18866
rect 2170 18802 2187 18866
rect 2251 18802 2268 18866
rect 2332 18802 2349 18866
rect 2413 18802 2430 18866
rect 2494 18802 2511 18866
rect 2575 18802 2592 18866
rect 2656 18802 2673 18866
rect 2737 18802 2754 18866
rect 2818 18802 2835 18866
rect 2899 18802 2916 18866
rect 2980 18802 2997 18866
rect 3061 18802 3078 18866
rect 3142 18802 3159 18866
rect 3223 18802 3240 18866
rect 3304 18802 3321 18866
rect 3385 18802 3402 18866
rect 3466 18802 3483 18866
rect 3547 18802 3563 18866
rect 3627 18802 3643 18866
rect 3707 18802 3723 18866
rect 3787 18802 3803 18866
rect 3867 18802 3883 18866
rect 3947 18802 3948 18866
rect 0 18782 3948 18802
rect 0 18718 162 18782
rect 226 18718 243 18782
rect 307 18718 324 18782
rect 388 18718 405 18782
rect 469 18718 486 18782
rect 550 18718 567 18782
rect 631 18718 648 18782
rect 712 18718 729 18782
rect 793 18718 810 18782
rect 874 18718 891 18782
rect 955 18718 972 18782
rect 1036 18718 1053 18782
rect 1117 18718 1134 18782
rect 1198 18718 1215 18782
rect 1279 18718 1296 18782
rect 1360 18718 1377 18782
rect 1441 18718 1458 18782
rect 1522 18718 1539 18782
rect 1603 18718 1620 18782
rect 1684 18718 1701 18782
rect 1765 18718 1782 18782
rect 1846 18718 1863 18782
rect 1927 18718 1944 18782
rect 2008 18718 2025 18782
rect 2089 18718 2106 18782
rect 2170 18718 2187 18782
rect 2251 18718 2268 18782
rect 2332 18718 2349 18782
rect 2413 18718 2430 18782
rect 2494 18718 2511 18782
rect 2575 18718 2592 18782
rect 2656 18718 2673 18782
rect 2737 18718 2754 18782
rect 2818 18718 2835 18782
rect 2899 18718 2916 18782
rect 2980 18718 2997 18782
rect 3061 18718 3078 18782
rect 3142 18718 3159 18782
rect 3223 18718 3240 18782
rect 3304 18718 3321 18782
rect 3385 18718 3402 18782
rect 3466 18718 3483 18782
rect 3547 18718 3563 18782
rect 3627 18718 3643 18782
rect 3707 18718 3723 18782
rect 3787 18718 3803 18782
rect 3867 18718 3883 18782
rect 3947 18718 3948 18782
rect 11064 18950 15000 18954
rect 11064 18886 11065 18950
rect 11129 18886 11145 18950
rect 11209 18886 11225 18950
rect 11289 18886 11305 18950
rect 11369 18886 11385 18950
rect 11449 18886 11465 18950
rect 11529 18886 11546 18950
rect 11610 18886 11627 18950
rect 11691 18886 11708 18950
rect 11772 18886 11789 18950
rect 11853 18886 11870 18950
rect 11934 18886 11951 18950
rect 12015 18886 12032 18950
rect 12096 18886 12113 18950
rect 12177 18886 12194 18950
rect 12258 18886 12275 18950
rect 12339 18886 12356 18950
rect 12420 18886 12437 18950
rect 12501 18886 12518 18950
rect 12582 18886 12599 18950
rect 12663 18886 12680 18950
rect 12744 18886 12761 18950
rect 12825 18886 12842 18950
rect 12906 18886 12923 18950
rect 12987 18886 13004 18950
rect 13068 18886 13085 18950
rect 13149 18886 13166 18950
rect 13230 18886 13247 18950
rect 13311 18886 13328 18950
rect 13392 18886 13409 18950
rect 13473 18886 13490 18950
rect 13554 18886 13571 18950
rect 13635 18886 13652 18950
rect 13716 18886 13733 18950
rect 13797 18886 13814 18950
rect 13878 18886 13895 18950
rect 13959 18886 13976 18950
rect 14040 18886 14057 18950
rect 14121 18886 14138 18950
rect 14202 18886 14219 18950
rect 14283 18886 14300 18950
rect 14364 18886 14381 18950
rect 14445 18886 14462 18950
rect 14526 18886 14543 18950
rect 14607 18886 14624 18950
rect 14688 18886 14705 18950
rect 14769 18886 14786 18950
rect 14850 18886 15000 18950
rect 11064 18866 15000 18886
rect 11064 18802 11065 18866
rect 11129 18802 11145 18866
rect 11209 18802 11225 18866
rect 11289 18802 11305 18866
rect 11369 18802 11385 18866
rect 11449 18802 11465 18866
rect 11529 18802 11546 18866
rect 11610 18802 11627 18866
rect 11691 18802 11708 18866
rect 11772 18802 11789 18866
rect 11853 18802 11870 18866
rect 11934 18802 11951 18866
rect 12015 18802 12032 18866
rect 12096 18802 12113 18866
rect 12177 18802 12194 18866
rect 12258 18802 12275 18866
rect 12339 18802 12356 18866
rect 12420 18802 12437 18866
rect 12501 18802 12518 18866
rect 12582 18802 12599 18866
rect 12663 18802 12680 18866
rect 12744 18802 12761 18866
rect 12825 18802 12842 18866
rect 12906 18802 12923 18866
rect 12987 18802 13004 18866
rect 13068 18802 13085 18866
rect 13149 18802 13166 18866
rect 13230 18802 13247 18866
rect 13311 18802 13328 18866
rect 13392 18802 13409 18866
rect 13473 18802 13490 18866
rect 13554 18802 13571 18866
rect 13635 18802 13652 18866
rect 13716 18802 13733 18866
rect 13797 18802 13814 18866
rect 13878 18802 13895 18866
rect 13959 18802 13976 18866
rect 14040 18802 14057 18866
rect 14121 18802 14138 18866
rect 14202 18802 14219 18866
rect 14283 18802 14300 18866
rect 14364 18802 14381 18866
rect 14445 18802 14462 18866
rect 14526 18802 14543 18866
rect 14607 18802 14624 18866
rect 14688 18802 14705 18866
rect 14769 18802 14786 18866
rect 14850 18802 15000 18866
rect 11064 18782 15000 18802
rect 0 18698 3948 18718
rect 0 18634 162 18698
rect 226 18634 243 18698
rect 307 18634 324 18698
rect 388 18634 405 18698
rect 469 18634 486 18698
rect 550 18634 567 18698
rect 631 18634 648 18698
rect 712 18634 729 18698
rect 793 18634 810 18698
rect 874 18634 891 18698
rect 955 18634 972 18698
rect 1036 18634 1053 18698
rect 1117 18634 1134 18698
rect 1198 18634 1215 18698
rect 1279 18634 1296 18698
rect 1360 18634 1377 18698
rect 1441 18634 1458 18698
rect 1522 18634 1539 18698
rect 1603 18634 1620 18698
rect 1684 18634 1701 18698
rect 1765 18634 1782 18698
rect 1846 18634 1863 18698
rect 1927 18634 1944 18698
rect 2008 18634 2025 18698
rect 2089 18634 2106 18698
rect 2170 18634 2187 18698
rect 2251 18634 2268 18698
rect 2332 18634 2349 18698
rect 2413 18634 2430 18698
rect 2494 18634 2511 18698
rect 2575 18634 2592 18698
rect 2656 18634 2673 18698
rect 2737 18634 2754 18698
rect 2818 18634 2835 18698
rect 2899 18634 2916 18698
rect 2980 18634 2997 18698
rect 3061 18634 3078 18698
rect 3142 18634 3159 18698
rect 3223 18634 3240 18698
rect 3304 18634 3321 18698
rect 3385 18634 3402 18698
rect 3466 18634 3483 18698
rect 3547 18634 3563 18698
rect 3627 18634 3643 18698
rect 3707 18634 3723 18698
rect 3787 18634 3803 18698
rect 3867 18634 3883 18698
rect 3947 18634 3948 18698
rect 0 18614 3948 18634
rect 0 18550 162 18614
rect 226 18550 243 18614
rect 307 18550 324 18614
rect 388 18550 405 18614
rect 469 18550 486 18614
rect 550 18550 567 18614
rect 631 18550 648 18614
rect 712 18550 729 18614
rect 793 18550 810 18614
rect 874 18550 891 18614
rect 955 18550 972 18614
rect 1036 18550 1053 18614
rect 1117 18550 1134 18614
rect 1198 18550 1215 18614
rect 1279 18550 1296 18614
rect 1360 18550 1377 18614
rect 1441 18550 1458 18614
rect 1522 18550 1539 18614
rect 1603 18550 1620 18614
rect 1684 18550 1701 18614
rect 1765 18550 1782 18614
rect 1846 18550 1863 18614
rect 1927 18550 1944 18614
rect 2008 18550 2025 18614
rect 2089 18550 2106 18614
rect 2170 18550 2187 18614
rect 2251 18550 2268 18614
rect 2332 18550 2349 18614
rect 2413 18550 2430 18614
rect 2494 18550 2511 18614
rect 2575 18550 2592 18614
rect 2656 18550 2673 18614
rect 2737 18550 2754 18614
rect 2818 18550 2835 18614
rect 2899 18550 2916 18614
rect 2980 18550 2997 18614
rect 3061 18550 3078 18614
rect 3142 18550 3159 18614
rect 3223 18550 3240 18614
rect 3304 18550 3321 18614
rect 3385 18550 3402 18614
rect 3466 18550 3483 18614
rect 3547 18550 3563 18614
rect 3627 18550 3643 18614
rect 3707 18550 3723 18614
rect 3787 18550 3803 18614
rect 3867 18550 3883 18614
rect 3947 18550 3948 18614
rect 3993 18765 4189 18766
rect 3993 18701 3994 18765
rect 4058 18701 4124 18765
rect 4188 18701 4189 18765
rect 3993 18643 4189 18701
rect 3993 18579 3994 18643
rect 4058 18579 4124 18643
rect 4188 18579 4189 18643
rect 3993 18578 4189 18579
rect 10823 18765 11019 18766
rect 10823 18701 10824 18765
rect 10888 18701 10954 18765
rect 11018 18701 11019 18765
rect 10823 18643 11019 18701
rect 10823 18579 10824 18643
rect 10888 18579 10954 18643
rect 11018 18579 11019 18643
rect 10823 18578 11019 18579
rect 11064 18718 11065 18782
rect 11129 18718 11145 18782
rect 11209 18718 11225 18782
rect 11289 18718 11305 18782
rect 11369 18718 11385 18782
rect 11449 18718 11465 18782
rect 11529 18718 11546 18782
rect 11610 18718 11627 18782
rect 11691 18718 11708 18782
rect 11772 18718 11789 18782
rect 11853 18718 11870 18782
rect 11934 18718 11951 18782
rect 12015 18718 12032 18782
rect 12096 18718 12113 18782
rect 12177 18718 12194 18782
rect 12258 18718 12275 18782
rect 12339 18718 12356 18782
rect 12420 18718 12437 18782
rect 12501 18718 12518 18782
rect 12582 18718 12599 18782
rect 12663 18718 12680 18782
rect 12744 18718 12761 18782
rect 12825 18718 12842 18782
rect 12906 18718 12923 18782
rect 12987 18718 13004 18782
rect 13068 18718 13085 18782
rect 13149 18718 13166 18782
rect 13230 18718 13247 18782
rect 13311 18718 13328 18782
rect 13392 18718 13409 18782
rect 13473 18718 13490 18782
rect 13554 18718 13571 18782
rect 13635 18718 13652 18782
rect 13716 18718 13733 18782
rect 13797 18718 13814 18782
rect 13878 18718 13895 18782
rect 13959 18718 13976 18782
rect 14040 18718 14057 18782
rect 14121 18718 14138 18782
rect 14202 18718 14219 18782
rect 14283 18718 14300 18782
rect 14364 18718 14381 18782
rect 14445 18718 14462 18782
rect 14526 18718 14543 18782
rect 14607 18718 14624 18782
rect 14688 18718 14705 18782
rect 14769 18718 14786 18782
rect 14850 18718 15000 18782
rect 11064 18698 15000 18718
rect 11064 18634 11065 18698
rect 11129 18634 11145 18698
rect 11209 18634 11225 18698
rect 11289 18634 11305 18698
rect 11369 18634 11385 18698
rect 11449 18634 11465 18698
rect 11529 18634 11546 18698
rect 11610 18634 11627 18698
rect 11691 18634 11708 18698
rect 11772 18634 11789 18698
rect 11853 18634 11870 18698
rect 11934 18634 11951 18698
rect 12015 18634 12032 18698
rect 12096 18634 12113 18698
rect 12177 18634 12194 18698
rect 12258 18634 12275 18698
rect 12339 18634 12356 18698
rect 12420 18634 12437 18698
rect 12501 18634 12518 18698
rect 12582 18634 12599 18698
rect 12663 18634 12680 18698
rect 12744 18634 12761 18698
rect 12825 18634 12842 18698
rect 12906 18634 12923 18698
rect 12987 18634 13004 18698
rect 13068 18634 13085 18698
rect 13149 18634 13166 18698
rect 13230 18634 13247 18698
rect 13311 18634 13328 18698
rect 13392 18634 13409 18698
rect 13473 18634 13490 18698
rect 13554 18634 13571 18698
rect 13635 18634 13652 18698
rect 13716 18634 13733 18698
rect 13797 18634 13814 18698
rect 13878 18634 13895 18698
rect 13959 18634 13976 18698
rect 14040 18634 14057 18698
rect 14121 18634 14138 18698
rect 14202 18634 14219 18698
rect 14283 18634 14300 18698
rect 14364 18634 14381 18698
rect 14445 18634 14462 18698
rect 14526 18634 14543 18698
rect 14607 18634 14624 18698
rect 14688 18634 14705 18698
rect 14769 18634 14786 18698
rect 14850 18634 15000 18698
rect 11064 18614 15000 18634
rect 0 18530 3948 18550
rect 0 18466 162 18530
rect 226 18466 243 18530
rect 307 18466 324 18530
rect 388 18466 405 18530
rect 469 18466 486 18530
rect 550 18466 567 18530
rect 631 18466 648 18530
rect 712 18466 729 18530
rect 793 18466 810 18530
rect 874 18466 891 18530
rect 955 18466 972 18530
rect 1036 18466 1053 18530
rect 1117 18466 1134 18530
rect 1198 18466 1215 18530
rect 1279 18466 1296 18530
rect 1360 18466 1377 18530
rect 1441 18466 1458 18530
rect 1522 18466 1539 18530
rect 1603 18466 1620 18530
rect 1684 18466 1701 18530
rect 1765 18466 1782 18530
rect 1846 18466 1863 18530
rect 1927 18466 1944 18530
rect 2008 18466 2025 18530
rect 2089 18466 2106 18530
rect 2170 18466 2187 18530
rect 2251 18466 2268 18530
rect 2332 18466 2349 18530
rect 2413 18466 2430 18530
rect 2494 18466 2511 18530
rect 2575 18466 2592 18530
rect 2656 18466 2673 18530
rect 2737 18466 2754 18530
rect 2818 18466 2835 18530
rect 2899 18466 2916 18530
rect 2980 18466 2997 18530
rect 3061 18466 3078 18530
rect 3142 18466 3159 18530
rect 3223 18466 3240 18530
rect 3304 18466 3321 18530
rect 3385 18466 3402 18530
rect 3466 18466 3483 18530
rect 3547 18466 3563 18530
rect 3627 18466 3643 18530
rect 3707 18466 3723 18530
rect 3787 18466 3803 18530
rect 3867 18466 3883 18530
rect 3947 18466 3948 18530
rect 11064 18550 11065 18614
rect 11129 18550 11145 18614
rect 11209 18550 11225 18614
rect 11289 18550 11305 18614
rect 11369 18550 11385 18614
rect 11449 18550 11465 18614
rect 11529 18550 11546 18614
rect 11610 18550 11627 18614
rect 11691 18550 11708 18614
rect 11772 18550 11789 18614
rect 11853 18550 11870 18614
rect 11934 18550 11951 18614
rect 12015 18550 12032 18614
rect 12096 18550 12113 18614
rect 12177 18550 12194 18614
rect 12258 18550 12275 18614
rect 12339 18550 12356 18614
rect 12420 18550 12437 18614
rect 12501 18550 12518 18614
rect 12582 18550 12599 18614
rect 12663 18550 12680 18614
rect 12744 18550 12761 18614
rect 12825 18550 12842 18614
rect 12906 18550 12923 18614
rect 12987 18550 13004 18614
rect 13068 18550 13085 18614
rect 13149 18550 13166 18614
rect 13230 18550 13247 18614
rect 13311 18550 13328 18614
rect 13392 18550 13409 18614
rect 13473 18550 13490 18614
rect 13554 18550 13571 18614
rect 13635 18550 13652 18614
rect 13716 18550 13733 18614
rect 13797 18550 13814 18614
rect 13878 18550 13895 18614
rect 13959 18550 13976 18614
rect 14040 18550 14057 18614
rect 14121 18550 14138 18614
rect 14202 18550 14219 18614
rect 14283 18550 14300 18614
rect 14364 18550 14381 18614
rect 14445 18550 14462 18614
rect 14526 18550 14543 18614
rect 14607 18550 14624 18614
rect 14688 18550 14705 18614
rect 14769 18550 14786 18614
rect 14850 18550 15000 18614
rect 11064 18530 15000 18550
rect 0 18446 3948 18466
rect 0 18382 162 18446
rect 226 18382 243 18446
rect 307 18382 324 18446
rect 388 18382 405 18446
rect 469 18382 486 18446
rect 550 18382 567 18446
rect 631 18382 648 18446
rect 712 18382 729 18446
rect 793 18382 810 18446
rect 874 18382 891 18446
rect 955 18382 972 18446
rect 1036 18382 1053 18446
rect 1117 18382 1134 18446
rect 1198 18382 1215 18446
rect 1279 18382 1296 18446
rect 1360 18382 1377 18446
rect 1441 18382 1458 18446
rect 1522 18382 1539 18446
rect 1603 18382 1620 18446
rect 1684 18382 1701 18446
rect 1765 18382 1782 18446
rect 1846 18382 1863 18446
rect 1927 18382 1944 18446
rect 2008 18382 2025 18446
rect 2089 18382 2106 18446
rect 2170 18382 2187 18446
rect 2251 18382 2268 18446
rect 2332 18382 2349 18446
rect 2413 18382 2430 18446
rect 2494 18382 2511 18446
rect 2575 18382 2592 18446
rect 2656 18382 2673 18446
rect 2737 18382 2754 18446
rect 2818 18382 2835 18446
rect 2899 18382 2916 18446
rect 2980 18382 2997 18446
rect 3061 18382 3078 18446
rect 3142 18382 3159 18446
rect 3223 18382 3240 18446
rect 3304 18382 3321 18446
rect 3385 18382 3402 18446
rect 3466 18382 3483 18446
rect 3547 18382 3563 18446
rect 3627 18382 3643 18446
rect 3707 18382 3723 18446
rect 3787 18382 3803 18446
rect 3867 18382 3883 18446
rect 3947 18382 3948 18446
rect 0 18362 3948 18382
rect 0 18298 162 18362
rect 226 18298 243 18362
rect 307 18298 324 18362
rect 388 18298 405 18362
rect 469 18298 486 18362
rect 550 18298 567 18362
rect 631 18298 648 18362
rect 712 18298 729 18362
rect 793 18298 810 18362
rect 874 18298 891 18362
rect 955 18298 972 18362
rect 1036 18298 1053 18362
rect 1117 18298 1134 18362
rect 1198 18298 1215 18362
rect 1279 18298 1296 18362
rect 1360 18298 1377 18362
rect 1441 18298 1458 18362
rect 1522 18298 1539 18362
rect 1603 18298 1620 18362
rect 1684 18298 1701 18362
rect 1765 18298 1782 18362
rect 1846 18298 1863 18362
rect 1927 18298 1944 18362
rect 2008 18298 2025 18362
rect 2089 18298 2106 18362
rect 2170 18298 2187 18362
rect 2251 18298 2268 18362
rect 2332 18298 2349 18362
rect 2413 18298 2430 18362
rect 2494 18298 2511 18362
rect 2575 18298 2592 18362
rect 2656 18298 2673 18362
rect 2737 18298 2754 18362
rect 2818 18298 2835 18362
rect 2899 18298 2916 18362
rect 2980 18298 2997 18362
rect 3061 18298 3078 18362
rect 3142 18298 3159 18362
rect 3223 18298 3240 18362
rect 3304 18298 3321 18362
rect 3385 18298 3402 18362
rect 3466 18298 3483 18362
rect 3547 18298 3563 18362
rect 3627 18298 3643 18362
rect 3707 18298 3723 18362
rect 3787 18298 3803 18362
rect 3867 18298 3883 18362
rect 3947 18298 3948 18362
rect 0 18278 3948 18298
rect 0 18214 162 18278
rect 226 18214 243 18278
rect 307 18214 324 18278
rect 388 18214 405 18278
rect 469 18214 486 18278
rect 550 18214 567 18278
rect 631 18214 648 18278
rect 712 18214 729 18278
rect 793 18214 810 18278
rect 874 18214 891 18278
rect 955 18214 972 18278
rect 1036 18214 1053 18278
rect 1117 18214 1134 18278
rect 1198 18214 1215 18278
rect 1279 18214 1296 18278
rect 1360 18214 1377 18278
rect 1441 18214 1458 18278
rect 1522 18214 1539 18278
rect 1603 18214 1620 18278
rect 1684 18214 1701 18278
rect 1765 18214 1782 18278
rect 1846 18214 1863 18278
rect 1927 18214 1944 18278
rect 2008 18214 2025 18278
rect 2089 18214 2106 18278
rect 2170 18214 2187 18278
rect 2251 18214 2268 18278
rect 2332 18214 2349 18278
rect 2413 18214 2430 18278
rect 2494 18214 2511 18278
rect 2575 18214 2592 18278
rect 2656 18214 2673 18278
rect 2737 18214 2754 18278
rect 2818 18214 2835 18278
rect 2899 18214 2916 18278
rect 2980 18214 2997 18278
rect 3061 18214 3078 18278
rect 3142 18214 3159 18278
rect 3223 18214 3240 18278
rect 3304 18214 3321 18278
rect 3385 18214 3402 18278
rect 3466 18214 3483 18278
rect 3547 18214 3563 18278
rect 3627 18214 3643 18278
rect 3707 18214 3723 18278
rect 3787 18214 3803 18278
rect 3867 18214 3883 18278
rect 3947 18214 3948 18278
rect 0 18194 3948 18214
rect 0 18130 162 18194
rect 226 18130 243 18194
rect 307 18130 324 18194
rect 388 18130 405 18194
rect 469 18130 486 18194
rect 550 18130 567 18194
rect 631 18130 648 18194
rect 712 18130 729 18194
rect 793 18130 810 18194
rect 874 18130 891 18194
rect 955 18130 972 18194
rect 1036 18130 1053 18194
rect 1117 18130 1134 18194
rect 1198 18130 1215 18194
rect 1279 18130 1296 18194
rect 1360 18130 1377 18194
rect 1441 18130 1458 18194
rect 1522 18130 1539 18194
rect 1603 18130 1620 18194
rect 1684 18130 1701 18194
rect 1765 18130 1782 18194
rect 1846 18130 1863 18194
rect 1927 18130 1944 18194
rect 2008 18130 2025 18194
rect 2089 18130 2106 18194
rect 2170 18130 2187 18194
rect 2251 18130 2268 18194
rect 2332 18130 2349 18194
rect 2413 18130 2430 18194
rect 2494 18130 2511 18194
rect 2575 18130 2592 18194
rect 2656 18130 2673 18194
rect 2737 18130 2754 18194
rect 2818 18130 2835 18194
rect 2899 18130 2916 18194
rect 2980 18130 2997 18194
rect 3061 18130 3078 18194
rect 3142 18130 3159 18194
rect 3223 18130 3240 18194
rect 3304 18130 3321 18194
rect 3385 18130 3402 18194
rect 3466 18130 3483 18194
rect 3547 18130 3563 18194
rect 3627 18130 3643 18194
rect 3707 18130 3723 18194
rect 3787 18130 3803 18194
rect 3867 18130 3883 18194
rect 3947 18130 3948 18194
rect 4015 18512 4420 18515
rect 4015 18448 4016 18512
rect 4080 18448 4129 18512
rect 4193 18448 4242 18512
rect 4306 18448 4355 18512
rect 4419 18448 4420 18512
rect 4015 18410 4420 18448
rect 4015 18346 4016 18410
rect 4080 18346 4129 18410
rect 4193 18346 4242 18410
rect 4306 18346 4355 18410
rect 4419 18346 4420 18410
rect 4015 18308 4420 18346
rect 4015 18244 4016 18308
rect 4080 18244 4129 18308
rect 4193 18244 4242 18308
rect 4306 18244 4355 18308
rect 4419 18244 4420 18308
rect 10592 18512 10997 18515
rect 10592 18448 10593 18512
rect 10657 18448 10706 18512
rect 10770 18448 10819 18512
rect 10883 18448 10932 18512
rect 10996 18448 10997 18512
rect 10592 18410 10997 18448
rect 10592 18346 10593 18410
rect 10657 18346 10706 18410
rect 10770 18346 10819 18410
rect 10883 18346 10932 18410
rect 10996 18346 10997 18410
rect 10592 18308 10997 18346
rect 4015 18206 4420 18244
rect 4015 18142 4016 18206
rect 4080 18142 4129 18206
rect 4193 18142 4242 18206
rect 4306 18142 4355 18206
rect 4419 18142 4420 18206
rect 4015 18139 4420 18142
rect 4477 18297 4663 18298
rect 4477 18233 4478 18297
rect 4542 18233 4598 18297
rect 4662 18233 4663 18297
rect 4477 18183 4663 18233
rect 0 18126 3948 18130
rect 0 18087 254 18126
rect 4477 18119 4478 18183
rect 4542 18119 4598 18183
rect 4662 18119 4663 18183
rect 4477 18118 4663 18119
rect 10349 18297 10535 18298
rect 10349 18233 10350 18297
rect 10414 18233 10470 18297
rect 10534 18233 10535 18297
rect 10349 18183 10535 18233
rect 10349 18119 10350 18183
rect 10414 18119 10470 18183
rect 10534 18119 10535 18183
rect 10592 18244 10593 18308
rect 10657 18244 10706 18308
rect 10770 18244 10819 18308
rect 10883 18244 10932 18308
rect 10996 18244 10997 18308
rect 10592 18206 10997 18244
rect 10592 18142 10593 18206
rect 10657 18142 10706 18206
rect 10770 18142 10819 18206
rect 10883 18142 10932 18206
rect 10996 18142 10997 18206
rect 10592 18139 10997 18142
rect 11064 18466 11065 18530
rect 11129 18466 11145 18530
rect 11209 18466 11225 18530
rect 11289 18466 11305 18530
rect 11369 18466 11385 18530
rect 11449 18466 11465 18530
rect 11529 18466 11546 18530
rect 11610 18466 11627 18530
rect 11691 18466 11708 18530
rect 11772 18466 11789 18530
rect 11853 18466 11870 18530
rect 11934 18466 11951 18530
rect 12015 18466 12032 18530
rect 12096 18466 12113 18530
rect 12177 18466 12194 18530
rect 12258 18466 12275 18530
rect 12339 18466 12356 18530
rect 12420 18466 12437 18530
rect 12501 18466 12518 18530
rect 12582 18466 12599 18530
rect 12663 18466 12680 18530
rect 12744 18466 12761 18530
rect 12825 18466 12842 18530
rect 12906 18466 12923 18530
rect 12987 18466 13004 18530
rect 13068 18466 13085 18530
rect 13149 18466 13166 18530
rect 13230 18466 13247 18530
rect 13311 18466 13328 18530
rect 13392 18466 13409 18530
rect 13473 18466 13490 18530
rect 13554 18466 13571 18530
rect 13635 18466 13652 18530
rect 13716 18466 13733 18530
rect 13797 18466 13814 18530
rect 13878 18466 13895 18530
rect 13959 18466 13976 18530
rect 14040 18466 14057 18530
rect 14121 18466 14138 18530
rect 14202 18466 14219 18530
rect 14283 18466 14300 18530
rect 14364 18466 14381 18530
rect 14445 18466 14462 18530
rect 14526 18466 14543 18530
rect 14607 18466 14624 18530
rect 14688 18466 14705 18530
rect 14769 18466 14786 18530
rect 14850 18466 15000 18530
rect 11064 18446 15000 18466
rect 11064 18382 11065 18446
rect 11129 18382 11145 18446
rect 11209 18382 11225 18446
rect 11289 18382 11305 18446
rect 11369 18382 11385 18446
rect 11449 18382 11465 18446
rect 11529 18382 11546 18446
rect 11610 18382 11627 18446
rect 11691 18382 11708 18446
rect 11772 18382 11789 18446
rect 11853 18382 11870 18446
rect 11934 18382 11951 18446
rect 12015 18382 12032 18446
rect 12096 18382 12113 18446
rect 12177 18382 12194 18446
rect 12258 18382 12275 18446
rect 12339 18382 12356 18446
rect 12420 18382 12437 18446
rect 12501 18382 12518 18446
rect 12582 18382 12599 18446
rect 12663 18382 12680 18446
rect 12744 18382 12761 18446
rect 12825 18382 12842 18446
rect 12906 18382 12923 18446
rect 12987 18382 13004 18446
rect 13068 18382 13085 18446
rect 13149 18382 13166 18446
rect 13230 18382 13247 18446
rect 13311 18382 13328 18446
rect 13392 18382 13409 18446
rect 13473 18382 13490 18446
rect 13554 18382 13571 18446
rect 13635 18382 13652 18446
rect 13716 18382 13733 18446
rect 13797 18382 13814 18446
rect 13878 18382 13895 18446
rect 13959 18382 13976 18446
rect 14040 18382 14057 18446
rect 14121 18382 14138 18446
rect 14202 18382 14219 18446
rect 14283 18382 14300 18446
rect 14364 18382 14381 18446
rect 14445 18382 14462 18446
rect 14526 18382 14543 18446
rect 14607 18382 14624 18446
rect 14688 18382 14705 18446
rect 14769 18382 14786 18446
rect 14850 18382 15000 18446
rect 11064 18362 15000 18382
rect 11064 18298 11065 18362
rect 11129 18298 11145 18362
rect 11209 18298 11225 18362
rect 11289 18298 11305 18362
rect 11369 18298 11385 18362
rect 11449 18298 11465 18362
rect 11529 18298 11546 18362
rect 11610 18298 11627 18362
rect 11691 18298 11708 18362
rect 11772 18298 11789 18362
rect 11853 18298 11870 18362
rect 11934 18298 11951 18362
rect 12015 18298 12032 18362
rect 12096 18298 12113 18362
rect 12177 18298 12194 18362
rect 12258 18298 12275 18362
rect 12339 18298 12356 18362
rect 12420 18298 12437 18362
rect 12501 18298 12518 18362
rect 12582 18298 12599 18362
rect 12663 18298 12680 18362
rect 12744 18298 12761 18362
rect 12825 18298 12842 18362
rect 12906 18298 12923 18362
rect 12987 18298 13004 18362
rect 13068 18298 13085 18362
rect 13149 18298 13166 18362
rect 13230 18298 13247 18362
rect 13311 18298 13328 18362
rect 13392 18298 13409 18362
rect 13473 18298 13490 18362
rect 13554 18298 13571 18362
rect 13635 18298 13652 18362
rect 13716 18298 13733 18362
rect 13797 18298 13814 18362
rect 13878 18298 13895 18362
rect 13959 18298 13976 18362
rect 14040 18298 14057 18362
rect 14121 18298 14138 18362
rect 14202 18298 14219 18362
rect 14283 18298 14300 18362
rect 14364 18298 14381 18362
rect 14445 18298 14462 18362
rect 14526 18298 14543 18362
rect 14607 18298 14624 18362
rect 14688 18298 14705 18362
rect 14769 18298 14786 18362
rect 14850 18298 15000 18362
rect 11064 18278 15000 18298
rect 11064 18214 11065 18278
rect 11129 18214 11145 18278
rect 11209 18214 11225 18278
rect 11289 18214 11305 18278
rect 11369 18214 11385 18278
rect 11449 18214 11465 18278
rect 11529 18214 11546 18278
rect 11610 18214 11627 18278
rect 11691 18214 11708 18278
rect 11772 18214 11789 18278
rect 11853 18214 11870 18278
rect 11934 18214 11951 18278
rect 12015 18214 12032 18278
rect 12096 18214 12113 18278
rect 12177 18214 12194 18278
rect 12258 18214 12275 18278
rect 12339 18214 12356 18278
rect 12420 18214 12437 18278
rect 12501 18214 12518 18278
rect 12582 18214 12599 18278
rect 12663 18214 12680 18278
rect 12744 18214 12761 18278
rect 12825 18214 12842 18278
rect 12906 18214 12923 18278
rect 12987 18214 13004 18278
rect 13068 18214 13085 18278
rect 13149 18214 13166 18278
rect 13230 18214 13247 18278
rect 13311 18214 13328 18278
rect 13392 18214 13409 18278
rect 13473 18214 13490 18278
rect 13554 18214 13571 18278
rect 13635 18214 13652 18278
rect 13716 18214 13733 18278
rect 13797 18214 13814 18278
rect 13878 18214 13895 18278
rect 13959 18214 13976 18278
rect 14040 18214 14057 18278
rect 14121 18214 14138 18278
rect 14202 18214 14219 18278
rect 14283 18214 14300 18278
rect 14364 18214 14381 18278
rect 14445 18214 14462 18278
rect 14526 18214 14543 18278
rect 14607 18214 14624 18278
rect 14688 18214 14705 18278
rect 14769 18214 14786 18278
rect 14850 18214 15000 18278
rect 11064 18194 15000 18214
rect 11064 18130 11065 18194
rect 11129 18130 11145 18194
rect 11209 18130 11225 18194
rect 11289 18130 11305 18194
rect 11369 18130 11385 18194
rect 11449 18130 11465 18194
rect 11529 18130 11546 18194
rect 11610 18130 11627 18194
rect 11691 18130 11708 18194
rect 11772 18130 11789 18194
rect 11853 18130 11870 18194
rect 11934 18130 11951 18194
rect 12015 18130 12032 18194
rect 12096 18130 12113 18194
rect 12177 18130 12194 18194
rect 12258 18130 12275 18194
rect 12339 18130 12356 18194
rect 12420 18130 12437 18194
rect 12501 18130 12518 18194
rect 12582 18130 12599 18194
rect 12663 18130 12680 18194
rect 12744 18130 12761 18194
rect 12825 18130 12842 18194
rect 12906 18130 12923 18194
rect 12987 18130 13004 18194
rect 13068 18130 13085 18194
rect 13149 18130 13166 18194
rect 13230 18130 13247 18194
rect 13311 18130 13328 18194
rect 13392 18130 13409 18194
rect 13473 18130 13490 18194
rect 13554 18130 13571 18194
rect 13635 18130 13652 18194
rect 13716 18130 13733 18194
rect 13797 18130 13814 18194
rect 13878 18130 13895 18194
rect 13959 18130 13976 18194
rect 14040 18130 14057 18194
rect 14121 18130 14138 18194
rect 14202 18130 14219 18194
rect 14283 18130 14300 18194
rect 14364 18130 14381 18194
rect 14445 18130 14462 18194
rect 14526 18130 14543 18194
rect 14607 18130 14624 18194
rect 14688 18130 14705 18194
rect 14769 18130 14786 18194
rect 14850 18130 15000 18194
rect 11064 18126 15000 18130
rect 10349 18118 10535 18119
rect 14746 18087 15000 18126
rect 0 18086 4880 18087
rect 0 14742 137 18086
rect 4841 14742 4880 18086
rect 0 14725 4880 14742
rect 0 14661 137 14725
rect 201 14661 217 14725
rect 281 14661 297 14725
rect 361 14661 377 14725
rect 441 14661 457 14725
rect 521 14661 537 14725
rect 601 14661 617 14725
rect 681 14661 697 14725
rect 761 14661 777 14725
rect 841 14661 857 14725
rect 921 14661 937 14725
rect 1001 14661 1017 14725
rect 1081 14661 1097 14725
rect 1161 14661 1177 14725
rect 1241 14661 1257 14725
rect 1321 14661 1337 14725
rect 1401 14661 1417 14725
rect 1481 14661 1497 14725
rect 1561 14661 1577 14725
rect 1641 14661 1657 14725
rect 1721 14661 1737 14725
rect 1801 14661 1817 14725
rect 1881 14661 1897 14725
rect 1961 14661 1977 14725
rect 2041 14661 2057 14725
rect 2121 14661 2137 14725
rect 2201 14661 2217 14725
rect 2281 14661 2297 14725
rect 2361 14661 2377 14725
rect 2441 14661 2457 14725
rect 2521 14661 2537 14725
rect 2601 14661 2617 14725
rect 2681 14661 2697 14725
rect 2761 14661 2777 14725
rect 2841 14661 2857 14725
rect 2921 14661 2937 14725
rect 3001 14661 3017 14725
rect 3081 14661 3097 14725
rect 3161 14661 3177 14725
rect 3241 14661 3257 14725
rect 3321 14661 3337 14725
rect 3401 14661 3417 14725
rect 3481 14661 3497 14725
rect 3561 14661 3577 14725
rect 3641 14661 3657 14725
rect 3721 14661 3737 14725
rect 3801 14661 3817 14725
rect 3881 14661 3897 14725
rect 3961 14661 3977 14725
rect 4041 14661 4057 14725
rect 4121 14661 4137 14725
rect 4201 14661 4217 14725
rect 4281 14661 4297 14725
rect 4361 14661 4377 14725
rect 4441 14661 4457 14725
rect 4521 14661 4537 14725
rect 4601 14661 4617 14725
rect 4681 14661 4697 14725
rect 4761 14661 4777 14725
rect 4841 14661 4880 14725
rect 0 14644 4880 14661
rect 0 14580 137 14644
rect 201 14580 217 14644
rect 281 14580 297 14644
rect 361 14580 377 14644
rect 441 14580 457 14644
rect 521 14580 537 14644
rect 601 14580 617 14644
rect 681 14580 697 14644
rect 761 14580 777 14644
rect 841 14580 857 14644
rect 921 14580 937 14644
rect 1001 14580 1017 14644
rect 1081 14580 1097 14644
rect 1161 14580 1177 14644
rect 1241 14580 1257 14644
rect 1321 14580 1337 14644
rect 1401 14580 1417 14644
rect 1481 14580 1497 14644
rect 1561 14580 1577 14644
rect 1641 14580 1657 14644
rect 1721 14580 1737 14644
rect 1801 14580 1817 14644
rect 1881 14580 1897 14644
rect 1961 14580 1977 14644
rect 2041 14580 2057 14644
rect 2121 14580 2137 14644
rect 2201 14580 2217 14644
rect 2281 14580 2297 14644
rect 2361 14580 2377 14644
rect 2441 14580 2457 14644
rect 2521 14580 2537 14644
rect 2601 14580 2617 14644
rect 2681 14580 2697 14644
rect 2761 14580 2777 14644
rect 2841 14580 2857 14644
rect 2921 14580 2937 14644
rect 3001 14580 3017 14644
rect 3081 14580 3097 14644
rect 3161 14580 3177 14644
rect 3241 14580 3257 14644
rect 3321 14580 3337 14644
rect 3401 14580 3417 14644
rect 3481 14580 3497 14644
rect 3561 14580 3577 14644
rect 3641 14580 3657 14644
rect 3721 14580 3737 14644
rect 3801 14580 3817 14644
rect 3881 14580 3897 14644
rect 3961 14580 3977 14644
rect 4041 14580 4057 14644
rect 4121 14580 4137 14644
rect 4201 14580 4217 14644
rect 4281 14580 4297 14644
rect 4361 14580 4377 14644
rect 4441 14580 4457 14644
rect 4521 14580 4537 14644
rect 4601 14580 4617 14644
rect 4681 14580 4697 14644
rect 4761 14580 4777 14644
rect 4841 14580 4880 14644
rect 0 14563 4880 14580
rect 0 14499 137 14563
rect 201 14499 217 14563
rect 281 14499 297 14563
rect 361 14499 377 14563
rect 441 14499 457 14563
rect 521 14499 537 14563
rect 601 14499 617 14563
rect 681 14499 697 14563
rect 761 14499 777 14563
rect 841 14499 857 14563
rect 921 14499 937 14563
rect 1001 14499 1017 14563
rect 1081 14499 1097 14563
rect 1161 14499 1177 14563
rect 1241 14499 1257 14563
rect 1321 14499 1337 14563
rect 1401 14499 1417 14563
rect 1481 14499 1497 14563
rect 1561 14499 1577 14563
rect 1641 14499 1657 14563
rect 1721 14499 1737 14563
rect 1801 14499 1817 14563
rect 1881 14499 1897 14563
rect 1961 14499 1977 14563
rect 2041 14499 2057 14563
rect 2121 14499 2137 14563
rect 2201 14499 2217 14563
rect 2281 14499 2297 14563
rect 2361 14499 2377 14563
rect 2441 14499 2457 14563
rect 2521 14499 2537 14563
rect 2601 14499 2617 14563
rect 2681 14499 2697 14563
rect 2761 14499 2777 14563
rect 2841 14499 2857 14563
rect 2921 14499 2937 14563
rect 3001 14499 3017 14563
rect 3081 14499 3097 14563
rect 3161 14499 3177 14563
rect 3241 14499 3257 14563
rect 3321 14499 3337 14563
rect 3401 14499 3417 14563
rect 3481 14499 3497 14563
rect 3561 14499 3577 14563
rect 3641 14499 3657 14563
rect 3721 14499 3737 14563
rect 3801 14499 3817 14563
rect 3881 14499 3897 14563
rect 3961 14499 3977 14563
rect 4041 14499 4057 14563
rect 4121 14499 4137 14563
rect 4201 14499 4217 14563
rect 4281 14499 4297 14563
rect 4361 14499 4377 14563
rect 4441 14499 4457 14563
rect 4521 14499 4537 14563
rect 4601 14499 4617 14563
rect 4681 14499 4697 14563
rect 4761 14499 4777 14563
rect 4841 14499 4880 14563
rect 0 14482 4880 14499
rect 0 14418 137 14482
rect 201 14418 217 14482
rect 281 14418 297 14482
rect 361 14418 377 14482
rect 441 14418 457 14482
rect 521 14418 537 14482
rect 601 14418 617 14482
rect 681 14418 697 14482
rect 761 14418 777 14482
rect 841 14418 857 14482
rect 921 14418 937 14482
rect 1001 14418 1017 14482
rect 1081 14418 1097 14482
rect 1161 14418 1177 14482
rect 1241 14418 1257 14482
rect 1321 14418 1337 14482
rect 1401 14418 1417 14482
rect 1481 14418 1497 14482
rect 1561 14418 1577 14482
rect 1641 14418 1657 14482
rect 1721 14418 1737 14482
rect 1801 14418 1817 14482
rect 1881 14418 1897 14482
rect 1961 14418 1977 14482
rect 2041 14418 2057 14482
rect 2121 14418 2137 14482
rect 2201 14418 2217 14482
rect 2281 14418 2297 14482
rect 2361 14418 2377 14482
rect 2441 14418 2457 14482
rect 2521 14418 2537 14482
rect 2601 14418 2617 14482
rect 2681 14418 2697 14482
rect 2761 14418 2777 14482
rect 2841 14418 2857 14482
rect 2921 14418 2937 14482
rect 3001 14418 3017 14482
rect 3081 14418 3097 14482
rect 3161 14418 3177 14482
rect 3241 14418 3257 14482
rect 3321 14418 3337 14482
rect 3401 14418 3417 14482
rect 3481 14418 3497 14482
rect 3561 14418 3577 14482
rect 3641 14418 3657 14482
rect 3721 14418 3737 14482
rect 3801 14418 3817 14482
rect 3881 14418 3897 14482
rect 3961 14418 3977 14482
rect 4041 14418 4057 14482
rect 4121 14418 4137 14482
rect 4201 14418 4217 14482
rect 4281 14418 4297 14482
rect 4361 14418 4377 14482
rect 4441 14418 4457 14482
rect 4521 14418 4537 14482
rect 4601 14418 4617 14482
rect 4681 14418 4697 14482
rect 4761 14418 4777 14482
rect 4841 14418 4880 14482
rect 0 14401 4880 14418
rect 0 14337 137 14401
rect 201 14337 217 14401
rect 281 14337 297 14401
rect 361 14337 377 14401
rect 441 14337 457 14401
rect 521 14337 537 14401
rect 601 14337 617 14401
rect 681 14337 697 14401
rect 761 14337 777 14401
rect 841 14337 857 14401
rect 921 14337 937 14401
rect 1001 14337 1017 14401
rect 1081 14337 1097 14401
rect 1161 14337 1177 14401
rect 1241 14337 1257 14401
rect 1321 14337 1337 14401
rect 1401 14337 1417 14401
rect 1481 14337 1497 14401
rect 1561 14337 1577 14401
rect 1641 14337 1657 14401
rect 1721 14337 1737 14401
rect 1801 14337 1817 14401
rect 1881 14337 1897 14401
rect 1961 14337 1977 14401
rect 2041 14337 2057 14401
rect 2121 14337 2137 14401
rect 2201 14337 2217 14401
rect 2281 14337 2297 14401
rect 2361 14337 2377 14401
rect 2441 14337 2457 14401
rect 2521 14337 2537 14401
rect 2601 14337 2617 14401
rect 2681 14337 2697 14401
rect 2761 14337 2777 14401
rect 2841 14337 2857 14401
rect 2921 14337 2937 14401
rect 3001 14337 3017 14401
rect 3081 14337 3097 14401
rect 3161 14337 3177 14401
rect 3241 14337 3257 14401
rect 3321 14337 3337 14401
rect 3401 14337 3417 14401
rect 3481 14337 3497 14401
rect 3561 14337 3577 14401
rect 3641 14337 3657 14401
rect 3721 14337 3737 14401
rect 3801 14337 3817 14401
rect 3881 14337 3897 14401
rect 3961 14337 3977 14401
rect 4041 14337 4057 14401
rect 4121 14337 4137 14401
rect 4201 14337 4217 14401
rect 4281 14337 4297 14401
rect 4361 14337 4377 14401
rect 4441 14337 4457 14401
rect 4521 14337 4537 14401
rect 4601 14337 4617 14401
rect 4681 14337 4697 14401
rect 4761 14337 4777 14401
rect 4841 14337 4880 14401
rect 0 14320 4880 14337
rect 0 14256 137 14320
rect 201 14256 217 14320
rect 281 14256 297 14320
rect 361 14256 377 14320
rect 441 14256 457 14320
rect 521 14256 537 14320
rect 601 14256 617 14320
rect 681 14256 697 14320
rect 761 14256 777 14320
rect 841 14256 857 14320
rect 921 14256 937 14320
rect 1001 14256 1017 14320
rect 1081 14256 1097 14320
rect 1161 14256 1177 14320
rect 1241 14256 1257 14320
rect 1321 14256 1337 14320
rect 1401 14256 1417 14320
rect 1481 14256 1497 14320
rect 1561 14256 1577 14320
rect 1641 14256 1657 14320
rect 1721 14256 1737 14320
rect 1801 14256 1817 14320
rect 1881 14256 1897 14320
rect 1961 14256 1977 14320
rect 2041 14256 2057 14320
rect 2121 14256 2137 14320
rect 2201 14256 2217 14320
rect 2281 14256 2297 14320
rect 2361 14256 2377 14320
rect 2441 14256 2457 14320
rect 2521 14256 2537 14320
rect 2601 14256 2617 14320
rect 2681 14256 2697 14320
rect 2761 14256 2777 14320
rect 2841 14256 2857 14320
rect 2921 14256 2937 14320
rect 3001 14256 3017 14320
rect 3081 14256 3097 14320
rect 3161 14256 3177 14320
rect 3241 14256 3257 14320
rect 3321 14256 3337 14320
rect 3401 14256 3417 14320
rect 3481 14256 3497 14320
rect 3561 14256 3577 14320
rect 3641 14256 3657 14320
rect 3721 14256 3737 14320
rect 3801 14256 3817 14320
rect 3881 14256 3897 14320
rect 3961 14256 3977 14320
rect 4041 14256 4057 14320
rect 4121 14256 4137 14320
rect 4201 14256 4217 14320
rect 4281 14256 4297 14320
rect 4361 14256 4377 14320
rect 4441 14256 4457 14320
rect 4521 14256 4537 14320
rect 4601 14256 4617 14320
rect 4681 14256 4697 14320
rect 4761 14256 4777 14320
rect 4841 14256 4880 14320
rect 0 14239 4880 14256
rect 0 14175 137 14239
rect 201 14175 217 14239
rect 281 14175 297 14239
rect 361 14175 377 14239
rect 441 14175 457 14239
rect 521 14175 537 14239
rect 601 14175 617 14239
rect 681 14175 697 14239
rect 761 14175 777 14239
rect 841 14175 857 14239
rect 921 14175 937 14239
rect 1001 14175 1017 14239
rect 1081 14175 1097 14239
rect 1161 14175 1177 14239
rect 1241 14175 1257 14239
rect 1321 14175 1337 14239
rect 1401 14175 1417 14239
rect 1481 14175 1497 14239
rect 1561 14175 1577 14239
rect 1641 14175 1657 14239
rect 1721 14175 1737 14239
rect 1801 14175 1817 14239
rect 1881 14175 1897 14239
rect 1961 14175 1977 14239
rect 2041 14175 2057 14239
rect 2121 14175 2137 14239
rect 2201 14175 2217 14239
rect 2281 14175 2297 14239
rect 2361 14175 2377 14239
rect 2441 14175 2457 14239
rect 2521 14175 2537 14239
rect 2601 14175 2617 14239
rect 2681 14175 2697 14239
rect 2761 14175 2777 14239
rect 2841 14175 2857 14239
rect 2921 14175 2937 14239
rect 3001 14175 3017 14239
rect 3081 14175 3097 14239
rect 3161 14175 3177 14239
rect 3241 14175 3257 14239
rect 3321 14175 3337 14239
rect 3401 14175 3417 14239
rect 3481 14175 3497 14239
rect 3561 14175 3577 14239
rect 3641 14175 3657 14239
rect 3721 14175 3737 14239
rect 3801 14175 3817 14239
rect 3881 14175 3897 14239
rect 3961 14175 3977 14239
rect 4041 14175 4057 14239
rect 4121 14175 4137 14239
rect 4201 14175 4217 14239
rect 4281 14175 4297 14239
rect 4361 14175 4377 14239
rect 4441 14175 4457 14239
rect 4521 14175 4537 14239
rect 4601 14175 4617 14239
rect 4681 14175 4697 14239
rect 4761 14175 4777 14239
rect 4841 14175 4880 14239
rect 0 14158 4880 14175
rect 0 14094 137 14158
rect 201 14094 217 14158
rect 281 14094 297 14158
rect 361 14094 377 14158
rect 441 14094 457 14158
rect 521 14094 537 14158
rect 601 14094 617 14158
rect 681 14094 697 14158
rect 761 14094 777 14158
rect 841 14094 857 14158
rect 921 14094 937 14158
rect 1001 14094 1017 14158
rect 1081 14094 1097 14158
rect 1161 14094 1177 14158
rect 1241 14094 1257 14158
rect 1321 14094 1337 14158
rect 1401 14094 1417 14158
rect 1481 14094 1497 14158
rect 1561 14094 1577 14158
rect 1641 14094 1657 14158
rect 1721 14094 1737 14158
rect 1801 14094 1817 14158
rect 1881 14094 1897 14158
rect 1961 14094 1977 14158
rect 2041 14094 2057 14158
rect 2121 14094 2137 14158
rect 2201 14094 2217 14158
rect 2281 14094 2297 14158
rect 2361 14094 2377 14158
rect 2441 14094 2457 14158
rect 2521 14094 2537 14158
rect 2601 14094 2617 14158
rect 2681 14094 2697 14158
rect 2761 14094 2777 14158
rect 2841 14094 2857 14158
rect 2921 14094 2937 14158
rect 3001 14094 3017 14158
rect 3081 14094 3097 14158
rect 3161 14094 3177 14158
rect 3241 14094 3257 14158
rect 3321 14094 3337 14158
rect 3401 14094 3417 14158
rect 3481 14094 3497 14158
rect 3561 14094 3577 14158
rect 3641 14094 3657 14158
rect 3721 14094 3737 14158
rect 3801 14094 3817 14158
rect 3881 14094 3897 14158
rect 3961 14094 3977 14158
rect 4041 14094 4057 14158
rect 4121 14094 4137 14158
rect 4201 14094 4217 14158
rect 4281 14094 4297 14158
rect 4361 14094 4377 14158
rect 4441 14094 4457 14158
rect 4521 14094 4537 14158
rect 4601 14094 4617 14158
rect 4681 14094 4697 14158
rect 4761 14094 4777 14158
rect 4841 14094 4880 14158
rect 0 14077 4880 14094
rect 0 14013 137 14077
rect 201 14013 217 14077
rect 281 14013 297 14077
rect 361 14013 377 14077
rect 441 14013 457 14077
rect 521 14013 537 14077
rect 601 14013 617 14077
rect 681 14013 697 14077
rect 761 14013 777 14077
rect 841 14013 857 14077
rect 921 14013 937 14077
rect 1001 14013 1017 14077
rect 1081 14013 1097 14077
rect 1161 14013 1177 14077
rect 1241 14013 1257 14077
rect 1321 14013 1337 14077
rect 1401 14013 1417 14077
rect 1481 14013 1497 14077
rect 1561 14013 1577 14077
rect 1641 14013 1657 14077
rect 1721 14013 1737 14077
rect 1801 14013 1817 14077
rect 1881 14013 1897 14077
rect 1961 14013 1977 14077
rect 2041 14013 2057 14077
rect 2121 14013 2137 14077
rect 2201 14013 2217 14077
rect 2281 14013 2297 14077
rect 2361 14013 2377 14077
rect 2441 14013 2457 14077
rect 2521 14013 2537 14077
rect 2601 14013 2617 14077
rect 2681 14013 2697 14077
rect 2761 14013 2777 14077
rect 2841 14013 2857 14077
rect 2921 14013 2937 14077
rect 3001 14013 3017 14077
rect 3081 14013 3097 14077
rect 3161 14013 3177 14077
rect 3241 14013 3257 14077
rect 3321 14013 3337 14077
rect 3401 14013 3417 14077
rect 3481 14013 3497 14077
rect 3561 14013 3577 14077
rect 3641 14013 3657 14077
rect 3721 14013 3737 14077
rect 3801 14013 3817 14077
rect 3881 14013 3897 14077
rect 3961 14013 3977 14077
rect 4041 14013 4057 14077
rect 4121 14013 4137 14077
rect 4201 14013 4217 14077
rect 4281 14013 4297 14077
rect 4361 14013 4377 14077
rect 4441 14013 4457 14077
rect 4521 14013 4537 14077
rect 4601 14013 4617 14077
rect 4681 14013 4697 14077
rect 4761 14013 4777 14077
rect 4841 14013 4880 14077
rect 0 14012 4880 14013
rect 10132 18086 15000 18087
rect 10132 14742 10143 18086
rect 14847 14742 15000 18086
rect 10132 14725 15000 14742
rect 10132 14661 10143 14725
rect 10207 14661 10223 14725
rect 10287 14661 10303 14725
rect 10367 14661 10383 14725
rect 10447 14661 10463 14725
rect 10527 14661 10543 14725
rect 10607 14661 10623 14725
rect 10687 14661 10703 14725
rect 10767 14661 10783 14725
rect 10847 14661 10863 14725
rect 10927 14661 10943 14725
rect 11007 14661 11023 14725
rect 11087 14661 11103 14725
rect 11167 14661 11183 14725
rect 11247 14661 11263 14725
rect 11327 14661 11343 14725
rect 11407 14661 11423 14725
rect 11487 14661 11503 14725
rect 11567 14661 11583 14725
rect 11647 14661 11663 14725
rect 11727 14661 11743 14725
rect 11807 14661 11823 14725
rect 11887 14661 11903 14725
rect 11967 14661 11983 14725
rect 12047 14661 12063 14725
rect 12127 14661 12143 14725
rect 12207 14661 12223 14725
rect 12287 14661 12303 14725
rect 12367 14661 12383 14725
rect 12447 14661 12463 14725
rect 12527 14661 12543 14725
rect 12607 14661 12623 14725
rect 12687 14661 12703 14725
rect 12767 14661 12783 14725
rect 12847 14661 12863 14725
rect 12927 14661 12943 14725
rect 13007 14661 13023 14725
rect 13087 14661 13103 14725
rect 13167 14661 13183 14725
rect 13247 14661 13263 14725
rect 13327 14661 13343 14725
rect 13407 14661 13423 14725
rect 13487 14661 13503 14725
rect 13567 14661 13583 14725
rect 13647 14661 13663 14725
rect 13727 14661 13743 14725
rect 13807 14661 13823 14725
rect 13887 14661 13903 14725
rect 13967 14661 13983 14725
rect 14047 14661 14063 14725
rect 14127 14661 14143 14725
rect 14207 14661 14223 14725
rect 14287 14661 14303 14725
rect 14367 14661 14383 14725
rect 14447 14661 14463 14725
rect 14527 14661 14543 14725
rect 14607 14661 14623 14725
rect 14687 14661 14703 14725
rect 14767 14661 14783 14725
rect 14847 14661 15000 14725
rect 10132 14644 15000 14661
rect 10132 14580 10143 14644
rect 10207 14580 10223 14644
rect 10287 14580 10303 14644
rect 10367 14580 10383 14644
rect 10447 14580 10463 14644
rect 10527 14580 10543 14644
rect 10607 14580 10623 14644
rect 10687 14580 10703 14644
rect 10767 14580 10783 14644
rect 10847 14580 10863 14644
rect 10927 14580 10943 14644
rect 11007 14580 11023 14644
rect 11087 14580 11103 14644
rect 11167 14580 11183 14644
rect 11247 14580 11263 14644
rect 11327 14580 11343 14644
rect 11407 14580 11423 14644
rect 11487 14580 11503 14644
rect 11567 14580 11583 14644
rect 11647 14580 11663 14644
rect 11727 14580 11743 14644
rect 11807 14580 11823 14644
rect 11887 14580 11903 14644
rect 11967 14580 11983 14644
rect 12047 14580 12063 14644
rect 12127 14580 12143 14644
rect 12207 14580 12223 14644
rect 12287 14580 12303 14644
rect 12367 14580 12383 14644
rect 12447 14580 12463 14644
rect 12527 14580 12543 14644
rect 12607 14580 12623 14644
rect 12687 14580 12703 14644
rect 12767 14580 12783 14644
rect 12847 14580 12863 14644
rect 12927 14580 12943 14644
rect 13007 14580 13023 14644
rect 13087 14580 13103 14644
rect 13167 14580 13183 14644
rect 13247 14580 13263 14644
rect 13327 14580 13343 14644
rect 13407 14580 13423 14644
rect 13487 14580 13503 14644
rect 13567 14580 13583 14644
rect 13647 14580 13663 14644
rect 13727 14580 13743 14644
rect 13807 14580 13823 14644
rect 13887 14580 13903 14644
rect 13967 14580 13983 14644
rect 14047 14580 14063 14644
rect 14127 14580 14143 14644
rect 14207 14580 14223 14644
rect 14287 14580 14303 14644
rect 14367 14580 14383 14644
rect 14447 14580 14463 14644
rect 14527 14580 14543 14644
rect 14607 14580 14623 14644
rect 14687 14580 14703 14644
rect 14767 14580 14783 14644
rect 14847 14580 15000 14644
rect 10132 14563 15000 14580
rect 10132 14499 10143 14563
rect 10207 14499 10223 14563
rect 10287 14499 10303 14563
rect 10367 14499 10383 14563
rect 10447 14499 10463 14563
rect 10527 14499 10543 14563
rect 10607 14499 10623 14563
rect 10687 14499 10703 14563
rect 10767 14499 10783 14563
rect 10847 14499 10863 14563
rect 10927 14499 10943 14563
rect 11007 14499 11023 14563
rect 11087 14499 11103 14563
rect 11167 14499 11183 14563
rect 11247 14499 11263 14563
rect 11327 14499 11343 14563
rect 11407 14499 11423 14563
rect 11487 14499 11503 14563
rect 11567 14499 11583 14563
rect 11647 14499 11663 14563
rect 11727 14499 11743 14563
rect 11807 14499 11823 14563
rect 11887 14499 11903 14563
rect 11967 14499 11983 14563
rect 12047 14499 12063 14563
rect 12127 14499 12143 14563
rect 12207 14499 12223 14563
rect 12287 14499 12303 14563
rect 12367 14499 12383 14563
rect 12447 14499 12463 14563
rect 12527 14499 12543 14563
rect 12607 14499 12623 14563
rect 12687 14499 12703 14563
rect 12767 14499 12783 14563
rect 12847 14499 12863 14563
rect 12927 14499 12943 14563
rect 13007 14499 13023 14563
rect 13087 14499 13103 14563
rect 13167 14499 13183 14563
rect 13247 14499 13263 14563
rect 13327 14499 13343 14563
rect 13407 14499 13423 14563
rect 13487 14499 13503 14563
rect 13567 14499 13583 14563
rect 13647 14499 13663 14563
rect 13727 14499 13743 14563
rect 13807 14499 13823 14563
rect 13887 14499 13903 14563
rect 13967 14499 13983 14563
rect 14047 14499 14063 14563
rect 14127 14499 14143 14563
rect 14207 14499 14223 14563
rect 14287 14499 14303 14563
rect 14367 14499 14383 14563
rect 14447 14499 14463 14563
rect 14527 14499 14543 14563
rect 14607 14499 14623 14563
rect 14687 14499 14703 14563
rect 14767 14499 14783 14563
rect 14847 14499 15000 14563
rect 10132 14482 15000 14499
rect 10132 14418 10143 14482
rect 10207 14418 10223 14482
rect 10287 14418 10303 14482
rect 10367 14418 10383 14482
rect 10447 14418 10463 14482
rect 10527 14418 10543 14482
rect 10607 14418 10623 14482
rect 10687 14418 10703 14482
rect 10767 14418 10783 14482
rect 10847 14418 10863 14482
rect 10927 14418 10943 14482
rect 11007 14418 11023 14482
rect 11087 14418 11103 14482
rect 11167 14418 11183 14482
rect 11247 14418 11263 14482
rect 11327 14418 11343 14482
rect 11407 14418 11423 14482
rect 11487 14418 11503 14482
rect 11567 14418 11583 14482
rect 11647 14418 11663 14482
rect 11727 14418 11743 14482
rect 11807 14418 11823 14482
rect 11887 14418 11903 14482
rect 11967 14418 11983 14482
rect 12047 14418 12063 14482
rect 12127 14418 12143 14482
rect 12207 14418 12223 14482
rect 12287 14418 12303 14482
rect 12367 14418 12383 14482
rect 12447 14418 12463 14482
rect 12527 14418 12543 14482
rect 12607 14418 12623 14482
rect 12687 14418 12703 14482
rect 12767 14418 12783 14482
rect 12847 14418 12863 14482
rect 12927 14418 12943 14482
rect 13007 14418 13023 14482
rect 13087 14418 13103 14482
rect 13167 14418 13183 14482
rect 13247 14418 13263 14482
rect 13327 14418 13343 14482
rect 13407 14418 13423 14482
rect 13487 14418 13503 14482
rect 13567 14418 13583 14482
rect 13647 14418 13663 14482
rect 13727 14418 13743 14482
rect 13807 14418 13823 14482
rect 13887 14418 13903 14482
rect 13967 14418 13983 14482
rect 14047 14418 14063 14482
rect 14127 14418 14143 14482
rect 14207 14418 14223 14482
rect 14287 14418 14303 14482
rect 14367 14418 14383 14482
rect 14447 14418 14463 14482
rect 14527 14418 14543 14482
rect 14607 14418 14623 14482
rect 14687 14418 14703 14482
rect 14767 14418 14783 14482
rect 14847 14418 15000 14482
rect 10132 14401 15000 14418
rect 10132 14337 10143 14401
rect 10207 14337 10223 14401
rect 10287 14337 10303 14401
rect 10367 14337 10383 14401
rect 10447 14337 10463 14401
rect 10527 14337 10543 14401
rect 10607 14337 10623 14401
rect 10687 14337 10703 14401
rect 10767 14337 10783 14401
rect 10847 14337 10863 14401
rect 10927 14337 10943 14401
rect 11007 14337 11023 14401
rect 11087 14337 11103 14401
rect 11167 14337 11183 14401
rect 11247 14337 11263 14401
rect 11327 14337 11343 14401
rect 11407 14337 11423 14401
rect 11487 14337 11503 14401
rect 11567 14337 11583 14401
rect 11647 14337 11663 14401
rect 11727 14337 11743 14401
rect 11807 14337 11823 14401
rect 11887 14337 11903 14401
rect 11967 14337 11983 14401
rect 12047 14337 12063 14401
rect 12127 14337 12143 14401
rect 12207 14337 12223 14401
rect 12287 14337 12303 14401
rect 12367 14337 12383 14401
rect 12447 14337 12463 14401
rect 12527 14337 12543 14401
rect 12607 14337 12623 14401
rect 12687 14337 12703 14401
rect 12767 14337 12783 14401
rect 12847 14337 12863 14401
rect 12927 14337 12943 14401
rect 13007 14337 13023 14401
rect 13087 14337 13103 14401
rect 13167 14337 13183 14401
rect 13247 14337 13263 14401
rect 13327 14337 13343 14401
rect 13407 14337 13423 14401
rect 13487 14337 13503 14401
rect 13567 14337 13583 14401
rect 13647 14337 13663 14401
rect 13727 14337 13743 14401
rect 13807 14337 13823 14401
rect 13887 14337 13903 14401
rect 13967 14337 13983 14401
rect 14047 14337 14063 14401
rect 14127 14337 14143 14401
rect 14207 14337 14223 14401
rect 14287 14337 14303 14401
rect 14367 14337 14383 14401
rect 14447 14337 14463 14401
rect 14527 14337 14543 14401
rect 14607 14337 14623 14401
rect 14687 14337 14703 14401
rect 14767 14337 14783 14401
rect 14847 14337 15000 14401
rect 10132 14320 15000 14337
rect 10132 14256 10143 14320
rect 10207 14256 10223 14320
rect 10287 14256 10303 14320
rect 10367 14256 10383 14320
rect 10447 14256 10463 14320
rect 10527 14256 10543 14320
rect 10607 14256 10623 14320
rect 10687 14256 10703 14320
rect 10767 14256 10783 14320
rect 10847 14256 10863 14320
rect 10927 14256 10943 14320
rect 11007 14256 11023 14320
rect 11087 14256 11103 14320
rect 11167 14256 11183 14320
rect 11247 14256 11263 14320
rect 11327 14256 11343 14320
rect 11407 14256 11423 14320
rect 11487 14256 11503 14320
rect 11567 14256 11583 14320
rect 11647 14256 11663 14320
rect 11727 14256 11743 14320
rect 11807 14256 11823 14320
rect 11887 14256 11903 14320
rect 11967 14256 11983 14320
rect 12047 14256 12063 14320
rect 12127 14256 12143 14320
rect 12207 14256 12223 14320
rect 12287 14256 12303 14320
rect 12367 14256 12383 14320
rect 12447 14256 12463 14320
rect 12527 14256 12543 14320
rect 12607 14256 12623 14320
rect 12687 14256 12703 14320
rect 12767 14256 12783 14320
rect 12847 14256 12863 14320
rect 12927 14256 12943 14320
rect 13007 14256 13023 14320
rect 13087 14256 13103 14320
rect 13167 14256 13183 14320
rect 13247 14256 13263 14320
rect 13327 14256 13343 14320
rect 13407 14256 13423 14320
rect 13487 14256 13503 14320
rect 13567 14256 13583 14320
rect 13647 14256 13663 14320
rect 13727 14256 13743 14320
rect 13807 14256 13823 14320
rect 13887 14256 13903 14320
rect 13967 14256 13983 14320
rect 14047 14256 14063 14320
rect 14127 14256 14143 14320
rect 14207 14256 14223 14320
rect 14287 14256 14303 14320
rect 14367 14256 14383 14320
rect 14447 14256 14463 14320
rect 14527 14256 14543 14320
rect 14607 14256 14623 14320
rect 14687 14256 14703 14320
rect 14767 14256 14783 14320
rect 14847 14256 15000 14320
rect 10132 14239 15000 14256
rect 10132 14175 10143 14239
rect 10207 14175 10223 14239
rect 10287 14175 10303 14239
rect 10367 14175 10383 14239
rect 10447 14175 10463 14239
rect 10527 14175 10543 14239
rect 10607 14175 10623 14239
rect 10687 14175 10703 14239
rect 10767 14175 10783 14239
rect 10847 14175 10863 14239
rect 10927 14175 10943 14239
rect 11007 14175 11023 14239
rect 11087 14175 11103 14239
rect 11167 14175 11183 14239
rect 11247 14175 11263 14239
rect 11327 14175 11343 14239
rect 11407 14175 11423 14239
rect 11487 14175 11503 14239
rect 11567 14175 11583 14239
rect 11647 14175 11663 14239
rect 11727 14175 11743 14239
rect 11807 14175 11823 14239
rect 11887 14175 11903 14239
rect 11967 14175 11983 14239
rect 12047 14175 12063 14239
rect 12127 14175 12143 14239
rect 12207 14175 12223 14239
rect 12287 14175 12303 14239
rect 12367 14175 12383 14239
rect 12447 14175 12463 14239
rect 12527 14175 12543 14239
rect 12607 14175 12623 14239
rect 12687 14175 12703 14239
rect 12767 14175 12783 14239
rect 12847 14175 12863 14239
rect 12927 14175 12943 14239
rect 13007 14175 13023 14239
rect 13087 14175 13103 14239
rect 13167 14175 13183 14239
rect 13247 14175 13263 14239
rect 13327 14175 13343 14239
rect 13407 14175 13423 14239
rect 13487 14175 13503 14239
rect 13567 14175 13583 14239
rect 13647 14175 13663 14239
rect 13727 14175 13743 14239
rect 13807 14175 13823 14239
rect 13887 14175 13903 14239
rect 13967 14175 13983 14239
rect 14047 14175 14063 14239
rect 14127 14175 14143 14239
rect 14207 14175 14223 14239
rect 14287 14175 14303 14239
rect 14367 14175 14383 14239
rect 14447 14175 14463 14239
rect 14527 14175 14543 14239
rect 14607 14175 14623 14239
rect 14687 14175 14703 14239
rect 14767 14175 14783 14239
rect 14847 14175 15000 14239
rect 10132 14158 15000 14175
rect 10132 14094 10143 14158
rect 10207 14094 10223 14158
rect 10287 14094 10303 14158
rect 10367 14094 10383 14158
rect 10447 14094 10463 14158
rect 10527 14094 10543 14158
rect 10607 14094 10623 14158
rect 10687 14094 10703 14158
rect 10767 14094 10783 14158
rect 10847 14094 10863 14158
rect 10927 14094 10943 14158
rect 11007 14094 11023 14158
rect 11087 14094 11103 14158
rect 11167 14094 11183 14158
rect 11247 14094 11263 14158
rect 11327 14094 11343 14158
rect 11407 14094 11423 14158
rect 11487 14094 11503 14158
rect 11567 14094 11583 14158
rect 11647 14094 11663 14158
rect 11727 14094 11743 14158
rect 11807 14094 11823 14158
rect 11887 14094 11903 14158
rect 11967 14094 11983 14158
rect 12047 14094 12063 14158
rect 12127 14094 12143 14158
rect 12207 14094 12223 14158
rect 12287 14094 12303 14158
rect 12367 14094 12383 14158
rect 12447 14094 12463 14158
rect 12527 14094 12543 14158
rect 12607 14094 12623 14158
rect 12687 14094 12703 14158
rect 12767 14094 12783 14158
rect 12847 14094 12863 14158
rect 12927 14094 12943 14158
rect 13007 14094 13023 14158
rect 13087 14094 13103 14158
rect 13167 14094 13183 14158
rect 13247 14094 13263 14158
rect 13327 14094 13343 14158
rect 13407 14094 13423 14158
rect 13487 14094 13503 14158
rect 13567 14094 13583 14158
rect 13647 14094 13663 14158
rect 13727 14094 13743 14158
rect 13807 14094 13823 14158
rect 13887 14094 13903 14158
rect 13967 14094 13983 14158
rect 14047 14094 14063 14158
rect 14127 14094 14143 14158
rect 14207 14094 14223 14158
rect 14287 14094 14303 14158
rect 14367 14094 14383 14158
rect 14447 14094 14463 14158
rect 14527 14094 14543 14158
rect 14607 14094 14623 14158
rect 14687 14094 14703 14158
rect 14767 14094 14783 14158
rect 14847 14094 15000 14158
rect 10132 14077 15000 14094
rect 10132 14013 10143 14077
rect 10207 14013 10223 14077
rect 10287 14013 10303 14077
rect 10367 14013 10383 14077
rect 10447 14013 10463 14077
rect 10527 14013 10543 14077
rect 10607 14013 10623 14077
rect 10687 14013 10703 14077
rect 10767 14013 10783 14077
rect 10847 14013 10863 14077
rect 10927 14013 10943 14077
rect 11007 14013 11023 14077
rect 11087 14013 11103 14077
rect 11167 14013 11183 14077
rect 11247 14013 11263 14077
rect 11327 14013 11343 14077
rect 11407 14013 11423 14077
rect 11487 14013 11503 14077
rect 11567 14013 11583 14077
rect 11647 14013 11663 14077
rect 11727 14013 11743 14077
rect 11807 14013 11823 14077
rect 11887 14013 11903 14077
rect 11967 14013 11983 14077
rect 12047 14013 12063 14077
rect 12127 14013 12143 14077
rect 12207 14013 12223 14077
rect 12287 14013 12303 14077
rect 12367 14013 12383 14077
rect 12447 14013 12463 14077
rect 12527 14013 12543 14077
rect 12607 14013 12623 14077
rect 12687 14013 12703 14077
rect 12767 14013 12783 14077
rect 12847 14013 12863 14077
rect 12927 14013 12943 14077
rect 13007 14013 13023 14077
rect 13087 14013 13103 14077
rect 13167 14013 13183 14077
rect 13247 14013 13263 14077
rect 13327 14013 13343 14077
rect 13407 14013 13423 14077
rect 13487 14013 13503 14077
rect 13567 14013 13583 14077
rect 13647 14013 13663 14077
rect 13727 14013 13743 14077
rect 13807 14013 13823 14077
rect 13887 14013 13903 14077
rect 13967 14013 13983 14077
rect 14047 14013 14063 14077
rect 14127 14013 14143 14077
rect 14207 14013 14223 14077
rect 14287 14013 14303 14077
rect 14367 14013 14383 14077
rect 14447 14013 14463 14077
rect 14527 14013 14543 14077
rect 14607 14013 14623 14077
rect 14687 14013 14703 14077
rect 14767 14013 14783 14077
rect 14847 14013 15000 14077
rect 10132 14012 15000 14013
rect 0 14007 254 14012
rect 14746 14007 15000 14012
rect 0 13704 4874 13707
rect 0 13640 105 13704
rect 169 13640 186 13704
rect 250 13640 267 13704
rect 331 13640 348 13704
rect 412 13640 429 13704
rect 493 13640 510 13704
rect 574 13640 591 13704
rect 655 13640 672 13704
rect 736 13640 753 13704
rect 817 13640 834 13704
rect 898 13640 915 13704
rect 979 13640 996 13704
rect 1060 13640 1077 13704
rect 1141 13640 1158 13704
rect 1222 13640 1239 13704
rect 1303 13640 1320 13704
rect 1384 13640 1401 13704
rect 1465 13640 1482 13704
rect 1546 13640 1563 13704
rect 1627 13640 1644 13704
rect 1708 13640 1725 13704
rect 1789 13640 1806 13704
rect 1870 13640 1887 13704
rect 1951 13640 1968 13704
rect 2032 13640 2049 13704
rect 2113 13640 2130 13704
rect 2194 13640 2211 13704
rect 2275 13640 2292 13704
rect 2356 13640 2373 13704
rect 2437 13640 2454 13704
rect 2518 13640 2535 13704
rect 2599 13640 2616 13704
rect 2680 13640 2697 13704
rect 2761 13640 2778 13704
rect 2842 13640 2859 13704
rect 2923 13640 2940 13704
rect 3004 13640 3021 13704
rect 3085 13640 3102 13704
rect 3166 13640 3183 13704
rect 3247 13640 3264 13704
rect 3328 13640 3345 13704
rect 3409 13640 3426 13704
rect 3490 13640 3507 13704
rect 3571 13640 3588 13704
rect 3652 13640 3669 13704
rect 3733 13640 3750 13704
rect 3814 13640 3831 13704
rect 3895 13640 3912 13704
rect 3976 13640 3993 13704
rect 4057 13640 4074 13704
rect 4138 13640 4155 13704
rect 4219 13640 4236 13704
rect 4300 13640 4317 13704
rect 4381 13640 4399 13704
rect 4463 13640 4481 13704
rect 4545 13640 4563 13704
rect 4627 13640 4645 13704
rect 4709 13640 4727 13704
rect 4791 13640 4809 13704
rect 4873 13640 4874 13704
rect 0 13622 4874 13640
rect 0 13558 105 13622
rect 169 13558 186 13622
rect 250 13558 267 13622
rect 331 13558 348 13622
rect 412 13558 429 13622
rect 493 13558 510 13622
rect 574 13558 591 13622
rect 655 13558 672 13622
rect 736 13558 753 13622
rect 817 13558 834 13622
rect 898 13558 915 13622
rect 979 13558 996 13622
rect 1060 13558 1077 13622
rect 1141 13558 1158 13622
rect 1222 13558 1239 13622
rect 1303 13558 1320 13622
rect 1384 13558 1401 13622
rect 1465 13558 1482 13622
rect 1546 13558 1563 13622
rect 1627 13558 1644 13622
rect 1708 13558 1725 13622
rect 1789 13558 1806 13622
rect 1870 13558 1887 13622
rect 1951 13558 1968 13622
rect 2032 13558 2049 13622
rect 2113 13558 2130 13622
rect 2194 13558 2211 13622
rect 2275 13558 2292 13622
rect 2356 13558 2373 13622
rect 2437 13558 2454 13622
rect 2518 13558 2535 13622
rect 2599 13558 2616 13622
rect 2680 13558 2697 13622
rect 2761 13558 2778 13622
rect 2842 13558 2859 13622
rect 2923 13558 2940 13622
rect 3004 13558 3021 13622
rect 3085 13558 3102 13622
rect 3166 13558 3183 13622
rect 3247 13558 3264 13622
rect 3328 13558 3345 13622
rect 3409 13558 3426 13622
rect 3490 13558 3507 13622
rect 3571 13558 3588 13622
rect 3652 13558 3669 13622
rect 3733 13558 3750 13622
rect 3814 13558 3831 13622
rect 3895 13558 3912 13622
rect 3976 13558 3993 13622
rect 4057 13558 4074 13622
rect 4138 13558 4155 13622
rect 4219 13558 4236 13622
rect 4300 13558 4317 13622
rect 4381 13558 4399 13622
rect 4463 13558 4481 13622
rect 4545 13558 4563 13622
rect 4627 13558 4645 13622
rect 4709 13558 4727 13622
rect 4791 13558 4809 13622
rect 4873 13558 4874 13622
rect 0 13540 4874 13558
rect 0 13476 105 13540
rect 169 13476 186 13540
rect 250 13476 267 13540
rect 331 13476 348 13540
rect 412 13476 429 13540
rect 493 13476 510 13540
rect 574 13476 591 13540
rect 655 13476 672 13540
rect 736 13476 753 13540
rect 817 13476 834 13540
rect 898 13476 915 13540
rect 979 13476 996 13540
rect 1060 13476 1077 13540
rect 1141 13476 1158 13540
rect 1222 13476 1239 13540
rect 1303 13476 1320 13540
rect 1384 13476 1401 13540
rect 1465 13476 1482 13540
rect 1546 13476 1563 13540
rect 1627 13476 1644 13540
rect 1708 13476 1725 13540
rect 1789 13476 1806 13540
rect 1870 13476 1887 13540
rect 1951 13476 1968 13540
rect 2032 13476 2049 13540
rect 2113 13476 2130 13540
rect 2194 13476 2211 13540
rect 2275 13476 2292 13540
rect 2356 13476 2373 13540
rect 2437 13476 2454 13540
rect 2518 13476 2535 13540
rect 2599 13476 2616 13540
rect 2680 13476 2697 13540
rect 2761 13476 2778 13540
rect 2842 13476 2859 13540
rect 2923 13476 2940 13540
rect 3004 13476 3021 13540
rect 3085 13476 3102 13540
rect 3166 13476 3183 13540
rect 3247 13476 3264 13540
rect 3328 13476 3345 13540
rect 3409 13476 3426 13540
rect 3490 13476 3507 13540
rect 3571 13476 3588 13540
rect 3652 13476 3669 13540
rect 3733 13476 3750 13540
rect 3814 13476 3831 13540
rect 3895 13476 3912 13540
rect 3976 13476 3993 13540
rect 4057 13476 4074 13540
rect 4138 13476 4155 13540
rect 4219 13476 4236 13540
rect 4300 13476 4317 13540
rect 4381 13476 4399 13540
rect 4463 13476 4481 13540
rect 4545 13476 4563 13540
rect 4627 13476 4645 13540
rect 4709 13476 4727 13540
rect 4791 13476 4809 13540
rect 4873 13476 4874 13540
rect 0 13458 4874 13476
rect 0 13394 105 13458
rect 169 13394 186 13458
rect 250 13394 267 13458
rect 331 13394 348 13458
rect 412 13394 429 13458
rect 493 13394 510 13458
rect 574 13394 591 13458
rect 655 13394 672 13458
rect 736 13394 753 13458
rect 817 13394 834 13458
rect 898 13394 915 13458
rect 979 13394 996 13458
rect 1060 13394 1077 13458
rect 1141 13394 1158 13458
rect 1222 13394 1239 13458
rect 1303 13394 1320 13458
rect 1384 13394 1401 13458
rect 1465 13394 1482 13458
rect 1546 13394 1563 13458
rect 1627 13394 1644 13458
rect 1708 13394 1725 13458
rect 1789 13394 1806 13458
rect 1870 13394 1887 13458
rect 1951 13394 1968 13458
rect 2032 13394 2049 13458
rect 2113 13394 2130 13458
rect 2194 13394 2211 13458
rect 2275 13394 2292 13458
rect 2356 13394 2373 13458
rect 2437 13394 2454 13458
rect 2518 13394 2535 13458
rect 2599 13394 2616 13458
rect 2680 13394 2697 13458
rect 2761 13394 2778 13458
rect 2842 13394 2859 13458
rect 2923 13394 2940 13458
rect 3004 13394 3021 13458
rect 3085 13394 3102 13458
rect 3166 13394 3183 13458
rect 3247 13394 3264 13458
rect 3328 13394 3345 13458
rect 3409 13394 3426 13458
rect 3490 13394 3507 13458
rect 3571 13394 3588 13458
rect 3652 13394 3669 13458
rect 3733 13394 3750 13458
rect 3814 13394 3831 13458
rect 3895 13394 3912 13458
rect 3976 13394 3993 13458
rect 4057 13394 4074 13458
rect 4138 13394 4155 13458
rect 4219 13394 4236 13458
rect 4300 13394 4317 13458
rect 4381 13394 4399 13458
rect 4463 13394 4481 13458
rect 4545 13394 4563 13458
rect 4627 13394 4645 13458
rect 4709 13394 4727 13458
rect 4791 13394 4809 13458
rect 4873 13394 4874 13458
rect 0 13376 4874 13394
rect 0 13312 105 13376
rect 169 13312 186 13376
rect 250 13312 267 13376
rect 331 13312 348 13376
rect 412 13312 429 13376
rect 493 13312 510 13376
rect 574 13312 591 13376
rect 655 13312 672 13376
rect 736 13312 753 13376
rect 817 13312 834 13376
rect 898 13312 915 13376
rect 979 13312 996 13376
rect 1060 13312 1077 13376
rect 1141 13312 1158 13376
rect 1222 13312 1239 13376
rect 1303 13312 1320 13376
rect 1384 13312 1401 13376
rect 1465 13312 1482 13376
rect 1546 13312 1563 13376
rect 1627 13312 1644 13376
rect 1708 13312 1725 13376
rect 1789 13312 1806 13376
rect 1870 13312 1887 13376
rect 1951 13312 1968 13376
rect 2032 13312 2049 13376
rect 2113 13312 2130 13376
rect 2194 13312 2211 13376
rect 2275 13312 2292 13376
rect 2356 13312 2373 13376
rect 2437 13312 2454 13376
rect 2518 13312 2535 13376
rect 2599 13312 2616 13376
rect 2680 13312 2697 13376
rect 2761 13312 2778 13376
rect 2842 13312 2859 13376
rect 2923 13312 2940 13376
rect 3004 13312 3021 13376
rect 3085 13312 3102 13376
rect 3166 13312 3183 13376
rect 3247 13312 3264 13376
rect 3328 13312 3345 13376
rect 3409 13312 3426 13376
rect 3490 13312 3507 13376
rect 3571 13312 3588 13376
rect 3652 13312 3669 13376
rect 3733 13312 3750 13376
rect 3814 13312 3831 13376
rect 3895 13312 3912 13376
rect 3976 13312 3993 13376
rect 4057 13312 4074 13376
rect 4138 13312 4155 13376
rect 4219 13312 4236 13376
rect 4300 13312 4317 13376
rect 4381 13312 4399 13376
rect 4463 13312 4481 13376
rect 4545 13312 4563 13376
rect 4627 13312 4645 13376
rect 4709 13312 4727 13376
rect 4791 13312 4809 13376
rect 4873 13312 4874 13376
rect 0 13294 4874 13312
rect 0 13230 105 13294
rect 169 13230 186 13294
rect 250 13230 267 13294
rect 331 13230 348 13294
rect 412 13230 429 13294
rect 493 13230 510 13294
rect 574 13230 591 13294
rect 655 13230 672 13294
rect 736 13230 753 13294
rect 817 13230 834 13294
rect 898 13230 915 13294
rect 979 13230 996 13294
rect 1060 13230 1077 13294
rect 1141 13230 1158 13294
rect 1222 13230 1239 13294
rect 1303 13230 1320 13294
rect 1384 13230 1401 13294
rect 1465 13230 1482 13294
rect 1546 13230 1563 13294
rect 1627 13230 1644 13294
rect 1708 13230 1725 13294
rect 1789 13230 1806 13294
rect 1870 13230 1887 13294
rect 1951 13230 1968 13294
rect 2032 13230 2049 13294
rect 2113 13230 2130 13294
rect 2194 13230 2211 13294
rect 2275 13230 2292 13294
rect 2356 13230 2373 13294
rect 2437 13230 2454 13294
rect 2518 13230 2535 13294
rect 2599 13230 2616 13294
rect 2680 13230 2697 13294
rect 2761 13230 2778 13294
rect 2842 13230 2859 13294
rect 2923 13230 2940 13294
rect 3004 13230 3021 13294
rect 3085 13230 3102 13294
rect 3166 13230 3183 13294
rect 3247 13230 3264 13294
rect 3328 13230 3345 13294
rect 3409 13230 3426 13294
rect 3490 13230 3507 13294
rect 3571 13230 3588 13294
rect 3652 13230 3669 13294
rect 3733 13230 3750 13294
rect 3814 13230 3831 13294
rect 3895 13230 3912 13294
rect 3976 13230 3993 13294
rect 4057 13230 4074 13294
rect 4138 13230 4155 13294
rect 4219 13230 4236 13294
rect 4300 13230 4317 13294
rect 4381 13230 4399 13294
rect 4463 13230 4481 13294
rect 4545 13230 4563 13294
rect 4627 13230 4645 13294
rect 4709 13230 4727 13294
rect 4791 13230 4809 13294
rect 4873 13230 4874 13294
rect 0 13212 4874 13230
rect 0 13148 105 13212
rect 169 13148 186 13212
rect 250 13148 267 13212
rect 331 13148 348 13212
rect 412 13148 429 13212
rect 493 13148 510 13212
rect 574 13148 591 13212
rect 655 13148 672 13212
rect 736 13148 753 13212
rect 817 13148 834 13212
rect 898 13148 915 13212
rect 979 13148 996 13212
rect 1060 13148 1077 13212
rect 1141 13148 1158 13212
rect 1222 13148 1239 13212
rect 1303 13148 1320 13212
rect 1384 13148 1401 13212
rect 1465 13148 1482 13212
rect 1546 13148 1563 13212
rect 1627 13148 1644 13212
rect 1708 13148 1725 13212
rect 1789 13148 1806 13212
rect 1870 13148 1887 13212
rect 1951 13148 1968 13212
rect 2032 13148 2049 13212
rect 2113 13148 2130 13212
rect 2194 13148 2211 13212
rect 2275 13148 2292 13212
rect 2356 13148 2373 13212
rect 2437 13148 2454 13212
rect 2518 13148 2535 13212
rect 2599 13148 2616 13212
rect 2680 13148 2697 13212
rect 2761 13148 2778 13212
rect 2842 13148 2859 13212
rect 2923 13148 2940 13212
rect 3004 13148 3021 13212
rect 3085 13148 3102 13212
rect 3166 13148 3183 13212
rect 3247 13148 3264 13212
rect 3328 13148 3345 13212
rect 3409 13148 3426 13212
rect 3490 13148 3507 13212
rect 3571 13148 3588 13212
rect 3652 13148 3669 13212
rect 3733 13148 3750 13212
rect 3814 13148 3831 13212
rect 3895 13148 3912 13212
rect 3976 13148 3993 13212
rect 4057 13148 4074 13212
rect 4138 13148 4155 13212
rect 4219 13148 4236 13212
rect 4300 13148 4317 13212
rect 4381 13148 4399 13212
rect 4463 13148 4481 13212
rect 4545 13148 4563 13212
rect 4627 13148 4645 13212
rect 4709 13148 4727 13212
rect 4791 13148 4809 13212
rect 4873 13148 4874 13212
rect 0 13130 4874 13148
rect 0 13066 105 13130
rect 169 13066 186 13130
rect 250 13066 267 13130
rect 331 13066 348 13130
rect 412 13066 429 13130
rect 493 13066 510 13130
rect 574 13066 591 13130
rect 655 13066 672 13130
rect 736 13066 753 13130
rect 817 13066 834 13130
rect 898 13066 915 13130
rect 979 13066 996 13130
rect 1060 13066 1077 13130
rect 1141 13066 1158 13130
rect 1222 13066 1239 13130
rect 1303 13066 1320 13130
rect 1384 13066 1401 13130
rect 1465 13066 1482 13130
rect 1546 13066 1563 13130
rect 1627 13066 1644 13130
rect 1708 13066 1725 13130
rect 1789 13066 1806 13130
rect 1870 13066 1887 13130
rect 1951 13066 1968 13130
rect 2032 13066 2049 13130
rect 2113 13066 2130 13130
rect 2194 13066 2211 13130
rect 2275 13066 2292 13130
rect 2356 13066 2373 13130
rect 2437 13066 2454 13130
rect 2518 13066 2535 13130
rect 2599 13066 2616 13130
rect 2680 13066 2697 13130
rect 2761 13066 2778 13130
rect 2842 13066 2859 13130
rect 2923 13066 2940 13130
rect 3004 13066 3021 13130
rect 3085 13066 3102 13130
rect 3166 13066 3183 13130
rect 3247 13066 3264 13130
rect 3328 13066 3345 13130
rect 3409 13066 3426 13130
rect 3490 13066 3507 13130
rect 3571 13066 3588 13130
rect 3652 13066 3669 13130
rect 3733 13066 3750 13130
rect 3814 13066 3831 13130
rect 3895 13066 3912 13130
rect 3976 13066 3993 13130
rect 4057 13066 4074 13130
rect 4138 13066 4155 13130
rect 4219 13066 4236 13130
rect 4300 13066 4317 13130
rect 4381 13066 4399 13130
rect 4463 13066 4481 13130
rect 4545 13066 4563 13130
rect 4627 13066 4645 13130
rect 4709 13066 4727 13130
rect 4791 13066 4809 13130
rect 4873 13066 4874 13130
rect 0 13048 4874 13066
rect 0 12984 105 13048
rect 169 12984 186 13048
rect 250 12984 267 13048
rect 331 12984 348 13048
rect 412 12984 429 13048
rect 493 12984 510 13048
rect 574 12984 591 13048
rect 655 12984 672 13048
rect 736 12984 753 13048
rect 817 12984 834 13048
rect 898 12984 915 13048
rect 979 12984 996 13048
rect 1060 12984 1077 13048
rect 1141 12984 1158 13048
rect 1222 12984 1239 13048
rect 1303 12984 1320 13048
rect 1384 12984 1401 13048
rect 1465 12984 1482 13048
rect 1546 12984 1563 13048
rect 1627 12984 1644 13048
rect 1708 12984 1725 13048
rect 1789 12984 1806 13048
rect 1870 12984 1887 13048
rect 1951 12984 1968 13048
rect 2032 12984 2049 13048
rect 2113 12984 2130 13048
rect 2194 12984 2211 13048
rect 2275 12984 2292 13048
rect 2356 12984 2373 13048
rect 2437 12984 2454 13048
rect 2518 12984 2535 13048
rect 2599 12984 2616 13048
rect 2680 12984 2697 13048
rect 2761 12984 2778 13048
rect 2842 12984 2859 13048
rect 2923 12984 2940 13048
rect 3004 12984 3021 13048
rect 3085 12984 3102 13048
rect 3166 12984 3183 13048
rect 3247 12984 3264 13048
rect 3328 12984 3345 13048
rect 3409 12984 3426 13048
rect 3490 12984 3507 13048
rect 3571 12984 3588 13048
rect 3652 12984 3669 13048
rect 3733 12984 3750 13048
rect 3814 12984 3831 13048
rect 3895 12984 3912 13048
rect 3976 12984 3993 13048
rect 4057 12984 4074 13048
rect 4138 12984 4155 13048
rect 4219 12984 4236 13048
rect 4300 12984 4317 13048
rect 4381 12984 4399 13048
rect 4463 12984 4481 13048
rect 4545 12984 4563 13048
rect 4627 12984 4645 13048
rect 4709 12984 4727 13048
rect 4791 12984 4809 13048
rect 4873 12984 4874 13048
rect 0 12966 4874 12984
rect 0 12902 105 12966
rect 169 12902 186 12966
rect 250 12902 267 12966
rect 331 12902 348 12966
rect 412 12902 429 12966
rect 493 12902 510 12966
rect 574 12902 591 12966
rect 655 12902 672 12966
rect 736 12902 753 12966
rect 817 12902 834 12966
rect 898 12902 915 12966
rect 979 12902 996 12966
rect 1060 12902 1077 12966
rect 1141 12902 1158 12966
rect 1222 12902 1239 12966
rect 1303 12902 1320 12966
rect 1384 12902 1401 12966
rect 1465 12902 1482 12966
rect 1546 12902 1563 12966
rect 1627 12902 1644 12966
rect 1708 12902 1725 12966
rect 1789 12902 1806 12966
rect 1870 12902 1887 12966
rect 1951 12902 1968 12966
rect 2032 12902 2049 12966
rect 2113 12902 2130 12966
rect 2194 12902 2211 12966
rect 2275 12902 2292 12966
rect 2356 12902 2373 12966
rect 2437 12902 2454 12966
rect 2518 12902 2535 12966
rect 2599 12902 2616 12966
rect 2680 12902 2697 12966
rect 2761 12902 2778 12966
rect 2842 12902 2859 12966
rect 2923 12902 2940 12966
rect 3004 12902 3021 12966
rect 3085 12902 3102 12966
rect 3166 12902 3183 12966
rect 3247 12902 3264 12966
rect 3328 12902 3345 12966
rect 3409 12902 3426 12966
rect 3490 12902 3507 12966
rect 3571 12902 3588 12966
rect 3652 12902 3669 12966
rect 3733 12902 3750 12966
rect 3814 12902 3831 12966
rect 3895 12902 3912 12966
rect 3976 12902 3993 12966
rect 4057 12902 4074 12966
rect 4138 12902 4155 12966
rect 4219 12902 4236 12966
rect 4300 12902 4317 12966
rect 4381 12902 4399 12966
rect 4463 12902 4481 12966
rect 4545 12902 4563 12966
rect 4627 12902 4645 12966
rect 4709 12902 4727 12966
rect 4791 12902 4809 12966
rect 4873 12902 4874 12966
rect 0 12884 4874 12902
rect 0 12820 105 12884
rect 169 12820 186 12884
rect 250 12820 267 12884
rect 331 12820 348 12884
rect 412 12820 429 12884
rect 493 12820 510 12884
rect 574 12820 591 12884
rect 655 12820 672 12884
rect 736 12820 753 12884
rect 817 12820 834 12884
rect 898 12820 915 12884
rect 979 12820 996 12884
rect 1060 12820 1077 12884
rect 1141 12820 1158 12884
rect 1222 12820 1239 12884
rect 1303 12820 1320 12884
rect 1384 12820 1401 12884
rect 1465 12820 1482 12884
rect 1546 12820 1563 12884
rect 1627 12820 1644 12884
rect 1708 12820 1725 12884
rect 1789 12820 1806 12884
rect 1870 12820 1887 12884
rect 1951 12820 1968 12884
rect 2032 12820 2049 12884
rect 2113 12820 2130 12884
rect 2194 12820 2211 12884
rect 2275 12820 2292 12884
rect 2356 12820 2373 12884
rect 2437 12820 2454 12884
rect 2518 12820 2535 12884
rect 2599 12820 2616 12884
rect 2680 12820 2697 12884
rect 2761 12820 2778 12884
rect 2842 12820 2859 12884
rect 2923 12820 2940 12884
rect 3004 12820 3021 12884
rect 3085 12820 3102 12884
rect 3166 12820 3183 12884
rect 3247 12820 3264 12884
rect 3328 12820 3345 12884
rect 3409 12820 3426 12884
rect 3490 12820 3507 12884
rect 3571 12820 3588 12884
rect 3652 12820 3669 12884
rect 3733 12820 3750 12884
rect 3814 12820 3831 12884
rect 3895 12820 3912 12884
rect 3976 12820 3993 12884
rect 4057 12820 4074 12884
rect 4138 12820 4155 12884
rect 4219 12820 4236 12884
rect 4300 12820 4317 12884
rect 4381 12820 4399 12884
rect 4463 12820 4481 12884
rect 4545 12820 4563 12884
rect 4627 12820 4645 12884
rect 4709 12820 4727 12884
rect 4791 12820 4809 12884
rect 4873 12820 4874 12884
rect 0 12817 4874 12820
rect 10083 13704 15000 13707
rect 10083 13640 10084 13704
rect 10148 13640 10165 13704
rect 10229 13640 10246 13704
rect 10310 13640 10327 13704
rect 10391 13640 10408 13704
rect 10472 13640 10489 13704
rect 10553 13640 10570 13704
rect 10634 13640 10651 13704
rect 10715 13640 10732 13704
rect 10796 13640 10813 13704
rect 10877 13640 10894 13704
rect 10958 13640 10975 13704
rect 11039 13640 11056 13704
rect 11120 13640 11137 13704
rect 11201 13640 11218 13704
rect 11282 13640 11299 13704
rect 11363 13640 11380 13704
rect 11444 13640 11461 13704
rect 11525 13640 11542 13704
rect 11606 13640 11623 13704
rect 11687 13640 11704 13704
rect 11768 13640 11785 13704
rect 11849 13640 11866 13704
rect 11930 13640 11947 13704
rect 12011 13640 12028 13704
rect 12092 13640 12109 13704
rect 12173 13640 12190 13704
rect 12254 13640 12271 13704
rect 12335 13640 12352 13704
rect 12416 13640 12433 13704
rect 12497 13640 12514 13704
rect 12578 13640 12595 13704
rect 12659 13640 12676 13704
rect 12740 13640 12757 13704
rect 12821 13640 12838 13704
rect 12902 13640 12919 13704
rect 12983 13640 13000 13704
rect 13064 13640 13081 13704
rect 13145 13640 13162 13704
rect 13226 13640 13243 13704
rect 13307 13640 13324 13704
rect 13388 13640 13405 13704
rect 13469 13640 13486 13704
rect 13550 13640 13567 13704
rect 13631 13640 13648 13704
rect 13712 13640 13729 13704
rect 13793 13640 13810 13704
rect 13874 13640 13891 13704
rect 13955 13640 13972 13704
rect 14036 13640 14053 13704
rect 14117 13640 14134 13704
rect 14198 13640 14215 13704
rect 14279 13640 14296 13704
rect 14360 13640 14378 13704
rect 14442 13640 14460 13704
rect 14524 13640 14542 13704
rect 14606 13640 14624 13704
rect 14688 13640 14706 13704
rect 14770 13640 14788 13704
rect 14852 13640 15000 13704
rect 10083 13622 15000 13640
rect 10083 13558 10084 13622
rect 10148 13558 10165 13622
rect 10229 13558 10246 13622
rect 10310 13558 10327 13622
rect 10391 13558 10408 13622
rect 10472 13558 10489 13622
rect 10553 13558 10570 13622
rect 10634 13558 10651 13622
rect 10715 13558 10732 13622
rect 10796 13558 10813 13622
rect 10877 13558 10894 13622
rect 10958 13558 10975 13622
rect 11039 13558 11056 13622
rect 11120 13558 11137 13622
rect 11201 13558 11218 13622
rect 11282 13558 11299 13622
rect 11363 13558 11380 13622
rect 11444 13558 11461 13622
rect 11525 13558 11542 13622
rect 11606 13558 11623 13622
rect 11687 13558 11704 13622
rect 11768 13558 11785 13622
rect 11849 13558 11866 13622
rect 11930 13558 11947 13622
rect 12011 13558 12028 13622
rect 12092 13558 12109 13622
rect 12173 13558 12190 13622
rect 12254 13558 12271 13622
rect 12335 13558 12352 13622
rect 12416 13558 12433 13622
rect 12497 13558 12514 13622
rect 12578 13558 12595 13622
rect 12659 13558 12676 13622
rect 12740 13558 12757 13622
rect 12821 13558 12838 13622
rect 12902 13558 12919 13622
rect 12983 13558 13000 13622
rect 13064 13558 13081 13622
rect 13145 13558 13162 13622
rect 13226 13558 13243 13622
rect 13307 13558 13324 13622
rect 13388 13558 13405 13622
rect 13469 13558 13486 13622
rect 13550 13558 13567 13622
rect 13631 13558 13648 13622
rect 13712 13558 13729 13622
rect 13793 13558 13810 13622
rect 13874 13558 13891 13622
rect 13955 13558 13972 13622
rect 14036 13558 14053 13622
rect 14117 13558 14134 13622
rect 14198 13558 14215 13622
rect 14279 13558 14296 13622
rect 14360 13558 14378 13622
rect 14442 13558 14460 13622
rect 14524 13558 14542 13622
rect 14606 13558 14624 13622
rect 14688 13558 14706 13622
rect 14770 13558 14788 13622
rect 14852 13558 15000 13622
rect 10083 13540 15000 13558
rect 10083 13476 10084 13540
rect 10148 13476 10165 13540
rect 10229 13476 10246 13540
rect 10310 13476 10327 13540
rect 10391 13476 10408 13540
rect 10472 13476 10489 13540
rect 10553 13476 10570 13540
rect 10634 13476 10651 13540
rect 10715 13476 10732 13540
rect 10796 13476 10813 13540
rect 10877 13476 10894 13540
rect 10958 13476 10975 13540
rect 11039 13476 11056 13540
rect 11120 13476 11137 13540
rect 11201 13476 11218 13540
rect 11282 13476 11299 13540
rect 11363 13476 11380 13540
rect 11444 13476 11461 13540
rect 11525 13476 11542 13540
rect 11606 13476 11623 13540
rect 11687 13476 11704 13540
rect 11768 13476 11785 13540
rect 11849 13476 11866 13540
rect 11930 13476 11947 13540
rect 12011 13476 12028 13540
rect 12092 13476 12109 13540
rect 12173 13476 12190 13540
rect 12254 13476 12271 13540
rect 12335 13476 12352 13540
rect 12416 13476 12433 13540
rect 12497 13476 12514 13540
rect 12578 13476 12595 13540
rect 12659 13476 12676 13540
rect 12740 13476 12757 13540
rect 12821 13476 12838 13540
rect 12902 13476 12919 13540
rect 12983 13476 13000 13540
rect 13064 13476 13081 13540
rect 13145 13476 13162 13540
rect 13226 13476 13243 13540
rect 13307 13476 13324 13540
rect 13388 13476 13405 13540
rect 13469 13476 13486 13540
rect 13550 13476 13567 13540
rect 13631 13476 13648 13540
rect 13712 13476 13729 13540
rect 13793 13476 13810 13540
rect 13874 13476 13891 13540
rect 13955 13476 13972 13540
rect 14036 13476 14053 13540
rect 14117 13476 14134 13540
rect 14198 13476 14215 13540
rect 14279 13476 14296 13540
rect 14360 13476 14378 13540
rect 14442 13476 14460 13540
rect 14524 13476 14542 13540
rect 14606 13476 14624 13540
rect 14688 13476 14706 13540
rect 14770 13476 14788 13540
rect 14852 13476 15000 13540
rect 10083 13458 15000 13476
rect 10083 13394 10084 13458
rect 10148 13394 10165 13458
rect 10229 13394 10246 13458
rect 10310 13394 10327 13458
rect 10391 13394 10408 13458
rect 10472 13394 10489 13458
rect 10553 13394 10570 13458
rect 10634 13394 10651 13458
rect 10715 13394 10732 13458
rect 10796 13394 10813 13458
rect 10877 13394 10894 13458
rect 10958 13394 10975 13458
rect 11039 13394 11056 13458
rect 11120 13394 11137 13458
rect 11201 13394 11218 13458
rect 11282 13394 11299 13458
rect 11363 13394 11380 13458
rect 11444 13394 11461 13458
rect 11525 13394 11542 13458
rect 11606 13394 11623 13458
rect 11687 13394 11704 13458
rect 11768 13394 11785 13458
rect 11849 13394 11866 13458
rect 11930 13394 11947 13458
rect 12011 13394 12028 13458
rect 12092 13394 12109 13458
rect 12173 13394 12190 13458
rect 12254 13394 12271 13458
rect 12335 13394 12352 13458
rect 12416 13394 12433 13458
rect 12497 13394 12514 13458
rect 12578 13394 12595 13458
rect 12659 13394 12676 13458
rect 12740 13394 12757 13458
rect 12821 13394 12838 13458
rect 12902 13394 12919 13458
rect 12983 13394 13000 13458
rect 13064 13394 13081 13458
rect 13145 13394 13162 13458
rect 13226 13394 13243 13458
rect 13307 13394 13324 13458
rect 13388 13394 13405 13458
rect 13469 13394 13486 13458
rect 13550 13394 13567 13458
rect 13631 13394 13648 13458
rect 13712 13394 13729 13458
rect 13793 13394 13810 13458
rect 13874 13394 13891 13458
rect 13955 13394 13972 13458
rect 14036 13394 14053 13458
rect 14117 13394 14134 13458
rect 14198 13394 14215 13458
rect 14279 13394 14296 13458
rect 14360 13394 14378 13458
rect 14442 13394 14460 13458
rect 14524 13394 14542 13458
rect 14606 13394 14624 13458
rect 14688 13394 14706 13458
rect 14770 13394 14788 13458
rect 14852 13394 15000 13458
rect 10083 13376 15000 13394
rect 10083 13312 10084 13376
rect 10148 13312 10165 13376
rect 10229 13312 10246 13376
rect 10310 13312 10327 13376
rect 10391 13312 10408 13376
rect 10472 13312 10489 13376
rect 10553 13312 10570 13376
rect 10634 13312 10651 13376
rect 10715 13312 10732 13376
rect 10796 13312 10813 13376
rect 10877 13312 10894 13376
rect 10958 13312 10975 13376
rect 11039 13312 11056 13376
rect 11120 13312 11137 13376
rect 11201 13312 11218 13376
rect 11282 13312 11299 13376
rect 11363 13312 11380 13376
rect 11444 13312 11461 13376
rect 11525 13312 11542 13376
rect 11606 13312 11623 13376
rect 11687 13312 11704 13376
rect 11768 13312 11785 13376
rect 11849 13312 11866 13376
rect 11930 13312 11947 13376
rect 12011 13312 12028 13376
rect 12092 13312 12109 13376
rect 12173 13312 12190 13376
rect 12254 13312 12271 13376
rect 12335 13312 12352 13376
rect 12416 13312 12433 13376
rect 12497 13312 12514 13376
rect 12578 13312 12595 13376
rect 12659 13312 12676 13376
rect 12740 13312 12757 13376
rect 12821 13312 12838 13376
rect 12902 13312 12919 13376
rect 12983 13312 13000 13376
rect 13064 13312 13081 13376
rect 13145 13312 13162 13376
rect 13226 13312 13243 13376
rect 13307 13312 13324 13376
rect 13388 13312 13405 13376
rect 13469 13312 13486 13376
rect 13550 13312 13567 13376
rect 13631 13312 13648 13376
rect 13712 13312 13729 13376
rect 13793 13312 13810 13376
rect 13874 13312 13891 13376
rect 13955 13312 13972 13376
rect 14036 13312 14053 13376
rect 14117 13312 14134 13376
rect 14198 13312 14215 13376
rect 14279 13312 14296 13376
rect 14360 13312 14378 13376
rect 14442 13312 14460 13376
rect 14524 13312 14542 13376
rect 14606 13312 14624 13376
rect 14688 13312 14706 13376
rect 14770 13312 14788 13376
rect 14852 13312 15000 13376
rect 10083 13294 15000 13312
rect 10083 13230 10084 13294
rect 10148 13230 10165 13294
rect 10229 13230 10246 13294
rect 10310 13230 10327 13294
rect 10391 13230 10408 13294
rect 10472 13230 10489 13294
rect 10553 13230 10570 13294
rect 10634 13230 10651 13294
rect 10715 13230 10732 13294
rect 10796 13230 10813 13294
rect 10877 13230 10894 13294
rect 10958 13230 10975 13294
rect 11039 13230 11056 13294
rect 11120 13230 11137 13294
rect 11201 13230 11218 13294
rect 11282 13230 11299 13294
rect 11363 13230 11380 13294
rect 11444 13230 11461 13294
rect 11525 13230 11542 13294
rect 11606 13230 11623 13294
rect 11687 13230 11704 13294
rect 11768 13230 11785 13294
rect 11849 13230 11866 13294
rect 11930 13230 11947 13294
rect 12011 13230 12028 13294
rect 12092 13230 12109 13294
rect 12173 13230 12190 13294
rect 12254 13230 12271 13294
rect 12335 13230 12352 13294
rect 12416 13230 12433 13294
rect 12497 13230 12514 13294
rect 12578 13230 12595 13294
rect 12659 13230 12676 13294
rect 12740 13230 12757 13294
rect 12821 13230 12838 13294
rect 12902 13230 12919 13294
rect 12983 13230 13000 13294
rect 13064 13230 13081 13294
rect 13145 13230 13162 13294
rect 13226 13230 13243 13294
rect 13307 13230 13324 13294
rect 13388 13230 13405 13294
rect 13469 13230 13486 13294
rect 13550 13230 13567 13294
rect 13631 13230 13648 13294
rect 13712 13230 13729 13294
rect 13793 13230 13810 13294
rect 13874 13230 13891 13294
rect 13955 13230 13972 13294
rect 14036 13230 14053 13294
rect 14117 13230 14134 13294
rect 14198 13230 14215 13294
rect 14279 13230 14296 13294
rect 14360 13230 14378 13294
rect 14442 13230 14460 13294
rect 14524 13230 14542 13294
rect 14606 13230 14624 13294
rect 14688 13230 14706 13294
rect 14770 13230 14788 13294
rect 14852 13230 15000 13294
rect 10083 13212 15000 13230
rect 10083 13148 10084 13212
rect 10148 13148 10165 13212
rect 10229 13148 10246 13212
rect 10310 13148 10327 13212
rect 10391 13148 10408 13212
rect 10472 13148 10489 13212
rect 10553 13148 10570 13212
rect 10634 13148 10651 13212
rect 10715 13148 10732 13212
rect 10796 13148 10813 13212
rect 10877 13148 10894 13212
rect 10958 13148 10975 13212
rect 11039 13148 11056 13212
rect 11120 13148 11137 13212
rect 11201 13148 11218 13212
rect 11282 13148 11299 13212
rect 11363 13148 11380 13212
rect 11444 13148 11461 13212
rect 11525 13148 11542 13212
rect 11606 13148 11623 13212
rect 11687 13148 11704 13212
rect 11768 13148 11785 13212
rect 11849 13148 11866 13212
rect 11930 13148 11947 13212
rect 12011 13148 12028 13212
rect 12092 13148 12109 13212
rect 12173 13148 12190 13212
rect 12254 13148 12271 13212
rect 12335 13148 12352 13212
rect 12416 13148 12433 13212
rect 12497 13148 12514 13212
rect 12578 13148 12595 13212
rect 12659 13148 12676 13212
rect 12740 13148 12757 13212
rect 12821 13148 12838 13212
rect 12902 13148 12919 13212
rect 12983 13148 13000 13212
rect 13064 13148 13081 13212
rect 13145 13148 13162 13212
rect 13226 13148 13243 13212
rect 13307 13148 13324 13212
rect 13388 13148 13405 13212
rect 13469 13148 13486 13212
rect 13550 13148 13567 13212
rect 13631 13148 13648 13212
rect 13712 13148 13729 13212
rect 13793 13148 13810 13212
rect 13874 13148 13891 13212
rect 13955 13148 13972 13212
rect 14036 13148 14053 13212
rect 14117 13148 14134 13212
rect 14198 13148 14215 13212
rect 14279 13148 14296 13212
rect 14360 13148 14378 13212
rect 14442 13148 14460 13212
rect 14524 13148 14542 13212
rect 14606 13148 14624 13212
rect 14688 13148 14706 13212
rect 14770 13148 14788 13212
rect 14852 13148 15000 13212
rect 10083 13130 15000 13148
rect 10083 13066 10084 13130
rect 10148 13066 10165 13130
rect 10229 13066 10246 13130
rect 10310 13066 10327 13130
rect 10391 13066 10408 13130
rect 10472 13066 10489 13130
rect 10553 13066 10570 13130
rect 10634 13066 10651 13130
rect 10715 13066 10732 13130
rect 10796 13066 10813 13130
rect 10877 13066 10894 13130
rect 10958 13066 10975 13130
rect 11039 13066 11056 13130
rect 11120 13066 11137 13130
rect 11201 13066 11218 13130
rect 11282 13066 11299 13130
rect 11363 13066 11380 13130
rect 11444 13066 11461 13130
rect 11525 13066 11542 13130
rect 11606 13066 11623 13130
rect 11687 13066 11704 13130
rect 11768 13066 11785 13130
rect 11849 13066 11866 13130
rect 11930 13066 11947 13130
rect 12011 13066 12028 13130
rect 12092 13066 12109 13130
rect 12173 13066 12190 13130
rect 12254 13066 12271 13130
rect 12335 13066 12352 13130
rect 12416 13066 12433 13130
rect 12497 13066 12514 13130
rect 12578 13066 12595 13130
rect 12659 13066 12676 13130
rect 12740 13066 12757 13130
rect 12821 13066 12838 13130
rect 12902 13066 12919 13130
rect 12983 13066 13000 13130
rect 13064 13066 13081 13130
rect 13145 13066 13162 13130
rect 13226 13066 13243 13130
rect 13307 13066 13324 13130
rect 13388 13066 13405 13130
rect 13469 13066 13486 13130
rect 13550 13066 13567 13130
rect 13631 13066 13648 13130
rect 13712 13066 13729 13130
rect 13793 13066 13810 13130
rect 13874 13066 13891 13130
rect 13955 13066 13972 13130
rect 14036 13066 14053 13130
rect 14117 13066 14134 13130
rect 14198 13066 14215 13130
rect 14279 13066 14296 13130
rect 14360 13066 14378 13130
rect 14442 13066 14460 13130
rect 14524 13066 14542 13130
rect 14606 13066 14624 13130
rect 14688 13066 14706 13130
rect 14770 13066 14788 13130
rect 14852 13066 15000 13130
rect 10083 13048 15000 13066
rect 10083 12984 10084 13048
rect 10148 12984 10165 13048
rect 10229 12984 10246 13048
rect 10310 12984 10327 13048
rect 10391 12984 10408 13048
rect 10472 12984 10489 13048
rect 10553 12984 10570 13048
rect 10634 12984 10651 13048
rect 10715 12984 10732 13048
rect 10796 12984 10813 13048
rect 10877 12984 10894 13048
rect 10958 12984 10975 13048
rect 11039 12984 11056 13048
rect 11120 12984 11137 13048
rect 11201 12984 11218 13048
rect 11282 12984 11299 13048
rect 11363 12984 11380 13048
rect 11444 12984 11461 13048
rect 11525 12984 11542 13048
rect 11606 12984 11623 13048
rect 11687 12984 11704 13048
rect 11768 12984 11785 13048
rect 11849 12984 11866 13048
rect 11930 12984 11947 13048
rect 12011 12984 12028 13048
rect 12092 12984 12109 13048
rect 12173 12984 12190 13048
rect 12254 12984 12271 13048
rect 12335 12984 12352 13048
rect 12416 12984 12433 13048
rect 12497 12984 12514 13048
rect 12578 12984 12595 13048
rect 12659 12984 12676 13048
rect 12740 12984 12757 13048
rect 12821 12984 12838 13048
rect 12902 12984 12919 13048
rect 12983 12984 13000 13048
rect 13064 12984 13081 13048
rect 13145 12984 13162 13048
rect 13226 12984 13243 13048
rect 13307 12984 13324 13048
rect 13388 12984 13405 13048
rect 13469 12984 13486 13048
rect 13550 12984 13567 13048
rect 13631 12984 13648 13048
rect 13712 12984 13729 13048
rect 13793 12984 13810 13048
rect 13874 12984 13891 13048
rect 13955 12984 13972 13048
rect 14036 12984 14053 13048
rect 14117 12984 14134 13048
rect 14198 12984 14215 13048
rect 14279 12984 14296 13048
rect 14360 12984 14378 13048
rect 14442 12984 14460 13048
rect 14524 12984 14542 13048
rect 14606 12984 14624 13048
rect 14688 12984 14706 13048
rect 14770 12984 14788 13048
rect 14852 12984 15000 13048
rect 10083 12966 15000 12984
rect 10083 12902 10084 12966
rect 10148 12902 10165 12966
rect 10229 12902 10246 12966
rect 10310 12902 10327 12966
rect 10391 12902 10408 12966
rect 10472 12902 10489 12966
rect 10553 12902 10570 12966
rect 10634 12902 10651 12966
rect 10715 12902 10732 12966
rect 10796 12902 10813 12966
rect 10877 12902 10894 12966
rect 10958 12902 10975 12966
rect 11039 12902 11056 12966
rect 11120 12902 11137 12966
rect 11201 12902 11218 12966
rect 11282 12902 11299 12966
rect 11363 12902 11380 12966
rect 11444 12902 11461 12966
rect 11525 12902 11542 12966
rect 11606 12902 11623 12966
rect 11687 12902 11704 12966
rect 11768 12902 11785 12966
rect 11849 12902 11866 12966
rect 11930 12902 11947 12966
rect 12011 12902 12028 12966
rect 12092 12902 12109 12966
rect 12173 12902 12190 12966
rect 12254 12902 12271 12966
rect 12335 12902 12352 12966
rect 12416 12902 12433 12966
rect 12497 12902 12514 12966
rect 12578 12902 12595 12966
rect 12659 12902 12676 12966
rect 12740 12902 12757 12966
rect 12821 12902 12838 12966
rect 12902 12902 12919 12966
rect 12983 12902 13000 12966
rect 13064 12902 13081 12966
rect 13145 12902 13162 12966
rect 13226 12902 13243 12966
rect 13307 12902 13324 12966
rect 13388 12902 13405 12966
rect 13469 12902 13486 12966
rect 13550 12902 13567 12966
rect 13631 12902 13648 12966
rect 13712 12902 13729 12966
rect 13793 12902 13810 12966
rect 13874 12902 13891 12966
rect 13955 12902 13972 12966
rect 14036 12902 14053 12966
rect 14117 12902 14134 12966
rect 14198 12902 14215 12966
rect 14279 12902 14296 12966
rect 14360 12902 14378 12966
rect 14442 12902 14460 12966
rect 14524 12902 14542 12966
rect 14606 12902 14624 12966
rect 14688 12902 14706 12966
rect 14770 12902 14788 12966
rect 14852 12902 15000 12966
rect 10083 12884 15000 12902
rect 10083 12820 10084 12884
rect 10148 12820 10165 12884
rect 10229 12820 10246 12884
rect 10310 12820 10327 12884
rect 10391 12820 10408 12884
rect 10472 12820 10489 12884
rect 10553 12820 10570 12884
rect 10634 12820 10651 12884
rect 10715 12820 10732 12884
rect 10796 12820 10813 12884
rect 10877 12820 10894 12884
rect 10958 12820 10975 12884
rect 11039 12820 11056 12884
rect 11120 12820 11137 12884
rect 11201 12820 11218 12884
rect 11282 12820 11299 12884
rect 11363 12820 11380 12884
rect 11444 12820 11461 12884
rect 11525 12820 11542 12884
rect 11606 12820 11623 12884
rect 11687 12820 11704 12884
rect 11768 12820 11785 12884
rect 11849 12820 11866 12884
rect 11930 12820 11947 12884
rect 12011 12820 12028 12884
rect 12092 12820 12109 12884
rect 12173 12820 12190 12884
rect 12254 12820 12271 12884
rect 12335 12820 12352 12884
rect 12416 12820 12433 12884
rect 12497 12820 12514 12884
rect 12578 12820 12595 12884
rect 12659 12820 12676 12884
rect 12740 12820 12757 12884
rect 12821 12820 12838 12884
rect 12902 12820 12919 12884
rect 12983 12820 13000 12884
rect 13064 12820 13081 12884
rect 13145 12820 13162 12884
rect 13226 12820 13243 12884
rect 13307 12820 13324 12884
rect 13388 12820 13405 12884
rect 13469 12820 13486 12884
rect 13550 12820 13567 12884
rect 13631 12820 13648 12884
rect 13712 12820 13729 12884
rect 13793 12820 13810 12884
rect 13874 12820 13891 12884
rect 13955 12820 13972 12884
rect 14036 12820 14053 12884
rect 14117 12820 14134 12884
rect 14198 12820 14215 12884
rect 14279 12820 14296 12884
rect 14360 12820 14378 12884
rect 14442 12820 14460 12884
rect 14524 12820 14542 12884
rect 14606 12820 14624 12884
rect 14688 12820 14706 12884
rect 14770 12820 14788 12884
rect 14852 12820 15000 12884
rect 10083 12817 15000 12820
rect 0 11647 254 12537
rect 14746 11647 15000 12537
rect 0 11281 254 11347
rect 14746 11281 15000 11347
rect 0 10625 254 11221
rect 14746 10625 15000 11221
rect 0 10329 254 10565
rect 14746 10329 15000 10565
rect 0 9673 254 10269
rect 14746 9673 15000 10269
rect 0 9547 254 9613
rect 14746 9547 15000 9613
rect 0 8317 254 9247
rect 14746 8317 15000 9247
rect 0 7347 254 8037
rect 14746 7347 15000 8037
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 5167 254 6097
rect 14746 5167 15000 6097
rect 0 4884 4874 4887
rect 0 4820 105 4884
rect 169 4820 186 4884
rect 250 4820 267 4884
rect 331 4820 348 4884
rect 412 4820 429 4884
rect 493 4820 510 4884
rect 574 4820 591 4884
rect 655 4820 672 4884
rect 736 4820 753 4884
rect 817 4820 834 4884
rect 898 4820 915 4884
rect 979 4820 996 4884
rect 1060 4820 1077 4884
rect 1141 4820 1158 4884
rect 1222 4820 1239 4884
rect 1303 4820 1320 4884
rect 1384 4820 1401 4884
rect 1465 4820 1482 4884
rect 1546 4820 1563 4884
rect 1627 4820 1644 4884
rect 1708 4820 1725 4884
rect 1789 4820 1806 4884
rect 1870 4820 1887 4884
rect 1951 4820 1968 4884
rect 2032 4820 2049 4884
rect 2113 4820 2130 4884
rect 2194 4820 2211 4884
rect 2275 4820 2292 4884
rect 2356 4820 2373 4884
rect 2437 4820 2454 4884
rect 2518 4820 2535 4884
rect 2599 4820 2616 4884
rect 2680 4820 2697 4884
rect 2761 4820 2778 4884
rect 2842 4820 2859 4884
rect 2923 4820 2940 4884
rect 3004 4820 3021 4884
rect 3085 4820 3102 4884
rect 3166 4820 3183 4884
rect 3247 4820 3264 4884
rect 3328 4820 3345 4884
rect 3409 4820 3426 4884
rect 3490 4820 3507 4884
rect 3571 4820 3588 4884
rect 3652 4820 3669 4884
rect 3733 4820 3750 4884
rect 3814 4820 3831 4884
rect 3895 4820 3912 4884
rect 3976 4820 3993 4884
rect 4057 4820 4074 4884
rect 4138 4820 4155 4884
rect 4219 4820 4236 4884
rect 4300 4820 4317 4884
rect 4381 4820 4399 4884
rect 4463 4820 4481 4884
rect 4545 4820 4563 4884
rect 4627 4820 4645 4884
rect 4709 4820 4727 4884
rect 4791 4820 4809 4884
rect 4873 4820 4874 4884
rect 0 4798 4874 4820
rect 0 4734 105 4798
rect 169 4734 186 4798
rect 250 4734 267 4798
rect 331 4734 348 4798
rect 412 4734 429 4798
rect 493 4734 510 4798
rect 574 4734 591 4798
rect 655 4734 672 4798
rect 736 4734 753 4798
rect 817 4734 834 4798
rect 898 4734 915 4798
rect 979 4734 996 4798
rect 1060 4734 1077 4798
rect 1141 4734 1158 4798
rect 1222 4734 1239 4798
rect 1303 4734 1320 4798
rect 1384 4734 1401 4798
rect 1465 4734 1482 4798
rect 1546 4734 1563 4798
rect 1627 4734 1644 4798
rect 1708 4734 1725 4798
rect 1789 4734 1806 4798
rect 1870 4734 1887 4798
rect 1951 4734 1968 4798
rect 2032 4734 2049 4798
rect 2113 4734 2130 4798
rect 2194 4734 2211 4798
rect 2275 4734 2292 4798
rect 2356 4734 2373 4798
rect 2437 4734 2454 4798
rect 2518 4734 2535 4798
rect 2599 4734 2616 4798
rect 2680 4734 2697 4798
rect 2761 4734 2778 4798
rect 2842 4734 2859 4798
rect 2923 4734 2940 4798
rect 3004 4734 3021 4798
rect 3085 4734 3102 4798
rect 3166 4734 3183 4798
rect 3247 4734 3264 4798
rect 3328 4734 3345 4798
rect 3409 4734 3426 4798
rect 3490 4734 3507 4798
rect 3571 4734 3588 4798
rect 3652 4734 3669 4798
rect 3733 4734 3750 4798
rect 3814 4734 3831 4798
rect 3895 4734 3912 4798
rect 3976 4734 3993 4798
rect 4057 4734 4074 4798
rect 4138 4734 4155 4798
rect 4219 4734 4236 4798
rect 4300 4734 4317 4798
rect 4381 4734 4399 4798
rect 4463 4734 4481 4798
rect 4545 4734 4563 4798
rect 4627 4734 4645 4798
rect 4709 4734 4727 4798
rect 4791 4734 4809 4798
rect 4873 4734 4874 4798
rect 0 4712 4874 4734
rect 0 4648 105 4712
rect 169 4648 186 4712
rect 250 4648 267 4712
rect 331 4648 348 4712
rect 412 4648 429 4712
rect 493 4648 510 4712
rect 574 4648 591 4712
rect 655 4648 672 4712
rect 736 4648 753 4712
rect 817 4648 834 4712
rect 898 4648 915 4712
rect 979 4648 996 4712
rect 1060 4648 1077 4712
rect 1141 4648 1158 4712
rect 1222 4648 1239 4712
rect 1303 4648 1320 4712
rect 1384 4648 1401 4712
rect 1465 4648 1482 4712
rect 1546 4648 1563 4712
rect 1627 4648 1644 4712
rect 1708 4648 1725 4712
rect 1789 4648 1806 4712
rect 1870 4648 1887 4712
rect 1951 4648 1968 4712
rect 2032 4648 2049 4712
rect 2113 4648 2130 4712
rect 2194 4648 2211 4712
rect 2275 4648 2292 4712
rect 2356 4648 2373 4712
rect 2437 4648 2454 4712
rect 2518 4648 2535 4712
rect 2599 4648 2616 4712
rect 2680 4648 2697 4712
rect 2761 4648 2778 4712
rect 2842 4648 2859 4712
rect 2923 4648 2940 4712
rect 3004 4648 3021 4712
rect 3085 4648 3102 4712
rect 3166 4648 3183 4712
rect 3247 4648 3264 4712
rect 3328 4648 3345 4712
rect 3409 4648 3426 4712
rect 3490 4648 3507 4712
rect 3571 4648 3588 4712
rect 3652 4648 3669 4712
rect 3733 4648 3750 4712
rect 3814 4648 3831 4712
rect 3895 4648 3912 4712
rect 3976 4648 3993 4712
rect 4057 4648 4074 4712
rect 4138 4648 4155 4712
rect 4219 4648 4236 4712
rect 4300 4648 4317 4712
rect 4381 4648 4399 4712
rect 4463 4648 4481 4712
rect 4545 4648 4563 4712
rect 4627 4648 4645 4712
rect 4709 4648 4727 4712
rect 4791 4648 4809 4712
rect 4873 4648 4874 4712
rect 0 4626 4874 4648
rect 0 4562 105 4626
rect 169 4562 186 4626
rect 250 4562 267 4626
rect 331 4562 348 4626
rect 412 4562 429 4626
rect 493 4562 510 4626
rect 574 4562 591 4626
rect 655 4562 672 4626
rect 736 4562 753 4626
rect 817 4562 834 4626
rect 898 4562 915 4626
rect 979 4562 996 4626
rect 1060 4562 1077 4626
rect 1141 4562 1158 4626
rect 1222 4562 1239 4626
rect 1303 4562 1320 4626
rect 1384 4562 1401 4626
rect 1465 4562 1482 4626
rect 1546 4562 1563 4626
rect 1627 4562 1644 4626
rect 1708 4562 1725 4626
rect 1789 4562 1806 4626
rect 1870 4562 1887 4626
rect 1951 4562 1968 4626
rect 2032 4562 2049 4626
rect 2113 4562 2130 4626
rect 2194 4562 2211 4626
rect 2275 4562 2292 4626
rect 2356 4562 2373 4626
rect 2437 4562 2454 4626
rect 2518 4562 2535 4626
rect 2599 4562 2616 4626
rect 2680 4562 2697 4626
rect 2761 4562 2778 4626
rect 2842 4562 2859 4626
rect 2923 4562 2940 4626
rect 3004 4562 3021 4626
rect 3085 4562 3102 4626
rect 3166 4562 3183 4626
rect 3247 4562 3264 4626
rect 3328 4562 3345 4626
rect 3409 4562 3426 4626
rect 3490 4562 3507 4626
rect 3571 4562 3588 4626
rect 3652 4562 3669 4626
rect 3733 4562 3750 4626
rect 3814 4562 3831 4626
rect 3895 4562 3912 4626
rect 3976 4562 3993 4626
rect 4057 4562 4074 4626
rect 4138 4562 4155 4626
rect 4219 4562 4236 4626
rect 4300 4562 4317 4626
rect 4381 4562 4399 4626
rect 4463 4562 4481 4626
rect 4545 4562 4563 4626
rect 4627 4562 4645 4626
rect 4709 4562 4727 4626
rect 4791 4562 4809 4626
rect 4873 4562 4874 4626
rect 0 4540 4874 4562
rect 0 4476 105 4540
rect 169 4476 186 4540
rect 250 4476 267 4540
rect 331 4476 348 4540
rect 412 4476 429 4540
rect 493 4476 510 4540
rect 574 4476 591 4540
rect 655 4476 672 4540
rect 736 4476 753 4540
rect 817 4476 834 4540
rect 898 4476 915 4540
rect 979 4476 996 4540
rect 1060 4476 1077 4540
rect 1141 4476 1158 4540
rect 1222 4476 1239 4540
rect 1303 4476 1320 4540
rect 1384 4476 1401 4540
rect 1465 4476 1482 4540
rect 1546 4476 1563 4540
rect 1627 4476 1644 4540
rect 1708 4476 1725 4540
rect 1789 4476 1806 4540
rect 1870 4476 1887 4540
rect 1951 4476 1968 4540
rect 2032 4476 2049 4540
rect 2113 4476 2130 4540
rect 2194 4476 2211 4540
rect 2275 4476 2292 4540
rect 2356 4476 2373 4540
rect 2437 4476 2454 4540
rect 2518 4476 2535 4540
rect 2599 4476 2616 4540
rect 2680 4476 2697 4540
rect 2761 4476 2778 4540
rect 2842 4476 2859 4540
rect 2923 4476 2940 4540
rect 3004 4476 3021 4540
rect 3085 4476 3102 4540
rect 3166 4476 3183 4540
rect 3247 4476 3264 4540
rect 3328 4476 3345 4540
rect 3409 4476 3426 4540
rect 3490 4476 3507 4540
rect 3571 4476 3588 4540
rect 3652 4476 3669 4540
rect 3733 4476 3750 4540
rect 3814 4476 3831 4540
rect 3895 4476 3912 4540
rect 3976 4476 3993 4540
rect 4057 4476 4074 4540
rect 4138 4476 4155 4540
rect 4219 4476 4236 4540
rect 4300 4476 4317 4540
rect 4381 4476 4399 4540
rect 4463 4476 4481 4540
rect 4545 4476 4563 4540
rect 4627 4476 4645 4540
rect 4709 4476 4727 4540
rect 4791 4476 4809 4540
rect 4873 4476 4874 4540
rect 0 4454 4874 4476
rect 0 4390 105 4454
rect 169 4390 186 4454
rect 250 4390 267 4454
rect 331 4390 348 4454
rect 412 4390 429 4454
rect 493 4390 510 4454
rect 574 4390 591 4454
rect 655 4390 672 4454
rect 736 4390 753 4454
rect 817 4390 834 4454
rect 898 4390 915 4454
rect 979 4390 996 4454
rect 1060 4390 1077 4454
rect 1141 4390 1158 4454
rect 1222 4390 1239 4454
rect 1303 4390 1320 4454
rect 1384 4390 1401 4454
rect 1465 4390 1482 4454
rect 1546 4390 1563 4454
rect 1627 4390 1644 4454
rect 1708 4390 1725 4454
rect 1789 4390 1806 4454
rect 1870 4390 1887 4454
rect 1951 4390 1968 4454
rect 2032 4390 2049 4454
rect 2113 4390 2130 4454
rect 2194 4390 2211 4454
rect 2275 4390 2292 4454
rect 2356 4390 2373 4454
rect 2437 4390 2454 4454
rect 2518 4390 2535 4454
rect 2599 4390 2616 4454
rect 2680 4390 2697 4454
rect 2761 4390 2778 4454
rect 2842 4390 2859 4454
rect 2923 4390 2940 4454
rect 3004 4390 3021 4454
rect 3085 4390 3102 4454
rect 3166 4390 3183 4454
rect 3247 4390 3264 4454
rect 3328 4390 3345 4454
rect 3409 4390 3426 4454
rect 3490 4390 3507 4454
rect 3571 4390 3588 4454
rect 3652 4390 3669 4454
rect 3733 4390 3750 4454
rect 3814 4390 3831 4454
rect 3895 4390 3912 4454
rect 3976 4390 3993 4454
rect 4057 4390 4074 4454
rect 4138 4390 4155 4454
rect 4219 4390 4236 4454
rect 4300 4390 4317 4454
rect 4381 4390 4399 4454
rect 4463 4390 4481 4454
rect 4545 4390 4563 4454
rect 4627 4390 4645 4454
rect 4709 4390 4727 4454
rect 4791 4390 4809 4454
rect 4873 4390 4874 4454
rect 0 4368 4874 4390
rect 0 4304 105 4368
rect 169 4304 186 4368
rect 250 4304 267 4368
rect 331 4304 348 4368
rect 412 4304 429 4368
rect 493 4304 510 4368
rect 574 4304 591 4368
rect 655 4304 672 4368
rect 736 4304 753 4368
rect 817 4304 834 4368
rect 898 4304 915 4368
rect 979 4304 996 4368
rect 1060 4304 1077 4368
rect 1141 4304 1158 4368
rect 1222 4304 1239 4368
rect 1303 4304 1320 4368
rect 1384 4304 1401 4368
rect 1465 4304 1482 4368
rect 1546 4304 1563 4368
rect 1627 4304 1644 4368
rect 1708 4304 1725 4368
rect 1789 4304 1806 4368
rect 1870 4304 1887 4368
rect 1951 4304 1968 4368
rect 2032 4304 2049 4368
rect 2113 4304 2130 4368
rect 2194 4304 2211 4368
rect 2275 4304 2292 4368
rect 2356 4304 2373 4368
rect 2437 4304 2454 4368
rect 2518 4304 2535 4368
rect 2599 4304 2616 4368
rect 2680 4304 2697 4368
rect 2761 4304 2778 4368
rect 2842 4304 2859 4368
rect 2923 4304 2940 4368
rect 3004 4304 3021 4368
rect 3085 4304 3102 4368
rect 3166 4304 3183 4368
rect 3247 4304 3264 4368
rect 3328 4304 3345 4368
rect 3409 4304 3426 4368
rect 3490 4304 3507 4368
rect 3571 4304 3588 4368
rect 3652 4304 3669 4368
rect 3733 4304 3750 4368
rect 3814 4304 3831 4368
rect 3895 4304 3912 4368
rect 3976 4304 3993 4368
rect 4057 4304 4074 4368
rect 4138 4304 4155 4368
rect 4219 4304 4236 4368
rect 4300 4304 4317 4368
rect 4381 4304 4399 4368
rect 4463 4304 4481 4368
rect 4545 4304 4563 4368
rect 4627 4304 4645 4368
rect 4709 4304 4727 4368
rect 4791 4304 4809 4368
rect 4873 4304 4874 4368
rect 0 4282 4874 4304
rect 0 4218 105 4282
rect 169 4218 186 4282
rect 250 4218 267 4282
rect 331 4218 348 4282
rect 412 4218 429 4282
rect 493 4218 510 4282
rect 574 4218 591 4282
rect 655 4218 672 4282
rect 736 4218 753 4282
rect 817 4218 834 4282
rect 898 4218 915 4282
rect 979 4218 996 4282
rect 1060 4218 1077 4282
rect 1141 4218 1158 4282
rect 1222 4218 1239 4282
rect 1303 4218 1320 4282
rect 1384 4218 1401 4282
rect 1465 4218 1482 4282
rect 1546 4218 1563 4282
rect 1627 4218 1644 4282
rect 1708 4218 1725 4282
rect 1789 4218 1806 4282
rect 1870 4218 1887 4282
rect 1951 4218 1968 4282
rect 2032 4218 2049 4282
rect 2113 4218 2130 4282
rect 2194 4218 2211 4282
rect 2275 4218 2292 4282
rect 2356 4218 2373 4282
rect 2437 4218 2454 4282
rect 2518 4218 2535 4282
rect 2599 4218 2616 4282
rect 2680 4218 2697 4282
rect 2761 4218 2778 4282
rect 2842 4218 2859 4282
rect 2923 4218 2940 4282
rect 3004 4218 3021 4282
rect 3085 4218 3102 4282
rect 3166 4218 3183 4282
rect 3247 4218 3264 4282
rect 3328 4218 3345 4282
rect 3409 4218 3426 4282
rect 3490 4218 3507 4282
rect 3571 4218 3588 4282
rect 3652 4218 3669 4282
rect 3733 4218 3750 4282
rect 3814 4218 3831 4282
rect 3895 4218 3912 4282
rect 3976 4218 3993 4282
rect 4057 4218 4074 4282
rect 4138 4218 4155 4282
rect 4219 4218 4236 4282
rect 4300 4218 4317 4282
rect 4381 4218 4399 4282
rect 4463 4218 4481 4282
rect 4545 4218 4563 4282
rect 4627 4218 4645 4282
rect 4709 4218 4727 4282
rect 4791 4218 4809 4282
rect 4873 4218 4874 4282
rect 0 4196 4874 4218
rect 0 4132 105 4196
rect 169 4132 186 4196
rect 250 4132 267 4196
rect 331 4132 348 4196
rect 412 4132 429 4196
rect 493 4132 510 4196
rect 574 4132 591 4196
rect 655 4132 672 4196
rect 736 4132 753 4196
rect 817 4132 834 4196
rect 898 4132 915 4196
rect 979 4132 996 4196
rect 1060 4132 1077 4196
rect 1141 4132 1158 4196
rect 1222 4132 1239 4196
rect 1303 4132 1320 4196
rect 1384 4132 1401 4196
rect 1465 4132 1482 4196
rect 1546 4132 1563 4196
rect 1627 4132 1644 4196
rect 1708 4132 1725 4196
rect 1789 4132 1806 4196
rect 1870 4132 1887 4196
rect 1951 4132 1968 4196
rect 2032 4132 2049 4196
rect 2113 4132 2130 4196
rect 2194 4132 2211 4196
rect 2275 4132 2292 4196
rect 2356 4132 2373 4196
rect 2437 4132 2454 4196
rect 2518 4132 2535 4196
rect 2599 4132 2616 4196
rect 2680 4132 2697 4196
rect 2761 4132 2778 4196
rect 2842 4132 2859 4196
rect 2923 4132 2940 4196
rect 3004 4132 3021 4196
rect 3085 4132 3102 4196
rect 3166 4132 3183 4196
rect 3247 4132 3264 4196
rect 3328 4132 3345 4196
rect 3409 4132 3426 4196
rect 3490 4132 3507 4196
rect 3571 4132 3588 4196
rect 3652 4132 3669 4196
rect 3733 4132 3750 4196
rect 3814 4132 3831 4196
rect 3895 4132 3912 4196
rect 3976 4132 3993 4196
rect 4057 4132 4074 4196
rect 4138 4132 4155 4196
rect 4219 4132 4236 4196
rect 4300 4132 4317 4196
rect 4381 4132 4399 4196
rect 4463 4132 4481 4196
rect 4545 4132 4563 4196
rect 4627 4132 4645 4196
rect 4709 4132 4727 4196
rect 4791 4132 4809 4196
rect 4873 4132 4874 4196
rect 0 4110 4874 4132
rect 0 4046 105 4110
rect 169 4046 186 4110
rect 250 4046 267 4110
rect 331 4046 348 4110
rect 412 4046 429 4110
rect 493 4046 510 4110
rect 574 4046 591 4110
rect 655 4046 672 4110
rect 736 4046 753 4110
rect 817 4046 834 4110
rect 898 4046 915 4110
rect 979 4046 996 4110
rect 1060 4046 1077 4110
rect 1141 4046 1158 4110
rect 1222 4046 1239 4110
rect 1303 4046 1320 4110
rect 1384 4046 1401 4110
rect 1465 4046 1482 4110
rect 1546 4046 1563 4110
rect 1627 4046 1644 4110
rect 1708 4046 1725 4110
rect 1789 4046 1806 4110
rect 1870 4046 1887 4110
rect 1951 4046 1968 4110
rect 2032 4046 2049 4110
rect 2113 4046 2130 4110
rect 2194 4046 2211 4110
rect 2275 4046 2292 4110
rect 2356 4046 2373 4110
rect 2437 4046 2454 4110
rect 2518 4046 2535 4110
rect 2599 4046 2616 4110
rect 2680 4046 2697 4110
rect 2761 4046 2778 4110
rect 2842 4046 2859 4110
rect 2923 4046 2940 4110
rect 3004 4046 3021 4110
rect 3085 4046 3102 4110
rect 3166 4046 3183 4110
rect 3247 4046 3264 4110
rect 3328 4046 3345 4110
rect 3409 4046 3426 4110
rect 3490 4046 3507 4110
rect 3571 4046 3588 4110
rect 3652 4046 3669 4110
rect 3733 4046 3750 4110
rect 3814 4046 3831 4110
rect 3895 4046 3912 4110
rect 3976 4046 3993 4110
rect 4057 4046 4074 4110
rect 4138 4046 4155 4110
rect 4219 4046 4236 4110
rect 4300 4046 4317 4110
rect 4381 4046 4399 4110
rect 4463 4046 4481 4110
rect 4545 4046 4563 4110
rect 4627 4046 4645 4110
rect 4709 4046 4727 4110
rect 4791 4046 4809 4110
rect 4873 4046 4874 4110
rect 0 4024 4874 4046
rect 0 3960 105 4024
rect 169 3960 186 4024
rect 250 3960 267 4024
rect 331 3960 348 4024
rect 412 3960 429 4024
rect 493 3960 510 4024
rect 574 3960 591 4024
rect 655 3960 672 4024
rect 736 3960 753 4024
rect 817 3960 834 4024
rect 898 3960 915 4024
rect 979 3960 996 4024
rect 1060 3960 1077 4024
rect 1141 3960 1158 4024
rect 1222 3960 1239 4024
rect 1303 3960 1320 4024
rect 1384 3960 1401 4024
rect 1465 3960 1482 4024
rect 1546 3960 1563 4024
rect 1627 3960 1644 4024
rect 1708 3960 1725 4024
rect 1789 3960 1806 4024
rect 1870 3960 1887 4024
rect 1951 3960 1968 4024
rect 2032 3960 2049 4024
rect 2113 3960 2130 4024
rect 2194 3960 2211 4024
rect 2275 3960 2292 4024
rect 2356 3960 2373 4024
rect 2437 3960 2454 4024
rect 2518 3960 2535 4024
rect 2599 3960 2616 4024
rect 2680 3960 2697 4024
rect 2761 3960 2778 4024
rect 2842 3960 2859 4024
rect 2923 3960 2940 4024
rect 3004 3960 3021 4024
rect 3085 3960 3102 4024
rect 3166 3960 3183 4024
rect 3247 3960 3264 4024
rect 3328 3960 3345 4024
rect 3409 3960 3426 4024
rect 3490 3960 3507 4024
rect 3571 3960 3588 4024
rect 3652 3960 3669 4024
rect 3733 3960 3750 4024
rect 3814 3960 3831 4024
rect 3895 3960 3912 4024
rect 3976 3960 3993 4024
rect 4057 3960 4074 4024
rect 4138 3960 4155 4024
rect 4219 3960 4236 4024
rect 4300 3960 4317 4024
rect 4381 3960 4399 4024
rect 4463 3960 4481 4024
rect 4545 3960 4563 4024
rect 4627 3960 4645 4024
rect 4709 3960 4727 4024
rect 4791 3960 4809 4024
rect 4873 3960 4874 4024
rect 0 3957 4874 3960
rect 10083 4884 15000 4887
rect 10083 4820 10084 4884
rect 10148 4820 10165 4884
rect 10229 4820 10246 4884
rect 10310 4820 10327 4884
rect 10391 4820 10408 4884
rect 10472 4820 10489 4884
rect 10553 4820 10570 4884
rect 10634 4820 10651 4884
rect 10715 4820 10732 4884
rect 10796 4820 10813 4884
rect 10877 4820 10894 4884
rect 10958 4820 10975 4884
rect 11039 4820 11056 4884
rect 11120 4820 11137 4884
rect 11201 4820 11218 4884
rect 11282 4820 11299 4884
rect 11363 4820 11380 4884
rect 11444 4820 11461 4884
rect 11525 4820 11542 4884
rect 11606 4820 11623 4884
rect 11687 4820 11704 4884
rect 11768 4820 11785 4884
rect 11849 4820 11866 4884
rect 11930 4820 11947 4884
rect 12011 4820 12028 4884
rect 12092 4820 12109 4884
rect 12173 4820 12190 4884
rect 12254 4820 12271 4884
rect 12335 4820 12352 4884
rect 12416 4820 12433 4884
rect 12497 4820 12514 4884
rect 12578 4820 12595 4884
rect 12659 4820 12676 4884
rect 12740 4820 12757 4884
rect 12821 4820 12838 4884
rect 12902 4820 12919 4884
rect 12983 4820 13000 4884
rect 13064 4820 13081 4884
rect 13145 4820 13162 4884
rect 13226 4820 13243 4884
rect 13307 4820 13324 4884
rect 13388 4820 13405 4884
rect 13469 4820 13486 4884
rect 13550 4820 13567 4884
rect 13631 4820 13648 4884
rect 13712 4820 13729 4884
rect 13793 4820 13810 4884
rect 13874 4820 13891 4884
rect 13955 4820 13972 4884
rect 14036 4820 14053 4884
rect 14117 4820 14134 4884
rect 14198 4820 14215 4884
rect 14279 4820 14296 4884
rect 14360 4820 14378 4884
rect 14442 4820 14460 4884
rect 14524 4820 14542 4884
rect 14606 4820 14624 4884
rect 14688 4820 14706 4884
rect 14770 4820 14788 4884
rect 14852 4820 15000 4884
rect 10083 4798 15000 4820
rect 10083 4734 10084 4798
rect 10148 4734 10165 4798
rect 10229 4734 10246 4798
rect 10310 4734 10327 4798
rect 10391 4734 10408 4798
rect 10472 4734 10489 4798
rect 10553 4734 10570 4798
rect 10634 4734 10651 4798
rect 10715 4734 10732 4798
rect 10796 4734 10813 4798
rect 10877 4734 10894 4798
rect 10958 4734 10975 4798
rect 11039 4734 11056 4798
rect 11120 4734 11137 4798
rect 11201 4734 11218 4798
rect 11282 4734 11299 4798
rect 11363 4734 11380 4798
rect 11444 4734 11461 4798
rect 11525 4734 11542 4798
rect 11606 4734 11623 4798
rect 11687 4734 11704 4798
rect 11768 4734 11785 4798
rect 11849 4734 11866 4798
rect 11930 4734 11947 4798
rect 12011 4734 12028 4798
rect 12092 4734 12109 4798
rect 12173 4734 12190 4798
rect 12254 4734 12271 4798
rect 12335 4734 12352 4798
rect 12416 4734 12433 4798
rect 12497 4734 12514 4798
rect 12578 4734 12595 4798
rect 12659 4734 12676 4798
rect 12740 4734 12757 4798
rect 12821 4734 12838 4798
rect 12902 4734 12919 4798
rect 12983 4734 13000 4798
rect 13064 4734 13081 4798
rect 13145 4734 13162 4798
rect 13226 4734 13243 4798
rect 13307 4734 13324 4798
rect 13388 4734 13405 4798
rect 13469 4734 13486 4798
rect 13550 4734 13567 4798
rect 13631 4734 13648 4798
rect 13712 4734 13729 4798
rect 13793 4734 13810 4798
rect 13874 4734 13891 4798
rect 13955 4734 13972 4798
rect 14036 4734 14053 4798
rect 14117 4734 14134 4798
rect 14198 4734 14215 4798
rect 14279 4734 14296 4798
rect 14360 4734 14378 4798
rect 14442 4734 14460 4798
rect 14524 4734 14542 4798
rect 14606 4734 14624 4798
rect 14688 4734 14706 4798
rect 14770 4734 14788 4798
rect 14852 4734 15000 4798
rect 10083 4712 15000 4734
rect 10083 4648 10084 4712
rect 10148 4648 10165 4712
rect 10229 4648 10246 4712
rect 10310 4648 10327 4712
rect 10391 4648 10408 4712
rect 10472 4648 10489 4712
rect 10553 4648 10570 4712
rect 10634 4648 10651 4712
rect 10715 4648 10732 4712
rect 10796 4648 10813 4712
rect 10877 4648 10894 4712
rect 10958 4648 10975 4712
rect 11039 4648 11056 4712
rect 11120 4648 11137 4712
rect 11201 4648 11218 4712
rect 11282 4648 11299 4712
rect 11363 4648 11380 4712
rect 11444 4648 11461 4712
rect 11525 4648 11542 4712
rect 11606 4648 11623 4712
rect 11687 4648 11704 4712
rect 11768 4648 11785 4712
rect 11849 4648 11866 4712
rect 11930 4648 11947 4712
rect 12011 4648 12028 4712
rect 12092 4648 12109 4712
rect 12173 4648 12190 4712
rect 12254 4648 12271 4712
rect 12335 4648 12352 4712
rect 12416 4648 12433 4712
rect 12497 4648 12514 4712
rect 12578 4648 12595 4712
rect 12659 4648 12676 4712
rect 12740 4648 12757 4712
rect 12821 4648 12838 4712
rect 12902 4648 12919 4712
rect 12983 4648 13000 4712
rect 13064 4648 13081 4712
rect 13145 4648 13162 4712
rect 13226 4648 13243 4712
rect 13307 4648 13324 4712
rect 13388 4648 13405 4712
rect 13469 4648 13486 4712
rect 13550 4648 13567 4712
rect 13631 4648 13648 4712
rect 13712 4648 13729 4712
rect 13793 4648 13810 4712
rect 13874 4648 13891 4712
rect 13955 4648 13972 4712
rect 14036 4648 14053 4712
rect 14117 4648 14134 4712
rect 14198 4648 14215 4712
rect 14279 4648 14296 4712
rect 14360 4648 14378 4712
rect 14442 4648 14460 4712
rect 14524 4648 14542 4712
rect 14606 4648 14624 4712
rect 14688 4648 14706 4712
rect 14770 4648 14788 4712
rect 14852 4648 15000 4712
rect 10083 4626 15000 4648
rect 10083 4562 10084 4626
rect 10148 4562 10165 4626
rect 10229 4562 10246 4626
rect 10310 4562 10327 4626
rect 10391 4562 10408 4626
rect 10472 4562 10489 4626
rect 10553 4562 10570 4626
rect 10634 4562 10651 4626
rect 10715 4562 10732 4626
rect 10796 4562 10813 4626
rect 10877 4562 10894 4626
rect 10958 4562 10975 4626
rect 11039 4562 11056 4626
rect 11120 4562 11137 4626
rect 11201 4562 11218 4626
rect 11282 4562 11299 4626
rect 11363 4562 11380 4626
rect 11444 4562 11461 4626
rect 11525 4562 11542 4626
rect 11606 4562 11623 4626
rect 11687 4562 11704 4626
rect 11768 4562 11785 4626
rect 11849 4562 11866 4626
rect 11930 4562 11947 4626
rect 12011 4562 12028 4626
rect 12092 4562 12109 4626
rect 12173 4562 12190 4626
rect 12254 4562 12271 4626
rect 12335 4562 12352 4626
rect 12416 4562 12433 4626
rect 12497 4562 12514 4626
rect 12578 4562 12595 4626
rect 12659 4562 12676 4626
rect 12740 4562 12757 4626
rect 12821 4562 12838 4626
rect 12902 4562 12919 4626
rect 12983 4562 13000 4626
rect 13064 4562 13081 4626
rect 13145 4562 13162 4626
rect 13226 4562 13243 4626
rect 13307 4562 13324 4626
rect 13388 4562 13405 4626
rect 13469 4562 13486 4626
rect 13550 4562 13567 4626
rect 13631 4562 13648 4626
rect 13712 4562 13729 4626
rect 13793 4562 13810 4626
rect 13874 4562 13891 4626
rect 13955 4562 13972 4626
rect 14036 4562 14053 4626
rect 14117 4562 14134 4626
rect 14198 4562 14215 4626
rect 14279 4562 14296 4626
rect 14360 4562 14378 4626
rect 14442 4562 14460 4626
rect 14524 4562 14542 4626
rect 14606 4562 14624 4626
rect 14688 4562 14706 4626
rect 14770 4562 14788 4626
rect 14852 4562 15000 4626
rect 10083 4540 15000 4562
rect 10083 4476 10084 4540
rect 10148 4476 10165 4540
rect 10229 4476 10246 4540
rect 10310 4476 10327 4540
rect 10391 4476 10408 4540
rect 10472 4476 10489 4540
rect 10553 4476 10570 4540
rect 10634 4476 10651 4540
rect 10715 4476 10732 4540
rect 10796 4476 10813 4540
rect 10877 4476 10894 4540
rect 10958 4476 10975 4540
rect 11039 4476 11056 4540
rect 11120 4476 11137 4540
rect 11201 4476 11218 4540
rect 11282 4476 11299 4540
rect 11363 4476 11380 4540
rect 11444 4476 11461 4540
rect 11525 4476 11542 4540
rect 11606 4476 11623 4540
rect 11687 4476 11704 4540
rect 11768 4476 11785 4540
rect 11849 4476 11866 4540
rect 11930 4476 11947 4540
rect 12011 4476 12028 4540
rect 12092 4476 12109 4540
rect 12173 4476 12190 4540
rect 12254 4476 12271 4540
rect 12335 4476 12352 4540
rect 12416 4476 12433 4540
rect 12497 4476 12514 4540
rect 12578 4476 12595 4540
rect 12659 4476 12676 4540
rect 12740 4476 12757 4540
rect 12821 4476 12838 4540
rect 12902 4476 12919 4540
rect 12983 4476 13000 4540
rect 13064 4476 13081 4540
rect 13145 4476 13162 4540
rect 13226 4476 13243 4540
rect 13307 4476 13324 4540
rect 13388 4476 13405 4540
rect 13469 4476 13486 4540
rect 13550 4476 13567 4540
rect 13631 4476 13648 4540
rect 13712 4476 13729 4540
rect 13793 4476 13810 4540
rect 13874 4476 13891 4540
rect 13955 4476 13972 4540
rect 14036 4476 14053 4540
rect 14117 4476 14134 4540
rect 14198 4476 14215 4540
rect 14279 4476 14296 4540
rect 14360 4476 14378 4540
rect 14442 4476 14460 4540
rect 14524 4476 14542 4540
rect 14606 4476 14624 4540
rect 14688 4476 14706 4540
rect 14770 4476 14788 4540
rect 14852 4476 15000 4540
rect 10083 4454 15000 4476
rect 10083 4390 10084 4454
rect 10148 4390 10165 4454
rect 10229 4390 10246 4454
rect 10310 4390 10327 4454
rect 10391 4390 10408 4454
rect 10472 4390 10489 4454
rect 10553 4390 10570 4454
rect 10634 4390 10651 4454
rect 10715 4390 10732 4454
rect 10796 4390 10813 4454
rect 10877 4390 10894 4454
rect 10958 4390 10975 4454
rect 11039 4390 11056 4454
rect 11120 4390 11137 4454
rect 11201 4390 11218 4454
rect 11282 4390 11299 4454
rect 11363 4390 11380 4454
rect 11444 4390 11461 4454
rect 11525 4390 11542 4454
rect 11606 4390 11623 4454
rect 11687 4390 11704 4454
rect 11768 4390 11785 4454
rect 11849 4390 11866 4454
rect 11930 4390 11947 4454
rect 12011 4390 12028 4454
rect 12092 4390 12109 4454
rect 12173 4390 12190 4454
rect 12254 4390 12271 4454
rect 12335 4390 12352 4454
rect 12416 4390 12433 4454
rect 12497 4390 12514 4454
rect 12578 4390 12595 4454
rect 12659 4390 12676 4454
rect 12740 4390 12757 4454
rect 12821 4390 12838 4454
rect 12902 4390 12919 4454
rect 12983 4390 13000 4454
rect 13064 4390 13081 4454
rect 13145 4390 13162 4454
rect 13226 4390 13243 4454
rect 13307 4390 13324 4454
rect 13388 4390 13405 4454
rect 13469 4390 13486 4454
rect 13550 4390 13567 4454
rect 13631 4390 13648 4454
rect 13712 4390 13729 4454
rect 13793 4390 13810 4454
rect 13874 4390 13891 4454
rect 13955 4390 13972 4454
rect 14036 4390 14053 4454
rect 14117 4390 14134 4454
rect 14198 4390 14215 4454
rect 14279 4390 14296 4454
rect 14360 4390 14378 4454
rect 14442 4390 14460 4454
rect 14524 4390 14542 4454
rect 14606 4390 14624 4454
rect 14688 4390 14706 4454
rect 14770 4390 14788 4454
rect 14852 4390 15000 4454
rect 10083 4368 15000 4390
rect 10083 4304 10084 4368
rect 10148 4304 10165 4368
rect 10229 4304 10246 4368
rect 10310 4304 10327 4368
rect 10391 4304 10408 4368
rect 10472 4304 10489 4368
rect 10553 4304 10570 4368
rect 10634 4304 10651 4368
rect 10715 4304 10732 4368
rect 10796 4304 10813 4368
rect 10877 4304 10894 4368
rect 10958 4304 10975 4368
rect 11039 4304 11056 4368
rect 11120 4304 11137 4368
rect 11201 4304 11218 4368
rect 11282 4304 11299 4368
rect 11363 4304 11380 4368
rect 11444 4304 11461 4368
rect 11525 4304 11542 4368
rect 11606 4304 11623 4368
rect 11687 4304 11704 4368
rect 11768 4304 11785 4368
rect 11849 4304 11866 4368
rect 11930 4304 11947 4368
rect 12011 4304 12028 4368
rect 12092 4304 12109 4368
rect 12173 4304 12190 4368
rect 12254 4304 12271 4368
rect 12335 4304 12352 4368
rect 12416 4304 12433 4368
rect 12497 4304 12514 4368
rect 12578 4304 12595 4368
rect 12659 4304 12676 4368
rect 12740 4304 12757 4368
rect 12821 4304 12838 4368
rect 12902 4304 12919 4368
rect 12983 4304 13000 4368
rect 13064 4304 13081 4368
rect 13145 4304 13162 4368
rect 13226 4304 13243 4368
rect 13307 4304 13324 4368
rect 13388 4304 13405 4368
rect 13469 4304 13486 4368
rect 13550 4304 13567 4368
rect 13631 4304 13648 4368
rect 13712 4304 13729 4368
rect 13793 4304 13810 4368
rect 13874 4304 13891 4368
rect 13955 4304 13972 4368
rect 14036 4304 14053 4368
rect 14117 4304 14134 4368
rect 14198 4304 14215 4368
rect 14279 4304 14296 4368
rect 14360 4304 14378 4368
rect 14442 4304 14460 4368
rect 14524 4304 14542 4368
rect 14606 4304 14624 4368
rect 14688 4304 14706 4368
rect 14770 4304 14788 4368
rect 14852 4304 15000 4368
rect 10083 4282 15000 4304
rect 10083 4218 10084 4282
rect 10148 4218 10165 4282
rect 10229 4218 10246 4282
rect 10310 4218 10327 4282
rect 10391 4218 10408 4282
rect 10472 4218 10489 4282
rect 10553 4218 10570 4282
rect 10634 4218 10651 4282
rect 10715 4218 10732 4282
rect 10796 4218 10813 4282
rect 10877 4218 10894 4282
rect 10958 4218 10975 4282
rect 11039 4218 11056 4282
rect 11120 4218 11137 4282
rect 11201 4218 11218 4282
rect 11282 4218 11299 4282
rect 11363 4218 11380 4282
rect 11444 4218 11461 4282
rect 11525 4218 11542 4282
rect 11606 4218 11623 4282
rect 11687 4218 11704 4282
rect 11768 4218 11785 4282
rect 11849 4218 11866 4282
rect 11930 4218 11947 4282
rect 12011 4218 12028 4282
rect 12092 4218 12109 4282
rect 12173 4218 12190 4282
rect 12254 4218 12271 4282
rect 12335 4218 12352 4282
rect 12416 4218 12433 4282
rect 12497 4218 12514 4282
rect 12578 4218 12595 4282
rect 12659 4218 12676 4282
rect 12740 4218 12757 4282
rect 12821 4218 12838 4282
rect 12902 4218 12919 4282
rect 12983 4218 13000 4282
rect 13064 4218 13081 4282
rect 13145 4218 13162 4282
rect 13226 4218 13243 4282
rect 13307 4218 13324 4282
rect 13388 4218 13405 4282
rect 13469 4218 13486 4282
rect 13550 4218 13567 4282
rect 13631 4218 13648 4282
rect 13712 4218 13729 4282
rect 13793 4218 13810 4282
rect 13874 4218 13891 4282
rect 13955 4218 13972 4282
rect 14036 4218 14053 4282
rect 14117 4218 14134 4282
rect 14198 4218 14215 4282
rect 14279 4218 14296 4282
rect 14360 4218 14378 4282
rect 14442 4218 14460 4282
rect 14524 4218 14542 4282
rect 14606 4218 14624 4282
rect 14688 4218 14706 4282
rect 14770 4218 14788 4282
rect 14852 4218 15000 4282
rect 10083 4196 15000 4218
rect 10083 4132 10084 4196
rect 10148 4132 10165 4196
rect 10229 4132 10246 4196
rect 10310 4132 10327 4196
rect 10391 4132 10408 4196
rect 10472 4132 10489 4196
rect 10553 4132 10570 4196
rect 10634 4132 10651 4196
rect 10715 4132 10732 4196
rect 10796 4132 10813 4196
rect 10877 4132 10894 4196
rect 10958 4132 10975 4196
rect 11039 4132 11056 4196
rect 11120 4132 11137 4196
rect 11201 4132 11218 4196
rect 11282 4132 11299 4196
rect 11363 4132 11380 4196
rect 11444 4132 11461 4196
rect 11525 4132 11542 4196
rect 11606 4132 11623 4196
rect 11687 4132 11704 4196
rect 11768 4132 11785 4196
rect 11849 4132 11866 4196
rect 11930 4132 11947 4196
rect 12011 4132 12028 4196
rect 12092 4132 12109 4196
rect 12173 4132 12190 4196
rect 12254 4132 12271 4196
rect 12335 4132 12352 4196
rect 12416 4132 12433 4196
rect 12497 4132 12514 4196
rect 12578 4132 12595 4196
rect 12659 4132 12676 4196
rect 12740 4132 12757 4196
rect 12821 4132 12838 4196
rect 12902 4132 12919 4196
rect 12983 4132 13000 4196
rect 13064 4132 13081 4196
rect 13145 4132 13162 4196
rect 13226 4132 13243 4196
rect 13307 4132 13324 4196
rect 13388 4132 13405 4196
rect 13469 4132 13486 4196
rect 13550 4132 13567 4196
rect 13631 4132 13648 4196
rect 13712 4132 13729 4196
rect 13793 4132 13810 4196
rect 13874 4132 13891 4196
rect 13955 4132 13972 4196
rect 14036 4132 14053 4196
rect 14117 4132 14134 4196
rect 14198 4132 14215 4196
rect 14279 4132 14296 4196
rect 14360 4132 14378 4196
rect 14442 4132 14460 4196
rect 14524 4132 14542 4196
rect 14606 4132 14624 4196
rect 14688 4132 14706 4196
rect 14770 4132 14788 4196
rect 14852 4132 15000 4196
rect 10083 4110 15000 4132
rect 10083 4046 10084 4110
rect 10148 4046 10165 4110
rect 10229 4046 10246 4110
rect 10310 4046 10327 4110
rect 10391 4046 10408 4110
rect 10472 4046 10489 4110
rect 10553 4046 10570 4110
rect 10634 4046 10651 4110
rect 10715 4046 10732 4110
rect 10796 4046 10813 4110
rect 10877 4046 10894 4110
rect 10958 4046 10975 4110
rect 11039 4046 11056 4110
rect 11120 4046 11137 4110
rect 11201 4046 11218 4110
rect 11282 4046 11299 4110
rect 11363 4046 11380 4110
rect 11444 4046 11461 4110
rect 11525 4046 11542 4110
rect 11606 4046 11623 4110
rect 11687 4046 11704 4110
rect 11768 4046 11785 4110
rect 11849 4046 11866 4110
rect 11930 4046 11947 4110
rect 12011 4046 12028 4110
rect 12092 4046 12109 4110
rect 12173 4046 12190 4110
rect 12254 4046 12271 4110
rect 12335 4046 12352 4110
rect 12416 4046 12433 4110
rect 12497 4046 12514 4110
rect 12578 4046 12595 4110
rect 12659 4046 12676 4110
rect 12740 4046 12757 4110
rect 12821 4046 12838 4110
rect 12902 4046 12919 4110
rect 12983 4046 13000 4110
rect 13064 4046 13081 4110
rect 13145 4046 13162 4110
rect 13226 4046 13243 4110
rect 13307 4046 13324 4110
rect 13388 4046 13405 4110
rect 13469 4046 13486 4110
rect 13550 4046 13567 4110
rect 13631 4046 13648 4110
rect 13712 4046 13729 4110
rect 13793 4046 13810 4110
rect 13874 4046 13891 4110
rect 13955 4046 13972 4110
rect 14036 4046 14053 4110
rect 14117 4046 14134 4110
rect 14198 4046 14215 4110
rect 14279 4046 14296 4110
rect 14360 4046 14378 4110
rect 14442 4046 14460 4110
rect 14524 4046 14542 4110
rect 14606 4046 14624 4110
rect 14688 4046 14706 4110
rect 14770 4046 14788 4110
rect 14852 4046 15000 4110
rect 10083 4024 15000 4046
rect 10083 3960 10084 4024
rect 10148 3960 10165 4024
rect 10229 3960 10246 4024
rect 10310 3960 10327 4024
rect 10391 3960 10408 4024
rect 10472 3960 10489 4024
rect 10553 3960 10570 4024
rect 10634 3960 10651 4024
rect 10715 3960 10732 4024
rect 10796 3960 10813 4024
rect 10877 3960 10894 4024
rect 10958 3960 10975 4024
rect 11039 3960 11056 4024
rect 11120 3960 11137 4024
rect 11201 3960 11218 4024
rect 11282 3960 11299 4024
rect 11363 3960 11380 4024
rect 11444 3960 11461 4024
rect 11525 3960 11542 4024
rect 11606 3960 11623 4024
rect 11687 3960 11704 4024
rect 11768 3960 11785 4024
rect 11849 3960 11866 4024
rect 11930 3960 11947 4024
rect 12011 3960 12028 4024
rect 12092 3960 12109 4024
rect 12173 3960 12190 4024
rect 12254 3960 12271 4024
rect 12335 3960 12352 4024
rect 12416 3960 12433 4024
rect 12497 3960 12514 4024
rect 12578 3960 12595 4024
rect 12659 3960 12676 4024
rect 12740 3960 12757 4024
rect 12821 3960 12838 4024
rect 12902 3960 12919 4024
rect 12983 3960 13000 4024
rect 13064 3960 13081 4024
rect 13145 3960 13162 4024
rect 13226 3960 13243 4024
rect 13307 3960 13324 4024
rect 13388 3960 13405 4024
rect 13469 3960 13486 4024
rect 13550 3960 13567 4024
rect 13631 3960 13648 4024
rect 13712 3960 13729 4024
rect 13793 3960 13810 4024
rect 13874 3960 13891 4024
rect 13955 3960 13972 4024
rect 14036 3960 14053 4024
rect 14117 3960 14134 4024
rect 14198 3960 14215 4024
rect 14279 3960 14296 4024
rect 14360 3960 14378 4024
rect 14442 3960 14460 4024
rect 14524 3960 14542 4024
rect 14606 3960 14624 4024
rect 14688 3960 14706 4024
rect 14770 3960 14788 4024
rect 14852 3960 15000 4024
rect 10083 3957 15000 3960
rect 0 2987 193 3677
rect 14807 2987 15000 3677
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 18997
rect 14746 14007 15000 18997
rect 0 12837 254 13687
rect 14746 12837 15000 13687
rect 0 11667 254 12517
rect 14746 11667 15000 12517
rect 0 9547 254 11347
rect 14746 9547 15000 11347
rect 0 8337 254 9227
rect 14746 8337 15000 9227
rect 0 7368 254 8017
rect 14746 7368 15000 8017
rect 0 6397 254 7047
rect 14746 6397 15000 7047
rect 0 5187 254 6077
rect 14746 5187 15000 6077
rect 0 3977 254 4867
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 14746 1797 15000 2687
rect 0 427 254 1477
rect 14746 427 15000 1477
use sky130_fd_io__com_bus_hookup  sky130_fd_io__com_bus_hookup_0
timestamp 1619729480
transform 1 0 0 0 1 549
box 0 -142 15000 39451
<< labels >>
flabel metal5 s 14746 35157 15000 40000 3 FreeSans 520 180 0 0 VSSIO
port 44 nsew signal default
flabel metal5 s 14746 7368 15000 8017 3 FreeSans 520 180 0 0 VSSA
port 28 nsew signal default
flabel metal5 s 0 3007 193 3657 3 FreeSans 520 0 0 0 VDDA
port 12 nsew signal default
flabel metal5 s 14746 14007 15000 18997 3 FreeSans 520 180 0 0 VDDIO
port 16 nsew signal default
flabel metal5 s 14746 3977 15000 4867 3 FreeSans 520 180 0 0 VDDIO
port 17 nsew signal default
flabel metal5 s 0 14007 254 18997 3 FreeSans 520 0 0 0 VDDIO
port 18 nsew signal default
flabel metal5 s 0 3977 254 4867 3 FreeSans 520 0 0 0 VDDIO
port 19 nsew signal default
flabel metal5 s 14746 427 15000 1477 3 FreeSans 520 180 0 0 VCCHIB
port 8 nsew signal default
flabel metal5 s 14746 12837 15000 13687 3 FreeSans 520 180 0 0 VDDIO_Q
port 24 nsew signal default
flabel metal5 s 0 12837 254 13687 3 FreeSans 520 0 0 0 VDDIO_Q
port 25 nsew signal default
flabel metal5 s 14746 9547 15000 11347 3 FreeSans 520 180 0 0 VSSA
port 29 nsew signal default
flabel metal5 s 14746 1797 15000 2687 3 FreeSans 520 180 0 0 VCCD
port 4 nsew signal default
flabel metal5 s 0 1797 254 2687 3 FreeSans 520 0 0 0 VCCD
port 5 nsew signal default
flabel metal5 s 0 427 254 1477 3 FreeSans 520 0 0 0 VCCHIB
port 9 nsew signal default
flabel metal5 s 14746 5187 15000 6077 3 FreeSans 520 180 0 0 VSSIO
port 45 nsew signal default
flabel metal5 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 46 nsew signal default
flabel metal5 s 0 5187 254 6077 3 FreeSans 520 0 0 0 VSSIO
port 47 nsew signal default
flabel metal5 s 14746 11667 15000 12517 3 FreeSans 520 180 0 0 VSSIO_Q
port 52 nsew signal default
flabel metal5 s 0 11667 254 12517 3 FreeSans 520 0 0 0 VSSIO_Q
port 53 nsew signal default
flabel metal5 s 14746 6397 15000 7047 3 FreeSans 520 180 0 0 VSWITCH
port 56 nsew signal default
flabel metal5 s 0 6397 254 7047 3 FreeSans 520 0 0 0 VSWITCH
port 57 nsew signal default
flabel metal5 s 0 9547 254 11347 3 FreeSans 520 0 0 0 VSSA
port 30 nsew signal default
flabel metal5 s 0 7368 254 8017 3 FreeSans 520 0 0 0 VSSA
port 31 nsew signal default
flabel metal5 s 14746 8337 15000 9227 3 FreeSans 520 180 0 0 VSSD
port 40 nsew signal default
flabel metal5 s 0 8337 254 9227 3 FreeSans 520 0 0 0 VSSD
port 41 nsew signal default
flabel metal5 s 14807 3007 15000 3657 3 FreeSans 520 180 0 0 VDDA
port 13 nsew signal default
flabel metal4 s 14746 5167 15000 6097 3 FreeSans 520 180 0 0 VSSIO
port 48 nsew signal default
flabel metal4 s 14746 3957 15000 4887 3 FreeSans 520 180 0 0 VDDIO
port 20 nsew signal default
flabel metal4 s 14746 10625 15000 11221 3 FreeSans 520 180 0 0 AMUXBUS_A
port 0 nsew signal default
flabel metal4 s 14746 14007 15000 19000 3 FreeSans 520 180 0 0 VDDIO
port 21 nsew signal default
flabel metal4 s 14746 1777 15000 2707 3 FreeSans 520 180 0 0 VCCD
port 6 nsew signal default
flabel metal4 s 0 3957 254 4887 3 FreeSans 520 0 0 0 VDDIO
port 22 nsew signal default
flabel metal4 s 0 14007 254 19000 3 FreeSans 520 0 0 0 VDDIO
port 23 nsew signal default
flabel metal4 s 14746 12817 15000 13707 3 FreeSans 520 180 0 0 VDDIO_Q
port 26 nsew signal default
flabel metal4 s 0 12817 254 13707 3 FreeSans 520 0 0 0 VDDIO_Q
port 27 nsew signal default
flabel metal4 s 0 9673 254 10269 3 FreeSans 520 0 0 0 AMUXBUS_B
port 2 nsew signal default
flabel metal4 s 14746 7347 15000 8037 3 FreeSans 520 180 0 0 VSSA
port 32 nsew signal default
flabel metal4 s 14746 9547 15000 9613 3 FreeSans 520 180 0 0 VSSA
port 33 nsew signal default
flabel metal4 s 14746 10329 15000 10565 3 FreeSans 520 180 0 0 VSSA
port 34 nsew signal default
flabel metal4 s 14746 11281 15000 11347 3 FreeSans 520 180 0 0 VSSA
port 35 nsew signal default
flabel metal4 s 0 10625 254 11221 3 FreeSans 520 0 0 0 AMUXBUS_A
port 1 nsew signal default
flabel metal4 s 14746 9673 15000 10269 3 FreeSans 520 180 0 0 AMUXBUS_B
port 3 nsew signal default
flabel metal4 s 0 1777 254 2707 3 FreeSans 520 0 0 0 VCCD
port 7 nsew signal default
flabel metal4 s 14746 407 15000 1497 3 FreeSans 520 180 0 0 VCCHIB
port 10 nsew signal default
flabel metal4 s 0 407 254 1497 3 FreeSans 520 0 0 0 VCCHIB
port 11 nsew signal default
flabel metal4 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 49 nsew signal default
flabel metal4 s 0 5167 254 6097 3 FreeSans 520 0 0 0 VSSIO
port 50 nsew signal default
flabel metal4 s 14746 11647 15000 12537 3 FreeSans 520 180 0 0 VSSIO_Q
port 54 nsew signal default
flabel metal4 s 0 11647 254 12537 3 FreeSans 520 0 0 0 VSSIO_Q
port 55 nsew signal default
flabel metal4 s 14746 6377 15000 7067 3 FreeSans 520 180 0 0 VSWITCH
port 58 nsew signal default
flabel metal4 s 0 6377 254 7067 3 FreeSans 520 0 0 0 VSWITCH
port 59 nsew signal default
flabel metal4 s 0 9547 254 9613 3 FreeSans 520 0 0 0 VSSA
port 36 nsew signal default
flabel metal4 s 0 10329 254 10565 3 FreeSans 520 0 0 0 VSSA
port 37 nsew signal default
flabel metal4 s 0 11281 254 11347 3 FreeSans 520 0 0 0 VSSA
port 38 nsew signal default
flabel metal4 s 0 7347 254 8037 3 FreeSans 520 0 0 0 VSSA
port 39 nsew signal default
flabel metal4 s 14746 8317 15000 9247 3 FreeSans 520 180 0 0 VSSD
port 42 nsew signal default
flabel metal4 s 0 8317 254 9247 3 FreeSans 520 0 0 0 VSSD
port 43 nsew signal default
flabel metal4 s 14746 35157 15000 40000 3 FreeSans 520 180 0 0 VSSIO
port 51 nsew signal default
flabel metal4 s 14807 2987 15000 3677 3 FreeSans 520 180 0 0 VDDA
port 14 nsew signal default
flabel metal4 s 0 2987 193 3677 3 FreeSans 520 0 0 0 VDDA
port 15 nsew signal default
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 15000 40000
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string LEFsymmetry X Y R90
string GDS_END 1262564
string GDS_START 637876
<< end >>
