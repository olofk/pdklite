magic
tech sky130A
magscale 1 2
timestamp 1640697677
<< locali >>
rect 191 1160 199 1194
rect 233 1160 271 1194
rect 305 1160 343 1194
rect 377 1160 415 1194
rect 449 1160 487 1194
rect 521 1160 529 1194
rect 191 20 199 54
rect 233 20 271 54
rect 305 20 343 54
rect 377 20 415 54
rect 449 20 487 54
rect 521 20 529 54
<< viali >>
rect 199 1160 233 1194
rect 271 1160 305 1194
rect 343 1160 377 1194
rect 415 1160 449 1194
rect 487 1160 521 1194
rect 199 20 233 54
rect 271 20 305 54
rect 343 20 377 54
rect 415 20 449 54
rect 487 20 521 54
<< obsli1 >>
rect 48 1020 82 1058
rect 48 948 82 986
rect 48 876 82 914
rect 48 804 82 842
rect 48 732 82 770
rect 48 660 82 698
rect 48 588 82 626
rect 48 516 82 554
rect 48 444 82 482
rect 48 372 82 410
rect 48 300 82 338
rect 48 228 82 266
rect 48 122 82 194
rect 159 98 193 1116
rect 251 98 285 1116
rect 343 98 377 1116
rect 435 98 469 1116
rect 527 98 561 1116
rect 638 1020 672 1058
rect 638 948 672 986
rect 638 876 672 914
rect 638 804 672 842
rect 638 732 672 770
rect 638 660 672 698
rect 638 588 672 626
rect 638 516 672 554
rect 638 444 672 482
rect 638 372 672 410
rect 638 300 672 338
rect 638 228 672 266
rect 638 122 672 194
<< obsli1c >>
rect 48 1058 82 1092
rect 48 986 82 1020
rect 48 914 82 948
rect 48 842 82 876
rect 48 770 82 804
rect 48 698 82 732
rect 48 626 82 660
rect 48 554 82 588
rect 48 482 82 516
rect 48 410 82 444
rect 48 338 82 372
rect 48 266 82 300
rect 48 194 82 228
rect 638 1058 672 1092
rect 638 986 672 1020
rect 638 914 672 948
rect 638 842 672 876
rect 638 770 672 804
rect 638 698 672 732
rect 638 626 672 660
rect 638 554 672 588
rect 638 482 672 516
rect 638 410 672 444
rect 638 338 672 372
rect 638 266 672 300
rect 638 194 672 228
<< metal1 >>
rect 187 1194 533 1214
rect 187 1160 199 1194
rect 233 1160 271 1194
rect 305 1160 343 1194
rect 377 1160 415 1194
rect 449 1160 487 1194
rect 521 1160 533 1194
rect 187 1148 533 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 110 94 194
rect 626 1092 684 1104
rect 626 1058 638 1092
rect 672 1058 684 1092
rect 626 1020 684 1058
rect 626 986 638 1020
rect 672 986 684 1020
rect 626 948 684 986
rect 626 914 638 948
rect 672 914 684 948
rect 626 876 684 914
rect 626 842 638 876
rect 672 842 684 876
rect 626 804 684 842
rect 626 770 638 804
rect 672 770 684 804
rect 626 732 684 770
rect 626 698 638 732
rect 672 698 684 732
rect 626 660 684 698
rect 626 626 638 660
rect 672 626 684 660
rect 626 588 684 626
rect 626 554 638 588
rect 672 554 684 588
rect 626 516 684 554
rect 626 482 638 516
rect 672 482 684 516
rect 626 444 684 482
rect 626 410 638 444
rect 672 410 684 444
rect 626 372 684 410
rect 626 338 638 372
rect 672 338 684 372
rect 626 300 684 338
rect 626 266 638 300
rect 672 266 684 300
rect 626 228 684 266
rect 626 194 638 228
rect 672 194 684 228
rect 626 110 684 194
rect 187 54 533 66
rect 187 20 199 54
rect 233 20 271 54
rect 305 20 343 54
rect 377 20 415 54
rect 449 20 487 54
rect 521 20 533 54
rect 187 0 533 20
<< obsm1 >>
rect 150 110 202 1104
rect 242 110 294 1104
rect 334 110 386 1104
rect 426 110 478 1104
rect 518 110 570 1104
<< metal2 >>
rect 10 632 710 1104
rect 10 110 710 582
<< labels >>
rlabel metal1 s 626 110 684 1104 6 BULK
port 1 nsew
rlabel metal1 s 36 110 94 1104 6 BULK
port 1 nsew
rlabel metal2 s 10 632 710 1104 6 DRAIN
port 2 nsew
rlabel viali s 487 1160 521 1194 6 GATE
port 3 nsew
rlabel viali s 487 20 521 54 6 GATE
port 3 nsew
rlabel viali s 415 1160 449 1194 6 GATE
port 3 nsew
rlabel viali s 415 20 449 54 6 GATE
port 3 nsew
rlabel viali s 343 1160 377 1194 6 GATE
port 3 nsew
rlabel viali s 343 20 377 54 6 GATE
port 3 nsew
rlabel viali s 271 1160 305 1194 6 GATE
port 3 nsew
rlabel viali s 271 20 305 54 6 GATE
port 3 nsew
rlabel viali s 199 1160 233 1194 6 GATE
port 3 nsew
rlabel viali s 199 20 233 54 6 GATE
port 3 nsew
rlabel locali s 191 1160 529 1194 6 GATE
port 3 nsew
rlabel locali s 191 20 529 54 6 GATE
port 3 nsew
rlabel metal1 s 187 1148 533 1214 6 GATE
port 3 nsew
rlabel metal1 s 187 0 533 66 6 GATE
port 3 nsew
rlabel metal2 s 10 110 710 582 6 SOURCE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 720 1214
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 9582762
string GDS_START 9560732
<< end >>
