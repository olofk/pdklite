magic
tech sky130A
magscale 1 2
timestamp 1640697850
use sky130_fd_pr__hvdfl1sd__example_55959141808102  sky130_fd_pr__hvdfl1sd__example_55959141808102_0
timestamp 1640697850
transform -1 0 -14 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 145 300 145 300 0 FreeSans 300 0 0 0 D
flabel comment s -42 267 -42 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 7394822
string GDS_START 7393838
<< end >>
