magic
tech sky130A
magscale 1 2
timestamp 1640697980
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 273 157 457 201
rect 1572 181 2198 203
rect 1386 157 2198 181
rect 1 21 2198 157
rect 29 -17 63 21
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 103 427 169 527
rect 18 195 88 325
rect 103 17 169 93
rect 291 427 357 527
rect 686 451 762 527
rect 354 201 436 325
rect 866 451 932 527
rect 1186 451 1268 527
rect 291 17 357 93
rect 722 187 804 213
rect 722 153 765 187
rect 799 153 804 187
rect 722 147 804 153
rect 1402 389 1468 527
rect 722 17 804 105
rect 948 17 1016 109
rect 1332 201 1398 213
rect 1332 187 1464 201
rect 1332 153 1409 187
rect 1443 153 1464 187
rect 1332 147 1464 153
rect 1604 296 1640 527
rect 1334 17 1466 113
rect 1604 17 1640 181
rect 1674 51 1740 493
rect 1774 296 1824 527
rect 1962 299 1996 527
rect 2030 333 2096 493
rect 2130 367 2183 527
rect 2030 299 2183 333
rect 1774 17 1824 181
rect 2072 169 2183 299
rect 2069 165 2183 169
rect 1946 17 2012 165
rect 2046 144 2183 165
rect 2046 51 2096 144
rect 2130 17 2183 110
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 765 153 799 187
rect 1409 153 1443 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< obsli1 >>
rect 35 393 69 493
rect 35 359 168 393
rect 122 161 168 359
rect 35 127 168 161
rect 35 69 69 127
rect 203 69 248 493
rect 391 393 425 493
rect 472 450 638 484
rect 286 359 425 393
rect 286 165 320 359
rect 470 315 570 391
rect 286 127 425 165
rect 470 141 514 315
rect 604 281 638 450
rect 798 417 832 475
rect 1022 433 1152 483
rect 1118 417 1152 433
rect 1308 417 1356 475
rect 672 367 942 417
rect 672 315 722 367
rect 824 281 874 313
rect 604 247 874 281
rect 604 239 688 247
rect 550 129 620 203
rect 391 61 425 127
rect 654 93 688 239
rect 908 213 942 367
rect 862 145 942 213
rect 980 331 1080 393
rect 1118 383 1356 417
rect 980 179 1014 331
rect 1048 213 1084 295
rect 1118 281 1152 383
rect 1502 353 1536 475
rect 1502 349 1566 353
rect 1186 315 1566 349
rect 1118 247 1494 281
rect 1164 179 1230 203
rect 980 145 1230 179
rect 485 53 688 93
rect 862 59 912 145
rect 1264 95 1298 247
rect 1428 235 1494 247
rect 1528 136 1566 315
rect 1128 61 1298 95
rect 1502 70 1566 136
rect 1862 265 1928 493
rect 1862 199 2038 265
rect 1862 51 1912 199
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 753 187 811 193
rect 753 153 765 187
rect 799 184 811 187
rect 1397 187 1455 193
rect 1397 184 1409 187
rect 799 156 1409 184
rect 799 153 811 156
rect 753 147 811 153
rect 1397 153 1409 156
rect 1443 153 1455 187
rect 1397 147 1455 153
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< obsm1 >>
rect 117 388 175 397
rect 477 388 535 397
rect 1029 388 1087 397
rect 117 360 1087 388
rect 117 351 175 360
rect 477 351 535 360
rect 1029 351 1087 360
rect 1037 252 1095 261
rect 584 224 1095 252
rect 584 193 627 224
rect 1037 215 1095 224
rect 201 184 259 193
rect 569 184 627 193
rect 201 156 627 184
rect 201 147 259 156
rect 569 147 627 156
<< labels >>
rlabel locali s 18 195 88 325 6 CLK
port 1 nsew clock input
rlabel locali s 354 201 436 325 6 D
port 2 nsew signal input
rlabel metal1 s 1397 147 1455 156 6 SET_B
port 3 nsew signal input
rlabel metal1 s 753 147 811 156 6 SET_B
port 3 nsew signal input
rlabel metal1 s 753 156 1455 184 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1397 184 1455 193 6 SET_B
port 3 nsew signal input
rlabel metal1 s 753 184 811 193 6 SET_B
port 3 nsew signal input
rlabel viali s 1409 153 1443 187 6 SET_B
port 3 nsew signal input
rlabel locali s 1332 147 1464 201 6 SET_B
port 3 nsew signal input
rlabel locali s 1332 201 1398 213 6 SET_B
port 3 nsew signal input
rlabel viali s 765 153 799 187 6 SET_B
port 3 nsew signal input
rlabel locali s 722 147 804 213 6 SET_B
port 3 nsew signal input
rlabel metal1 s 0 -48 2208 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 2145 -17 2179 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 2053 -17 2087 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1961 -17 1995 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1869 -17 1903 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1777 -17 1811 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1685 -17 1719 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1593 -17 1627 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1501 -17 1535 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1409 -17 1443 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1317 -17 1351 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1225 -17 1259 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1133 -17 1167 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 1041 -17 1075 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 949 -17 983 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 857 -17 891 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 765 -17 799 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 673 -17 707 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 581 -17 615 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 489 -17 523 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 397 -17 431 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 305 -17 339 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 213 -17 247 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 121 -17 155 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 29 -17 63 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 2208 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 2130 17 2183 110 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1946 17 2012 165 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1774 17 1824 181 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1604 17 1640 181 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 1334 17 1466 113 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 948 17 1016 109 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 722 17 804 105 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 291 17 357 93 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 103 17 169 93 6 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 2198 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1386 157 2198 181 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1572 181 2198 203 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 273 157 457 201 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 2246 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 2208 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 2145 527 2179 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 2053 527 2087 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1961 527 1995 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1869 527 1903 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1777 527 1811 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1685 527 1719 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1593 527 1627 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1501 527 1535 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1409 527 1443 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1317 527 1351 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1225 527 1259 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1133 527 1167 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 1041 527 1075 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 949 527 983 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 857 527 891 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 765 527 799 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 673 527 707 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 581 527 615 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 489 527 523 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 397 527 431 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 305 527 339 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 213 527 247 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 121 527 155 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 29 527 63 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 2130 367 2183 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1962 299 1996 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1774 296 1824 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1604 296 1640 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1402 389 1468 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1186 451 1268 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 866 451 932 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 686 451 762 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 291 427 357 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 427 169 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 2208 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 2046 51 2096 144 6 Q
port 8 nsew signal output
rlabel locali s 2046 144 2183 165 6 Q
port 8 nsew signal output
rlabel locali s 2069 165 2183 169 6 Q
port 8 nsew signal output
rlabel locali s 2072 169 2183 299 6 Q
port 8 nsew signal output
rlabel locali s 2030 299 2183 333 6 Q
port 8 nsew signal output
rlabel locali s 2030 333 2096 493 6 Q
port 8 nsew signal output
rlabel locali s 1674 51 1740 493 6 Q_N
port 9 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2208 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2515242
string GDS_START 2496374
<< end >>
