magic
tech sky130A
magscale 1 2
timestamp 1619729485
<< obsli1 >>
rect 214 200 14555 39939
<< obsm1 >>
rect 37 194 14724 39945
<< metal2 >>
rect 5179 0 5579 107
<< obsm2 >>
rect 53 163 14858 39015
rect 53 0 5123 163
rect 5635 0 14858 163
<< metal3 >>
rect 2810 34321 5002 39020
rect 5186 35070 7364 39020
rect 2810 34261 3100 34321
rect 4300 34261 5002 34321
rect 3100 33826 5002 34261
rect 3100 20936 4300 33826
rect 7246 35052 7364 35070
rect 5186 34962 7364 35052
rect 7246 34952 7364 34962
rect 7108 34932 7246 34952
rect 5186 34842 7246 34932
rect 7108 34814 7246 34842
rect 6958 34812 7108 34814
rect 5186 34692 7108 34812
rect 6958 34664 7108 34692
rect 6845 34662 6958 34664
rect 5186 34572 6958 34662
rect 6845 34551 6958 34572
rect 6386 34542 6845 34551
rect 5186 34092 6845 34542
rect 5186 20972 6386 34092
rect 7593 34152 9771 38004
rect 7593 34122 8571 34152
rect 7593 34092 9771 34122
rect 8571 22124 9771 34092
rect 5186 20936 7379 20972
rect 3100 20099 7379 20936
rect 3100 20051 5614 20099
rect 6386 20069 7379 20099
rect 3100 20021 3661 20051
rect 4300 20050 5614 20051
rect 5625 20050 7379 20069
rect 5186 20021 5607 20050
rect 3100 19931 5607 20021
rect 3100 19879 3661 19931
rect 5186 19901 5607 19931
rect 3669 19879 5607 19901
rect 3661 19631 5607 19879
rect 3661 19601 4207 19631
rect 5186 19629 5607 19631
rect 5614 20009 7379 20050
rect 5614 19979 6035 20009
rect 6386 19979 7379 20009
rect 5614 19665 7379 19979
rect 5614 19629 6035 19665
rect 6389 19635 7379 19665
rect 6059 19629 7379 19635
rect 5607 19601 5905 19629
rect 3661 19391 5905 19601
rect 3661 19333 4207 19391
rect 4207 19331 4749 19333
rect 5607 19331 5905 19391
rect 4207 18791 5905 19331
rect 6035 19275 7379 19629
rect 4749 18620 5905 18791
rect 4749 18493 6047 18620
rect 6389 18620 7379 19275
rect 4749 18478 5027 18493
rect 5905 18478 6047 18493
rect 6247 18478 7379 18620
rect 4749 18288 7379 18478
rect 4749 18230 5027 18288
rect 6389 18258 7379 18288
rect 5029 18230 7379 18258
rect 5027 18138 7379 18230
rect 5027 18108 5179 18138
rect 6389 18108 7379 18138
rect 5027 18078 7379 18108
rect 5179 0 7379 18078
rect 7578 21630 9771 22124
rect 9955 34936 12189 38008
rect 11857 34934 12189 34936
rect 9955 34604 12189 34934
rect 9955 33887 11857 34604
rect 9955 33857 10657 33887
rect 9955 33827 11857 33857
rect 10657 22088 11857 33827
rect 10199 21630 11857 22088
rect 7578 21611 8571 21630
rect 9343 21611 10199 21630
rect 10221 21622 11857 21630
rect 7578 21563 10199 21611
rect 10657 21592 11857 21622
rect 10208 21563 11857 21592
rect 7578 21221 11857 21563
rect 7578 21191 8571 21221
rect 9343 21202 11857 21221
rect 9048 21191 9343 21202
rect 7578 20907 9343 21191
rect 9476 21143 9771 21202
rect 9772 21173 11857 21202
rect 10208 21143 11857 21173
rect 9476 20907 11857 21143
rect 8568 20877 9048 20907
rect 7578 20427 9048 20877
rect 9052 20873 9476 20907
rect 9502 20903 11857 20907
rect 10208 20873 11857 20903
rect 7578 20043 8568 20427
rect 7578 20021 8710 20043
rect 8568 19991 8710 20021
rect 7578 19901 8710 19991
rect 9052 20043 11857 20873
rect 12300 20259 14858 34664
rect 8910 20033 11857 20043
rect 8910 20003 9052 20033
rect 10208 20003 11857 20033
rect 8910 19943 11857 20003
rect 11984 20257 14858 20259
rect 11984 20227 12300 20257
rect 11984 19943 14858 20227
rect 8910 19901 10208 19943
rect 7578 19660 10208 19901
rect 11271 19897 11984 19943
rect 11998 19927 14858 19943
rect 9778 19650 10208 19660
rect 7578 19230 10208 19650
rect 11271 19230 14858 19897
rect 7578 0 9778 19230
rect 10078 19177 11271 19230
rect 11278 19207 14858 19230
rect 10078 0 14858 19177
<< obsm3 >>
rect 48 34181 2730 35070
rect 48 19799 3020 34181
rect 5082 33746 5106 35070
rect 7444 34872 7513 35070
rect 7326 34734 7513 34872
rect 7188 34584 7513 34734
rect 4380 21016 5106 33746
rect 7038 34471 7513 34584
rect 6925 34012 7513 34471
rect 6466 22204 8491 34012
rect 6466 21052 7498 22204
rect 48 19253 3581 19799
rect 48 18711 4127 19253
rect 48 18150 4669 18711
rect 5985 18700 6309 19195
rect 6127 18558 6167 18700
rect 48 17998 4947 18150
rect 48 0 5099 17998
rect 7459 0 7498 21052
rect 9851 33747 9875 35070
rect 12269 34744 14858 35070
rect 9851 22168 10577 33747
rect 9851 21710 10119 22168
rect 8648 20123 8972 20347
rect 8790 19981 8830 20123
rect 11937 20339 12220 34524
rect 10288 19310 11191 19863
rect 9858 0 9998 19150
<< metal4 >>
rect 0 10625 15000 11221
rect 0 9673 15000 10269
<< obsm4 >>
rect 0 11301 15000 40000
rect 0 10349 15000 10545
rect 0 407 15000 9593
<< metal5 >>
rect 1220 20802 13760 33325
rect 14746 14007 15000 18997
rect 14746 12837 15000 13687
rect 14746 11667 15000 12517
rect 14746 9547 15000 11347
rect 14746 8337 15000 9227
rect 14746 6397 15000 7047
rect 14746 5187 15000 6077
rect 14807 3007 15000 3657
rect 14746 1797 15000 2687
rect 14746 427 15000 1477
<< obsm5 >>
rect 0 33645 15000 40000
rect 0 20482 900 33645
rect 14080 20482 15000 33645
rect 0 19317 15000 20482
rect 0 8017 14426 19317
rect 0 7367 15000 8017
rect 0 4867 14426 7367
rect 0 3977 15000 4867
rect 0 3007 14487 3977
rect 0 427 14426 3007
<< labels >>
rlabel metal4 s 0 10625 15000 11221 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 9673 15000 10269 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal5 s 1220 20802 13760 33325 6 G_PAD
port 3 nsew signal bidirectional
rlabel metal3 s 7578 0 9778 19230 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20021 8568 20043 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20043 8568 20427 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20427 8568 20457 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20457 8598 20487 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20487 8628 20517 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20517 8658 20547 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20547 8688 20577 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20577 8718 20607 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20607 8748 20637 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20637 8778 20667 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20667 8808 20697 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20697 8838 20727 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20727 8868 20757 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20757 8898 20787 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20787 8928 20817 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20817 8958 20847 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20847 8988 20877 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20907 9048 20937 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20937 9078 20967 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20967 9108 20997 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 20997 9138 21027 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 21027 9168 21057 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 21057 9198 21087 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 21087 9228 21117 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 21117 9258 21131 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 21131 8571 22124 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19230 9778 19260 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19260 9808 19290 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19290 9838 19320 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19320 9868 19350 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19350 9898 19380 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19380 9928 19410 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19410 9958 19440 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19440 9988 19470 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19470 10018 19500 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19500 10048 19530 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19530 10078 19560 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19560 10108 19590 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19590 10138 19620 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19620 10168 19650 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19660 10208 19901 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19901 8680 19931 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19931 8650 19961 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7578 19961 8620 19991 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7593 34092 8571 35070 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7593 35070 9771 38004 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7608 21131 9272 21161 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7611 35052 9771 35070 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7638 21161 9302 21191 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7641 35022 9771 35052 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7671 34992 9771 35022 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7698 21221 9362 21251 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7701 34962 9771 34992 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7728 21251 9392 21281 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7731 34932 9771 34962 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7758 21281 9422 21311 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7761 34902 9771 34932 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7788 21311 9452 21341 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7791 34872 9771 34902 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7818 21341 9482 21371 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7821 34842 9771 34872 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7848 21371 9512 21401 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7851 34812 9771 34842 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7878 21401 9542 21431 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7881 34782 9771 34812 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7908 21431 9572 21461 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7911 34752 9771 34782 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7938 21461 9602 21491 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7941 34722 9771 34752 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7968 21491 9632 21521 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7971 34692 9771 34722 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 7998 21521 9662 21551 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8001 34662 9771 34692 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8028 21551 9692 21581 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8031 34632 9771 34662 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8058 21581 9722 21611 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8061 34602 9771 34632 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8091 34572 9771 34602 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8107 21630 9771 21660 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8121 34542 9771 34572 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8137 21660 9771 21690 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8151 34512 9771 34542 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8167 21690 9771 21720 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8181 34482 9771 34512 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8197 21720 9771 21750 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8211 34452 9771 34482 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8227 21750 9771 21780 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8241 34422 9771 34452 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8257 21780 9771 21810 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8271 34392 9771 34422 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8287 21810 9771 21840 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8301 34362 9771 34392 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8317 21840 9771 21870 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8331 34332 9771 34362 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8347 21870 9771 21900 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8361 34302 9771 34332 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8377 21900 9771 21930 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8391 34272 9771 34302 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8407 21930 9771 21960 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8421 34242 9771 34272 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8437 21960 9771 21990 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8451 34212 9771 34242 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8467 21990 9771 22020 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8481 34182 9771 34212 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8497 22020 9771 22050 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8511 34152 9771 34182 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8527 22050 9771 22080 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8568 20427 9048 20907 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8568 19901 8710 20043 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8571 21630 9771 22124 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8571 22124 9771 34092 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8571 34092 9771 34122 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8910 19901 9052 20043 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8931 19901 10208 19922 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8952 19922 10208 19943 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 8982 19943 10208 19973 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9012 19973 10238 20003 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9048 20907 9343 21202 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20033 10298 20043 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20043 10308 20073 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20073 10338 20103 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20103 10368 20133 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20133 10398 20163 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20163 10428 20193 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20193 10458 20223 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20223 10488 20253 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20253 10518 20283 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20283 10548 20313 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20313 10578 20343 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20343 10608 20373 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20373 10638 20403 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20403 10668 20433 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20433 10698 20463 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20463 10728 20483 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9052 20483 9476 20907 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9082 20483 10748 20513 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9112 20513 10778 20543 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9142 20543 10808 20573 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9172 20573 10838 20603 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9202 20603 10868 20633 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9232 20633 10898 20663 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9262 20663 10928 20693 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9292 20693 10958 20723 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9322 20723 10988 20753 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9343 21202 9771 21630 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9352 20753 11018 20783 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9382 20783 11048 20813 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9412 20813 11078 20843 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9442 20843 11108 20873 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9476 20907 9771 21202 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9502 20903 11168 20933 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9532 20933 11198 20963 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9562 20963 11228 20993 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9592 20993 11258 21023 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9622 21023 11288 21053 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9652 21053 11318 21083 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9682 21083 11348 21113 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9712 21113 11378 21143 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9771 21202 10199 21630 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9772 21173 11438 21203 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9778 19230 10208 19660 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9802 21203 11468 21233 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9832 21233 11498 21263 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9862 21263 11528 21293 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9892 21293 11558 21323 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9922 21323 11588 21353 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9952 21353 11618 21383 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 33827 10657 34529 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34529 11857 34604 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34529 11857 34634 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34634 11887 34664 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34664 11917 34694 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34694 11947 34724 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34724 11977 34754 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34754 12007 34784 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34784 12037 34814 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34814 12067 34844 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34844 12097 34874 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34874 12127 34904 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34904 12157 34934 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9955 34936 12189 38008 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9967 34517 11857 34529 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9982 21383 11648 21413 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 9997 34487 11857 34517 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10012 21413 11678 21443 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10027 34457 11857 34487 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10042 21443 11708 21473 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10057 34427 11857 34457 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10072 21473 11738 21503 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10087 34397 11857 34427 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10102 21503 11768 21533 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10117 34367 11857 34397 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10132 21533 11798 21563 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10147 34337 11857 34367 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10177 34307 11857 34337 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10199 21630 10657 22088 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10207 34277 11857 34307 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10208 19943 11857 21592 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10221 21622 11857 21652 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10237 34247 11857 34277 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10251 21652 11857 21682 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10267 34217 11857 34247 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10281 21682 11857 21712 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10297 34187 11857 34217 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10311 21712 11857 21742 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10327 34157 11857 34187 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10341 21742 11857 21772 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10357 34127 11857 34157 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10371 21772 11857 21802 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10387 34097 11857 34127 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10401 21802 11857 21832 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10417 34067 11857 34097 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10431 21832 11857 21862 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10447 34037 11857 34067 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10461 21862 11857 21892 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10477 34007 11857 34037 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10491 21892 11857 21922 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10507 33977 11857 34007 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10521 21922 11857 21952 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10537 33947 11857 33977 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10551 21952 11857 21982 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10567 33917 11857 33947 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10581 21982 11857 22012 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10597 33887 11857 33917 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10611 22012 11857 22042 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10657 21592 11857 22088 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10657 22088 11857 33827 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10657 33827 11857 33857 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 11857 34604 12189 34936 6 DRN_HVC
port 4 nsew power bidirectional
rlabel metal3 s 10078 0 14858 18037 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10078 18037 11271 19230 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10108 18037 14858 18067 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10138 18067 14858 18097 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10168 18097 14858 18127 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10198 18127 14858 18157 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10228 18157 14858 18187 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10258 18187 14858 18217 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10288 18217 14858 18247 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10318 18247 14858 18277 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10348 18277 14858 18307 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10378 18307 14858 18337 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10408 18337 14858 18367 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10438 18367 14858 18397 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10468 18397 14858 18427 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10498 18427 14858 18457 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10528 18457 14858 18487 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10558 18487 14858 18517 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10588 18517 14858 18547 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10618 18547 14858 18577 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10648 18577 14858 18607 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10678 18607 14858 18637 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10708 18637 14858 18667 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10738 18667 14858 18697 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10768 18697 14858 18727 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10798 18727 14858 18757 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10828 18757 14858 18787 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10858 18787 14858 18817 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10888 18817 14858 18847 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10918 18847 14858 18877 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10948 18877 14858 18907 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 10978 18907 14858 18937 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11008 18937 14858 18967 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11038 18967 14858 18997 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11068 18997 14858 19027 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11098 19027 14858 19057 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11128 19057 14858 19087 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11158 19087 14858 19117 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11188 19117 14858 19147 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11218 19147 14858 19177 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11271 19230 11984 19943 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11278 19207 14858 19237 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11308 19237 14858 19267 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11338 19267 14858 19297 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11368 19297 14858 19327 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11398 19327 14858 19357 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11428 19357 14858 19387 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11458 19387 14858 19417 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11488 19417 14858 19447 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11518 19447 14858 19477 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11548 19477 14858 19507 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11578 19507 14858 19537 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11608 19537 14858 19567 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11638 19567 14858 19597 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11668 19597 14858 19627 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11698 19627 14858 19657 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11728 19657 14858 19687 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11758 19687 14858 19717 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11788 19717 14858 19747 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11818 19747 14858 19777 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11848 19777 14858 19807 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11878 19807 14858 19837 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11908 19837 14858 19867 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11938 19867 14858 19897 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11984 19943 12300 20259 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 11998 19927 14858 19957 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 12028 19957 14858 19987 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 12058 19987 14858 20017 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 12088 20017 14858 20047 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 12118 20047 14858 20077 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 12148 20077 14858 20107 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 12178 20107 14858 20137 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 12208 20137 14858 20167 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 12238 20167 14858 20197 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 12268 20197 14858 20227 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 12300 20257 14858 20259 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal3 s 12300 20259 14858 34664 6 G_CORE
port 5 nsew ground bidirectional
rlabel metal2 s 5179 0 5579 107 6 OGC_HVC
port 6 nsew power bidirectional
rlabel metal3 s 2810 34261 3100 34551 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2810 34551 5002 39020 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2811 34550 5002 34551 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2822 34539 5002 34550 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2833 34528 5002 34539 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2860 34501 4975 34528 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2890 34471 4945 34501 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2920 34441 4915 34471 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2950 34411 4885 34441 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 2980 34381 4855 34411 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3010 34351 4825 34381 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3040 34321 4795 34351 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20440 4766 20470 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20470 4736 20500 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20500 4706 20530 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20530 4676 20560 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20560 4646 20590 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20590 4616 20620 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20620 4586 20650 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20650 4556 20680 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20680 4526 20710 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20710 4496 20740 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20740 4466 20770 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20770 4436 20800 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20800 4406 20830 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20830 4376 20860 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20860 4346 20890 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20890 4316 20920 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20920 4300 20936 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 20936 4300 33826 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 31694 4300 33856 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 33856 4330 33886 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 33886 4360 33916 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 33916 4390 33946 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 33946 4420 33976 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 33976 4450 34006 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34006 4480 34036 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34036 4510 34066 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34066 4540 34096 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34096 4570 34126 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34126 4600 34156 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34156 4630 34186 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34186 4660 34216 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34216 4690 34246 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 34246 4720 34261 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3100 19879 3661 20440 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3129 20411 4796 20440 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3159 20381 4825 20411 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3189 20351 4855 20381 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3219 20321 4885 20351 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3249 20291 4915 20321 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3279 20261 4945 20291 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3309 20231 4975 20261 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3339 20201 5005 20231 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3369 20171 5035 20201 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3399 20141 5065 20171 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3429 20111 5095 20141 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3459 20081 5125 20111 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3489 20051 5155 20081 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3549 19991 5215 20021 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3579 19961 5245 19991 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3609 19931 5275 19961 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3661 19333 4207 19879 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3669 19871 5335 19901 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3699 19841 5365 19871 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3729 19811 5395 19841 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3759 19781 5425 19811 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3789 19751 5455 19781 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3819 19721 5485 19751 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3849 19691 5515 19721 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3879 19661 5545 19691 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3909 19631 5575 19661 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3969 19571 5635 19601 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 3999 19541 5665 19571 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4029 19511 5695 19541 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4059 19481 5725 19511 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4089 19451 5755 19481 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4119 19421 5785 19451 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4149 19391 5815 19421 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4207 18791 4749 19333 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4239 19301 5905 19331 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4269 19271 5905 19301 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4299 19241 5905 19271 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4300 20050 5186 20936 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4300 33826 5002 34528 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4329 19211 5905 19241 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4359 19181 5905 19211 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4389 19151 5905 19181 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4419 19121 5905 19151 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4449 19091 5905 19121 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4479 19061 5905 19091 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4509 19031 5905 19061 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4539 19001 5905 19031 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4569 18971 5905 19001 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4599 18941 5905 18971 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4629 18911 5905 18941 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4659 18881 5905 18911 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4689 18851 5905 18881 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4749 18230 5027 18508 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4749 18508 5905 19331 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4749 18508 5987 18538 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4749 18538 5957 18568 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4749 18568 5927 18598 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4749 18598 5905 18620 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4749 18620 5905 18791 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4764 18493 6017 18508 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4789 18468 7379 18478 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4819 18438 7379 18468 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4849 18408 7379 18438 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4879 18378 7379 18408 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4909 18348 7379 18378 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4939 18318 7379 18348 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 4969 18288 7379 18318 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5027 18078 5179 18230 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5029 18228 7379 18258 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5059 18198 7379 18228 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5089 18168 7379 18198 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5119 18138 7379 18168 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5179 0 7379 18078 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5179 18078 7379 18108 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20050 5614 20478 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20478 6850 20508 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20508 6820 20538 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20538 6790 20568 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20568 6760 20598 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20598 6730 20628 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20628 6700 20658 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20658 6670 20688 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20688 6640 20718 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20718 6610 20748 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20748 6580 20778 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20778 6550 20808 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20808 6520 20838 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20838 6490 20868 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20868 6460 20898 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20898 6430 20928 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20928 6400 20958 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20958 6386 20972 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 20972 6386 34092 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 31694 6386 34122 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34122 6416 34152 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34152 6446 34182 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34182 6476 34212 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34212 6506 34242 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34242 6536 34272 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34272 6566 34302 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34302 6596 34332 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34332 6626 34362 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34362 6656 34392 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34392 6686 34422 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34422 6716 34452 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34452 6746 34482 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34482 6776 34512 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34512 6806 34542 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34572 6866 34602 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34602 6896 34632 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34632 6926 34662 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34692 6986 34722 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34722 7016 34752 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34752 7046 34782 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34782 7076 34812 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34842 7136 34872 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34872 7166 34902 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34902 7196 34932 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34962 7256 34992 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 34992 7286 35022 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 35022 7316 35052 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 35070 7364 39020 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5186 19629 5607 20050 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5205 20459 6880 20478 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5235 20429 6899 20459 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5265 20399 6929 20429 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5295 20369 6959 20399 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5325 20339 6989 20369 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5355 20309 7019 20339 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5385 20279 7049 20309 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5415 20249 7079 20279 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5445 20219 7109 20249 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5475 20189 7139 20219 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5505 20159 7169 20189 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5535 20129 7199 20159 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5565 20099 7229 20129 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5607 19331 5905 19629 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5614 19629 6035 20050 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5625 20039 7289 20069 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5655 20009 7319 20039 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5699 19965 7379 19979 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5729 19935 7379 19965 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5759 19905 7379 19935 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5789 19875 7379 19905 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5819 19845 7379 19875 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5849 19815 7379 19845 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5879 19785 7379 19815 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5905 18478 6047 18620 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5909 19755 7379 19785 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5939 19725 7379 19755 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5969 19695 7379 19725 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 5999 19665 7379 19695 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6035 19275 6389 19629 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6059 19605 7379 19635 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6089 19575 7379 19605 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6119 19545 7379 19575 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6149 19515 7379 19545 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6179 19485 7379 19515 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6209 19455 7379 19485 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6239 19425 7379 19455 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6247 18478 6389 18620 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6269 19395 7379 19425 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6277 18478 7379 18508 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6299 19365 7379 19395 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6307 18508 7379 18538 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6329 19335 7379 19365 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6337 18538 7379 18568 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6386 34092 6845 34551 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6386 19979 7379 20972 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6389 17894 7379 19979 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6389 18598 7379 18620 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6389 18620 7379 19275 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6845 34551 6958 34664 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 6958 34664 7108 34814 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 7108 34814 7246 34952 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal3 s 7246 34952 7364 35070 6 SRC_BDY_HVC
port 7 nsew ground bidirectional
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 8 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 9 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 10 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 11 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 12 nsew power bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 13 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 14 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 15 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 16 nsew ground bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 17 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 15000 40000
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 31544388
string GDS_START 27543042
<< end >>
