magic
tech sky130A
magscale 1 2
timestamp 1640697996
<< nwell >>
rect -66 377 738 897
<< pwell >>
rect 60 43 653 283
rect -26 -43 698 43
<< locali >>
rect 240 415 274 751
rect 596 415 647 751
rect 240 381 647 415
rect 25 301 199 367
rect 377 162 455 345
rect 491 162 545 345
rect 596 265 647 381
rect 581 99 647 265
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 18 735 204 751
rect 18 701 22 735
rect 56 701 94 735
rect 128 701 166 735
rect 200 701 204 735
rect 18 435 204 701
rect 310 735 560 751
rect 344 701 382 735
rect 416 701 454 735
rect 488 701 526 735
rect 310 451 560 701
rect 18 113 341 265
rect 18 79 19 113
rect 53 79 91 113
rect 125 79 163 113
rect 197 79 235 113
rect 269 79 307 113
rect 18 73 341 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 22 701 56 735
rect 94 701 128 735
rect 166 701 200 735
rect 310 701 344 735
rect 382 701 416 735
rect 454 701 488 735
rect 526 701 560 735
rect 19 79 53 113
rect 91 79 125 113
rect 163 79 197 113
rect 235 79 269 113
rect 307 79 341 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 831 672 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 0 791 672 797
rect 0 735 672 763
rect 0 701 22 735
rect 56 701 94 735
rect 128 701 166 735
rect 200 701 310 735
rect 344 701 382 735
rect 416 701 454 735
rect 488 701 526 735
rect 560 701 672 735
rect 0 689 672 701
rect 0 113 672 125
rect 0 79 19 113
rect 53 79 91 113
rect 125 79 163 113
rect 197 79 235 113
rect 269 79 307 113
rect 341 79 672 113
rect 0 51 672 79
rect 0 17 672 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -23 672 -17
<< labels >>
rlabel locali s 491 162 545 345 6 A
port 1 nsew signal input
rlabel locali s 377 162 455 345 6 B
port 2 nsew signal input
rlabel locali s 25 301 199 367 6 C
port 3 nsew signal input
rlabel metal1 s 0 51 672 125 6 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 -23 672 23 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s -26 -43 698 43 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s 60 43 653 283 6 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 791 672 837 6 VPB
port 6 nsew power bidirectional
rlabel nwell s -66 377 738 897 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 689 672 763 6 VPWR
port 7 nsew power bidirectional
rlabel locali s 581 99 647 265 6 Y
port 8 nsew signal output
rlabel locali s 596 265 647 381 6 Y
port 8 nsew signal output
rlabel locali s 240 381 647 415 6 Y
port 8 nsew signal output
rlabel locali s 596 415 647 751 6 Y
port 8 nsew signal output
rlabel locali s 240 415 274 751 6 Y
port 8 nsew signal output
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 672 814
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_END 204742
string GDS_START 195378
<< end >>
