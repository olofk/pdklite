magic
tech sky130A
magscale 1 2
timestamp 1619729573
<< checkpaint >>
rect -1326 -1283 1806 2157
<< nwell >>
rect -66 377 546 897
<< pwell >>
rect 0 -17 480 17
<< mvnmos >>
rect 133 111 233 261
rect 275 111 375 261
<< mvpmos >>
rect 133 443 233 743
rect 289 443 389 743
<< mvndiff >>
rect 76 253 133 261
rect 76 219 88 253
rect 122 219 133 253
rect 76 153 133 219
rect 76 119 88 153
rect 122 119 133 153
rect 76 111 133 119
rect 233 111 275 261
rect 375 253 432 261
rect 375 219 386 253
rect 420 219 432 253
rect 375 153 432 219
rect 375 119 386 153
rect 420 119 432 153
rect 375 111 432 119
<< mvpdiff >>
rect 76 735 133 743
rect 76 701 88 735
rect 122 701 133 735
rect 76 652 133 701
rect 76 618 88 652
rect 122 618 133 652
rect 76 568 133 618
rect 76 534 88 568
rect 122 534 133 568
rect 76 485 133 534
rect 76 451 88 485
rect 122 451 133 485
rect 76 443 133 451
rect 233 735 289 743
rect 233 701 244 735
rect 278 701 289 735
rect 233 652 289 701
rect 233 618 244 652
rect 278 618 289 652
rect 233 568 289 618
rect 233 534 244 568
rect 278 534 289 568
rect 233 485 289 534
rect 233 451 244 485
rect 278 451 289 485
rect 233 443 289 451
rect 389 735 446 743
rect 389 701 400 735
rect 434 701 446 735
rect 389 652 446 701
rect 389 618 400 652
rect 434 618 446 652
rect 389 568 446 618
rect 389 534 400 568
rect 434 534 446 568
rect 389 485 446 534
rect 389 451 400 485
rect 434 451 446 485
rect 389 443 446 451
<< mvndiffc >>
rect 88 219 122 253
rect 88 119 122 153
rect 386 219 420 253
rect 386 119 420 153
<< mvpdiffc >>
rect 88 701 122 735
rect 88 618 122 652
rect 88 534 122 568
rect 88 451 122 485
rect 244 701 278 735
rect 244 618 278 652
rect 244 534 278 568
rect 244 451 278 485
rect 400 701 434 735
rect 400 618 434 652
rect 400 534 434 568
rect 400 451 434 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 480 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
<< poly >>
rect 133 743 233 769
rect 289 743 389 769
rect 133 371 233 443
rect 289 417 389 443
rect 133 337 153 371
rect 187 337 233 371
rect 133 261 233 337
rect 275 355 459 417
rect 275 321 405 355
rect 439 321 459 355
rect 275 287 459 321
rect 275 261 375 287
rect 133 85 233 111
rect 275 85 375 111
<< polycont >>
rect 153 337 187 371
rect 405 321 439 355
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 480 831
rect 18 735 208 751
rect 18 701 24 735
rect 58 701 88 735
rect 130 701 168 735
rect 202 701 208 735
rect 18 652 208 701
rect 18 618 88 652
rect 122 618 208 652
rect 18 568 208 618
rect 18 534 88 568
rect 122 534 208 568
rect 18 485 208 534
rect 18 451 88 485
rect 122 451 208 485
rect 18 435 208 451
rect 244 735 294 751
rect 278 701 294 735
rect 244 652 294 701
rect 278 618 294 652
rect 244 568 294 618
rect 278 534 294 568
rect 244 485 294 534
rect 278 451 294 485
rect 25 371 203 387
rect 25 337 153 371
rect 187 337 203 371
rect 25 310 203 337
rect 244 339 294 451
rect 332 735 450 751
rect 332 701 338 735
rect 372 701 400 735
rect 444 701 450 735
rect 332 652 450 701
rect 332 618 400 652
rect 434 618 450 652
rect 332 568 450 618
rect 332 534 400 568
rect 434 534 450 568
rect 332 485 450 534
rect 332 451 400 485
rect 434 451 450 485
rect 332 435 450 451
rect 395 355 455 371
rect 244 305 359 339
rect 395 321 405 355
rect 439 321 455 355
rect 395 305 455 321
rect 316 269 359 305
rect 18 253 280 269
rect 18 219 88 253
rect 122 219 280 253
rect 316 253 436 269
rect 316 235 386 253
rect 18 153 280 219
rect 18 119 88 153
rect 122 119 280 153
rect 18 113 280 119
rect 18 79 24 113
rect 58 79 96 113
rect 130 79 168 113
rect 202 79 240 113
rect 274 79 280 113
rect 370 219 386 235
rect 420 219 436 253
rect 370 153 436 219
rect 370 119 386 153
rect 420 119 436 153
rect 370 103 436 119
rect 18 73 280 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 24 701 58 735
rect 96 701 122 735
rect 122 701 130 735
rect 168 701 202 735
rect 338 701 372 735
rect 410 701 434 735
rect 434 701 444 735
rect 24 79 58 113
rect 96 79 130 113
rect 168 79 202 113
rect 240 79 274 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 831 480 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 480 831
rect 0 791 480 797
rect 0 735 480 763
rect 0 701 24 735
rect 58 701 96 735
rect 130 701 168 735
rect 202 701 338 735
rect 372 701 410 735
rect 444 701 480 735
rect 0 689 480 701
rect 0 113 480 125
rect 0 79 24 113
rect 58 79 96 113
rect 130 79 168 113
rect 202 79 240 113
rect 274 79 480 113
rect 0 51 480 79
rect 0 17 480 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -23 480 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand2_1
flabel metal1 s 0 51 480 125 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 0 480 23 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 0 689 480 763 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 791 480 814 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 480 814
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string LEFsymmetry X Y
string GDS_END 709384
string GDS_START 702626
<< end >>
