magic
tech sky130A
magscale 1 2
timestamp 1640697980
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 37 67 504 203
rect 37 21 407 67
rect 37 17 63 21
rect 29 -17 63 17
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 17 289 109 491
rect 323 425 389 527
rect 17 165 51 289
rect 213 199 261 323
rect 295 199 363 323
rect 397 199 467 323
rect 17 131 289 165
rect 17 51 121 131
rect 155 17 221 97
rect 255 62 289 131
rect 323 17 389 165
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< obsli1 >>
rect 143 357 535 391
rect 143 249 177 357
rect 85 215 177 249
rect 501 165 535 357
rect 436 131 535 165
rect 436 81 470 131
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 295 199 363 323 6 A
port 1 nsew signal input
rlabel locali s 213 199 261 323 6 B
port 2 nsew signal input
rlabel locali s 397 199 467 323 6 C_N
port 3 nsew signal input
rlabel metal1 s 0 -48 552 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 489 -17 523 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 397 -17 431 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 305 -17 339 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 213 -17 247 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 121 -17 155 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel viali s 29 -17 63 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 552 17 8 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 323 17 389 165 6 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 155 17 221 97 6 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s 37 17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 37 21 407 67 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 37 67 504 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 590 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 489 527 523 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 397 527 431 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 305 527 339 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 213 527 247 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 121 527 155 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel viali s 29 527 63 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 323 425 389 527 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 552 561 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 255 62 289 131 6 Y
port 8 nsew signal output
rlabel locali s 17 51 121 131 6 Y
port 8 nsew signal output
rlabel locali s 17 131 289 165 6 Y
port 8 nsew signal output
rlabel locali s 17 165 51 289 6 Y
port 8 nsew signal output
rlabel locali s 17 289 109 491 6 Y
port 8 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 552 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1128596
string GDS_START 1123852
<< end >>
