magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect 10461 367 39030 17423
<< nwell >>
rect 35513 13137 37645 15191
rect 13104 2287 15158 2497
rect 12349 2212 15158 2287
rect 12349 2006 15303 2212
rect 11967 1823 15303 2006
rect 11967 1790 15861 1823
rect 11997 1657 15861 1790
<< pwell >>
rect 11721 3640 14647 3674
rect 12520 2566 12880 2600
rect 18139 1657 23641 1691
<< mvnmos >>
rect 11794 2966 11894 3566
rect 11950 2966 12050 3566
rect 12106 2966 12206 3566
rect 12262 2966 12362 3566
rect 12418 2966 12518 3566
rect 12574 2966 12674 3566
rect 12730 2966 12830 3566
rect 12886 2966 12986 3566
rect 13042 2966 13142 3566
rect 13198 2966 13298 3566
rect 13354 2966 13454 3566
rect 13510 2966 13610 3566
rect 13787 2966 13907 3566
rect 14087 2966 14207 3566
rect 14263 2966 14363 3566
rect 14419 2966 14519 3566
rect 12468 2408 12668 2492
rect 12724 2408 12924 2492
<< mvpmos >>
rect 35579 14972 37579 15072
rect 35579 14816 37579 14916
rect 35579 14660 37579 14760
rect 35579 14504 37579 14604
rect 35579 14348 37579 14448
rect 35579 14192 37579 14292
rect 35579 14036 37579 14136
rect 35579 13880 37579 13980
rect 35579 13724 37579 13824
rect 35579 13568 37579 13668
rect 35579 13412 37579 13512
rect 35579 13256 37579 13356
rect 12468 2137 12668 2221
rect 12724 2137 12924 2221
rect 12086 1856 12486 1940
rect 12542 1856 12942 1940
rect 13223 1831 13323 2431
rect 13379 1831 13479 2431
rect 13535 1831 13635 2431
rect 13691 1831 13791 2431
rect 13847 1831 13947 2431
rect 14003 1831 14103 2431
rect 14159 1831 14259 2431
rect 14315 1831 14415 2431
rect 14471 1831 14571 2431
rect 14627 1831 14727 2431
rect 14783 1831 14883 2431
rect 14939 1831 15039 2431
<< mvndiff >>
rect 11741 3554 11794 3566
rect 11741 3520 11749 3554
rect 11783 3520 11794 3554
rect 11741 3486 11794 3520
rect 11741 3452 11749 3486
rect 11783 3452 11794 3486
rect 11741 3418 11794 3452
rect 11741 3384 11749 3418
rect 11783 3384 11794 3418
rect 11741 3350 11794 3384
rect 11741 3316 11749 3350
rect 11783 3316 11794 3350
rect 11741 3282 11794 3316
rect 11741 3248 11749 3282
rect 11783 3248 11794 3282
rect 11741 3214 11794 3248
rect 11741 3180 11749 3214
rect 11783 3180 11794 3214
rect 11741 3146 11794 3180
rect 11741 3112 11749 3146
rect 11783 3112 11794 3146
rect 11741 3078 11794 3112
rect 11741 3044 11749 3078
rect 11783 3044 11794 3078
rect 11741 2966 11794 3044
rect 11894 3554 11950 3566
rect 11894 3520 11905 3554
rect 11939 3520 11950 3554
rect 11894 3486 11950 3520
rect 11894 3452 11905 3486
rect 11939 3452 11950 3486
rect 11894 3418 11950 3452
rect 11894 3384 11905 3418
rect 11939 3384 11950 3418
rect 11894 3350 11950 3384
rect 11894 3316 11905 3350
rect 11939 3316 11950 3350
rect 11894 3282 11950 3316
rect 11894 3248 11905 3282
rect 11939 3248 11950 3282
rect 11894 3214 11950 3248
rect 11894 3180 11905 3214
rect 11939 3180 11950 3214
rect 11894 3146 11950 3180
rect 11894 3112 11905 3146
rect 11939 3112 11950 3146
rect 11894 3078 11950 3112
rect 11894 3044 11905 3078
rect 11939 3044 11950 3078
rect 11894 2966 11950 3044
rect 12050 3554 12106 3566
rect 12050 3520 12061 3554
rect 12095 3520 12106 3554
rect 12050 3486 12106 3520
rect 12050 3452 12061 3486
rect 12095 3452 12106 3486
rect 12050 3418 12106 3452
rect 12050 3384 12061 3418
rect 12095 3384 12106 3418
rect 12050 3350 12106 3384
rect 12050 3316 12061 3350
rect 12095 3316 12106 3350
rect 12050 3282 12106 3316
rect 12050 3248 12061 3282
rect 12095 3248 12106 3282
rect 12050 3214 12106 3248
rect 12050 3180 12061 3214
rect 12095 3180 12106 3214
rect 12050 3146 12106 3180
rect 12050 3112 12061 3146
rect 12095 3112 12106 3146
rect 12050 3078 12106 3112
rect 12050 3044 12061 3078
rect 12095 3044 12106 3078
rect 12050 2966 12106 3044
rect 12206 3554 12262 3566
rect 12206 3520 12217 3554
rect 12251 3520 12262 3554
rect 12206 3486 12262 3520
rect 12206 3452 12217 3486
rect 12251 3452 12262 3486
rect 12206 3418 12262 3452
rect 12206 3384 12217 3418
rect 12251 3384 12262 3418
rect 12206 3350 12262 3384
rect 12206 3316 12217 3350
rect 12251 3316 12262 3350
rect 12206 3282 12262 3316
rect 12206 3248 12217 3282
rect 12251 3248 12262 3282
rect 12206 3214 12262 3248
rect 12206 3180 12217 3214
rect 12251 3180 12262 3214
rect 12206 3146 12262 3180
rect 12206 3112 12217 3146
rect 12251 3112 12262 3146
rect 12206 3078 12262 3112
rect 12206 3044 12217 3078
rect 12251 3044 12262 3078
rect 12206 2966 12262 3044
rect 12362 3554 12418 3566
rect 12362 3520 12373 3554
rect 12407 3520 12418 3554
rect 12362 3486 12418 3520
rect 12362 3452 12373 3486
rect 12407 3452 12418 3486
rect 12362 3418 12418 3452
rect 12362 3384 12373 3418
rect 12407 3384 12418 3418
rect 12362 3350 12418 3384
rect 12362 3316 12373 3350
rect 12407 3316 12418 3350
rect 12362 3282 12418 3316
rect 12362 3248 12373 3282
rect 12407 3248 12418 3282
rect 12362 3214 12418 3248
rect 12362 3180 12373 3214
rect 12407 3180 12418 3214
rect 12362 3146 12418 3180
rect 12362 3112 12373 3146
rect 12407 3112 12418 3146
rect 12362 3078 12418 3112
rect 12362 3044 12373 3078
rect 12407 3044 12418 3078
rect 12362 2966 12418 3044
rect 12518 3554 12574 3566
rect 12518 3520 12529 3554
rect 12563 3520 12574 3554
rect 12518 3486 12574 3520
rect 12518 3452 12529 3486
rect 12563 3452 12574 3486
rect 12518 3418 12574 3452
rect 12518 3384 12529 3418
rect 12563 3384 12574 3418
rect 12518 3350 12574 3384
rect 12518 3316 12529 3350
rect 12563 3316 12574 3350
rect 12518 3282 12574 3316
rect 12518 3248 12529 3282
rect 12563 3248 12574 3282
rect 12518 3214 12574 3248
rect 12518 3180 12529 3214
rect 12563 3180 12574 3214
rect 12518 3146 12574 3180
rect 12518 3112 12529 3146
rect 12563 3112 12574 3146
rect 12518 3078 12574 3112
rect 12518 3044 12529 3078
rect 12563 3044 12574 3078
rect 12518 2966 12574 3044
rect 12674 3554 12730 3566
rect 12674 3520 12685 3554
rect 12719 3520 12730 3554
rect 12674 3486 12730 3520
rect 12674 3452 12685 3486
rect 12719 3452 12730 3486
rect 12674 3418 12730 3452
rect 12674 3384 12685 3418
rect 12719 3384 12730 3418
rect 12674 3350 12730 3384
rect 12674 3316 12685 3350
rect 12719 3316 12730 3350
rect 12674 3282 12730 3316
rect 12674 3248 12685 3282
rect 12719 3248 12730 3282
rect 12674 3214 12730 3248
rect 12674 3180 12685 3214
rect 12719 3180 12730 3214
rect 12674 3146 12730 3180
rect 12674 3112 12685 3146
rect 12719 3112 12730 3146
rect 12674 3078 12730 3112
rect 12674 3044 12685 3078
rect 12719 3044 12730 3078
rect 12674 2966 12730 3044
rect 12830 3554 12886 3566
rect 12830 3520 12841 3554
rect 12875 3520 12886 3554
rect 12830 3486 12886 3520
rect 12830 3452 12841 3486
rect 12875 3452 12886 3486
rect 12830 3418 12886 3452
rect 12830 3384 12841 3418
rect 12875 3384 12886 3418
rect 12830 3350 12886 3384
rect 12830 3316 12841 3350
rect 12875 3316 12886 3350
rect 12830 3282 12886 3316
rect 12830 3248 12841 3282
rect 12875 3248 12886 3282
rect 12830 3214 12886 3248
rect 12830 3180 12841 3214
rect 12875 3180 12886 3214
rect 12830 3146 12886 3180
rect 12830 3112 12841 3146
rect 12875 3112 12886 3146
rect 12830 3078 12886 3112
rect 12830 3044 12841 3078
rect 12875 3044 12886 3078
rect 12830 2966 12886 3044
rect 12986 3554 13042 3566
rect 12986 3520 12997 3554
rect 13031 3520 13042 3554
rect 12986 3486 13042 3520
rect 12986 3452 12997 3486
rect 13031 3452 13042 3486
rect 12986 3418 13042 3452
rect 12986 3384 12997 3418
rect 13031 3384 13042 3418
rect 12986 3350 13042 3384
rect 12986 3316 12997 3350
rect 13031 3316 13042 3350
rect 12986 3282 13042 3316
rect 12986 3248 12997 3282
rect 13031 3248 13042 3282
rect 12986 3214 13042 3248
rect 12986 3180 12997 3214
rect 13031 3180 13042 3214
rect 12986 3146 13042 3180
rect 12986 3112 12997 3146
rect 13031 3112 13042 3146
rect 12986 3078 13042 3112
rect 12986 3044 12997 3078
rect 13031 3044 13042 3078
rect 12986 2966 13042 3044
rect 13142 3554 13198 3566
rect 13142 3520 13153 3554
rect 13187 3520 13198 3554
rect 13142 3486 13198 3520
rect 13142 3452 13153 3486
rect 13187 3452 13198 3486
rect 13142 3418 13198 3452
rect 13142 3384 13153 3418
rect 13187 3384 13198 3418
rect 13142 3350 13198 3384
rect 13142 3316 13153 3350
rect 13187 3316 13198 3350
rect 13142 3282 13198 3316
rect 13142 3248 13153 3282
rect 13187 3248 13198 3282
rect 13142 3214 13198 3248
rect 13142 3180 13153 3214
rect 13187 3180 13198 3214
rect 13142 3146 13198 3180
rect 13142 3112 13153 3146
rect 13187 3112 13198 3146
rect 13142 3078 13198 3112
rect 13142 3044 13153 3078
rect 13187 3044 13198 3078
rect 13142 2966 13198 3044
rect 13298 3554 13354 3566
rect 13298 3520 13309 3554
rect 13343 3520 13354 3554
rect 13298 3486 13354 3520
rect 13298 3452 13309 3486
rect 13343 3452 13354 3486
rect 13298 3418 13354 3452
rect 13298 3384 13309 3418
rect 13343 3384 13354 3418
rect 13298 3350 13354 3384
rect 13298 3316 13309 3350
rect 13343 3316 13354 3350
rect 13298 3282 13354 3316
rect 13298 3248 13309 3282
rect 13343 3248 13354 3282
rect 13298 3214 13354 3248
rect 13298 3180 13309 3214
rect 13343 3180 13354 3214
rect 13298 3146 13354 3180
rect 13298 3112 13309 3146
rect 13343 3112 13354 3146
rect 13298 3078 13354 3112
rect 13298 3044 13309 3078
rect 13343 3044 13354 3078
rect 13298 2966 13354 3044
rect 13454 3554 13510 3566
rect 13454 3520 13465 3554
rect 13499 3520 13510 3554
rect 13454 3486 13510 3520
rect 13454 3452 13465 3486
rect 13499 3452 13510 3486
rect 13454 3418 13510 3452
rect 13454 3384 13465 3418
rect 13499 3384 13510 3418
rect 13454 3350 13510 3384
rect 13454 3316 13465 3350
rect 13499 3316 13510 3350
rect 13454 3282 13510 3316
rect 13454 3248 13465 3282
rect 13499 3248 13510 3282
rect 13454 3214 13510 3248
rect 13454 3180 13465 3214
rect 13499 3180 13510 3214
rect 13454 3146 13510 3180
rect 13454 3112 13465 3146
rect 13499 3112 13510 3146
rect 13454 3078 13510 3112
rect 13454 3044 13465 3078
rect 13499 3044 13510 3078
rect 13454 2966 13510 3044
rect 13610 3554 13663 3566
rect 13610 3520 13621 3554
rect 13655 3520 13663 3554
rect 13610 3486 13663 3520
rect 13610 3452 13621 3486
rect 13655 3452 13663 3486
rect 13610 3418 13663 3452
rect 13610 3384 13621 3418
rect 13655 3384 13663 3418
rect 13610 3350 13663 3384
rect 13610 3316 13621 3350
rect 13655 3316 13663 3350
rect 13610 3282 13663 3316
rect 13610 3248 13621 3282
rect 13655 3248 13663 3282
rect 13610 3214 13663 3248
rect 13610 3180 13621 3214
rect 13655 3180 13663 3214
rect 13610 3146 13663 3180
rect 13610 3112 13621 3146
rect 13655 3112 13663 3146
rect 13610 3078 13663 3112
rect 13610 3044 13621 3078
rect 13655 3044 13663 3078
rect 13610 2966 13663 3044
rect 13734 3554 13787 3566
rect 13734 3520 13742 3554
rect 13776 3520 13787 3554
rect 13734 3486 13787 3520
rect 13734 3452 13742 3486
rect 13776 3452 13787 3486
rect 13734 3418 13787 3452
rect 13734 3384 13742 3418
rect 13776 3384 13787 3418
rect 13734 3350 13787 3384
rect 13734 3316 13742 3350
rect 13776 3316 13787 3350
rect 13734 3282 13787 3316
rect 13734 3248 13742 3282
rect 13776 3248 13787 3282
rect 13734 3214 13787 3248
rect 13734 3180 13742 3214
rect 13776 3180 13787 3214
rect 13734 3146 13787 3180
rect 13734 3112 13742 3146
rect 13776 3112 13787 3146
rect 13734 3078 13787 3112
rect 13734 3044 13742 3078
rect 13776 3044 13787 3078
rect 13734 2966 13787 3044
rect 13907 3554 13960 3566
rect 13907 3520 13918 3554
rect 13952 3520 13960 3554
rect 13907 3486 13960 3520
rect 13907 3452 13918 3486
rect 13952 3452 13960 3486
rect 13907 3418 13960 3452
rect 13907 3384 13918 3418
rect 13952 3384 13960 3418
rect 13907 3350 13960 3384
rect 13907 3316 13918 3350
rect 13952 3316 13960 3350
rect 13907 3282 13960 3316
rect 13907 3248 13918 3282
rect 13952 3248 13960 3282
rect 13907 3214 13960 3248
rect 13907 3180 13918 3214
rect 13952 3180 13960 3214
rect 13907 3146 13960 3180
rect 13907 3112 13918 3146
rect 13952 3112 13960 3146
rect 13907 3078 13960 3112
rect 13907 3044 13918 3078
rect 13952 3044 13960 3078
rect 13907 2966 13960 3044
rect 14034 3554 14087 3566
rect 14034 3520 14042 3554
rect 14076 3520 14087 3554
rect 14034 3486 14087 3520
rect 14034 3452 14042 3486
rect 14076 3452 14087 3486
rect 14034 3418 14087 3452
rect 14034 3384 14042 3418
rect 14076 3384 14087 3418
rect 14034 3350 14087 3384
rect 14034 3316 14042 3350
rect 14076 3316 14087 3350
rect 14034 3282 14087 3316
rect 14034 3248 14042 3282
rect 14076 3248 14087 3282
rect 14034 3214 14087 3248
rect 14034 3180 14042 3214
rect 14076 3180 14087 3214
rect 14034 3146 14087 3180
rect 14034 3112 14042 3146
rect 14076 3112 14087 3146
rect 14034 3078 14087 3112
rect 14034 3044 14042 3078
rect 14076 3044 14087 3078
rect 14034 2966 14087 3044
rect 14207 3554 14263 3566
rect 14207 3520 14218 3554
rect 14252 3520 14263 3554
rect 14207 3486 14263 3520
rect 14207 3452 14218 3486
rect 14252 3452 14263 3486
rect 14207 3418 14263 3452
rect 14207 3384 14218 3418
rect 14252 3384 14263 3418
rect 14207 3350 14263 3384
rect 14207 3316 14218 3350
rect 14252 3316 14263 3350
rect 14207 3282 14263 3316
rect 14207 3248 14218 3282
rect 14252 3248 14263 3282
rect 14207 3214 14263 3248
rect 14207 3180 14218 3214
rect 14252 3180 14263 3214
rect 14207 3146 14263 3180
rect 14207 3112 14218 3146
rect 14252 3112 14263 3146
rect 14207 3078 14263 3112
rect 14207 3044 14218 3078
rect 14252 3044 14263 3078
rect 14207 2966 14263 3044
rect 14363 3554 14419 3566
rect 14363 3520 14374 3554
rect 14408 3520 14419 3554
rect 14363 3486 14419 3520
rect 14363 3452 14374 3486
rect 14408 3452 14419 3486
rect 14363 3418 14419 3452
rect 14363 3384 14374 3418
rect 14408 3384 14419 3418
rect 14363 3350 14419 3384
rect 14363 3316 14374 3350
rect 14408 3316 14419 3350
rect 14363 3282 14419 3316
rect 14363 3248 14374 3282
rect 14408 3248 14419 3282
rect 14363 3214 14419 3248
rect 14363 3180 14374 3214
rect 14408 3180 14419 3214
rect 14363 3146 14419 3180
rect 14363 3112 14374 3146
rect 14408 3112 14419 3146
rect 14363 3078 14419 3112
rect 14363 3044 14374 3078
rect 14408 3044 14419 3078
rect 14363 2966 14419 3044
rect 14519 3554 14572 3566
rect 14519 3520 14530 3554
rect 14564 3520 14572 3554
rect 14519 3486 14572 3520
rect 14519 3452 14530 3486
rect 14564 3452 14572 3486
rect 14519 3418 14572 3452
rect 14519 3384 14530 3418
rect 14564 3384 14572 3418
rect 14519 3350 14572 3384
rect 14519 3316 14530 3350
rect 14564 3316 14572 3350
rect 14519 3282 14572 3316
rect 14519 3248 14530 3282
rect 14564 3248 14572 3282
rect 14519 3214 14572 3248
rect 14519 3180 14530 3214
rect 14564 3180 14572 3214
rect 14519 3146 14572 3180
rect 14519 3112 14530 3146
rect 14564 3112 14572 3146
rect 14519 3078 14572 3112
rect 14519 3044 14530 3078
rect 14564 3044 14572 3078
rect 14519 2966 14572 3044
rect 12415 2480 12468 2492
rect 12415 2446 12423 2480
rect 12457 2446 12468 2480
rect 12415 2408 12468 2446
rect 12668 2480 12724 2492
rect 12668 2446 12679 2480
rect 12713 2446 12724 2480
rect 12668 2408 12724 2446
rect 12924 2480 12977 2492
rect 12924 2446 12935 2480
rect 12969 2446 12977 2480
rect 12924 2408 12977 2446
<< mvpdiff >>
rect 35579 15117 37579 15125
rect 35579 15083 35591 15117
rect 35625 15083 35659 15117
rect 35693 15083 35727 15117
rect 35761 15083 35795 15117
rect 35829 15083 35863 15117
rect 35897 15083 35931 15117
rect 35965 15083 35999 15117
rect 36033 15083 36067 15117
rect 36101 15083 36135 15117
rect 36169 15083 36203 15117
rect 36237 15083 36271 15117
rect 36305 15083 36339 15117
rect 36373 15083 36407 15117
rect 36441 15083 36475 15117
rect 36509 15083 36543 15117
rect 36577 15083 36611 15117
rect 36645 15083 36679 15117
rect 36713 15083 36747 15117
rect 36781 15083 36815 15117
rect 36849 15083 36883 15117
rect 36917 15083 36951 15117
rect 36985 15083 37019 15117
rect 37053 15083 37087 15117
rect 37121 15083 37155 15117
rect 37189 15083 37223 15117
rect 37257 15083 37291 15117
rect 37325 15083 37359 15117
rect 37393 15083 37427 15117
rect 37461 15083 37495 15117
rect 37529 15083 37579 15117
rect 35579 15072 37579 15083
rect 35579 14961 37579 14972
rect 35579 14927 35591 14961
rect 35625 14927 35659 14961
rect 35693 14927 35727 14961
rect 35761 14927 35795 14961
rect 35829 14927 35863 14961
rect 35897 14927 35931 14961
rect 35965 14927 35999 14961
rect 36033 14927 36067 14961
rect 36101 14927 36135 14961
rect 36169 14927 36203 14961
rect 36237 14927 36271 14961
rect 36305 14927 36339 14961
rect 36373 14927 36407 14961
rect 36441 14927 36475 14961
rect 36509 14927 36543 14961
rect 36577 14927 36611 14961
rect 36645 14927 36679 14961
rect 36713 14927 36747 14961
rect 36781 14927 36815 14961
rect 36849 14927 36883 14961
rect 36917 14927 36951 14961
rect 36985 14927 37019 14961
rect 37053 14927 37087 14961
rect 37121 14927 37155 14961
rect 37189 14927 37223 14961
rect 37257 14927 37291 14961
rect 37325 14927 37359 14961
rect 37393 14927 37427 14961
rect 37461 14927 37495 14961
rect 37529 14927 37579 14961
rect 35579 14916 37579 14927
rect 35579 14805 37579 14816
rect 35579 14771 35591 14805
rect 35625 14771 35659 14805
rect 35693 14771 35727 14805
rect 35761 14771 35795 14805
rect 35829 14771 35863 14805
rect 35897 14771 35931 14805
rect 35965 14771 35999 14805
rect 36033 14771 36067 14805
rect 36101 14771 36135 14805
rect 36169 14771 36203 14805
rect 36237 14771 36271 14805
rect 36305 14771 36339 14805
rect 36373 14771 36407 14805
rect 36441 14771 36475 14805
rect 36509 14771 36543 14805
rect 36577 14771 36611 14805
rect 36645 14771 36679 14805
rect 36713 14771 36747 14805
rect 36781 14771 36815 14805
rect 36849 14771 36883 14805
rect 36917 14771 36951 14805
rect 36985 14771 37019 14805
rect 37053 14771 37087 14805
rect 37121 14771 37155 14805
rect 37189 14771 37223 14805
rect 37257 14771 37291 14805
rect 37325 14771 37359 14805
rect 37393 14771 37427 14805
rect 37461 14771 37495 14805
rect 37529 14771 37579 14805
rect 35579 14760 37579 14771
rect 35579 14649 37579 14660
rect 35579 14615 35591 14649
rect 35625 14615 35659 14649
rect 35693 14615 35727 14649
rect 35761 14615 35795 14649
rect 35829 14615 35863 14649
rect 35897 14615 35931 14649
rect 35965 14615 35999 14649
rect 36033 14615 36067 14649
rect 36101 14615 36135 14649
rect 36169 14615 36203 14649
rect 36237 14615 36271 14649
rect 36305 14615 36339 14649
rect 36373 14615 36407 14649
rect 36441 14615 36475 14649
rect 36509 14615 36543 14649
rect 36577 14615 36611 14649
rect 36645 14615 36679 14649
rect 36713 14615 36747 14649
rect 36781 14615 36815 14649
rect 36849 14615 36883 14649
rect 36917 14615 36951 14649
rect 36985 14615 37019 14649
rect 37053 14615 37087 14649
rect 37121 14615 37155 14649
rect 37189 14615 37223 14649
rect 37257 14615 37291 14649
rect 37325 14615 37359 14649
rect 37393 14615 37427 14649
rect 37461 14615 37495 14649
rect 37529 14615 37579 14649
rect 35579 14604 37579 14615
rect 35579 14493 37579 14504
rect 35579 14459 35591 14493
rect 35625 14459 35659 14493
rect 35693 14459 35727 14493
rect 35761 14459 35795 14493
rect 35829 14459 35863 14493
rect 35897 14459 35931 14493
rect 35965 14459 35999 14493
rect 36033 14459 36067 14493
rect 36101 14459 36135 14493
rect 36169 14459 36203 14493
rect 36237 14459 36271 14493
rect 36305 14459 36339 14493
rect 36373 14459 36407 14493
rect 36441 14459 36475 14493
rect 36509 14459 36543 14493
rect 36577 14459 36611 14493
rect 36645 14459 36679 14493
rect 36713 14459 36747 14493
rect 36781 14459 36815 14493
rect 36849 14459 36883 14493
rect 36917 14459 36951 14493
rect 36985 14459 37019 14493
rect 37053 14459 37087 14493
rect 37121 14459 37155 14493
rect 37189 14459 37223 14493
rect 37257 14459 37291 14493
rect 37325 14459 37359 14493
rect 37393 14459 37427 14493
rect 37461 14459 37495 14493
rect 37529 14459 37579 14493
rect 35579 14448 37579 14459
rect 35579 14337 37579 14348
rect 35579 14303 35591 14337
rect 35625 14303 35659 14337
rect 35693 14303 35727 14337
rect 35761 14303 35795 14337
rect 35829 14303 35863 14337
rect 35897 14303 35931 14337
rect 35965 14303 35999 14337
rect 36033 14303 36067 14337
rect 36101 14303 36135 14337
rect 36169 14303 36203 14337
rect 36237 14303 36271 14337
rect 36305 14303 36339 14337
rect 36373 14303 36407 14337
rect 36441 14303 36475 14337
rect 36509 14303 36543 14337
rect 36577 14303 36611 14337
rect 36645 14303 36679 14337
rect 36713 14303 36747 14337
rect 36781 14303 36815 14337
rect 36849 14303 36883 14337
rect 36917 14303 36951 14337
rect 36985 14303 37019 14337
rect 37053 14303 37087 14337
rect 37121 14303 37155 14337
rect 37189 14303 37223 14337
rect 37257 14303 37291 14337
rect 37325 14303 37359 14337
rect 37393 14303 37427 14337
rect 37461 14303 37495 14337
rect 37529 14303 37579 14337
rect 35579 14292 37579 14303
rect 35579 14181 37579 14192
rect 35579 14147 35591 14181
rect 35625 14147 35659 14181
rect 35693 14147 35727 14181
rect 35761 14147 35795 14181
rect 35829 14147 35863 14181
rect 35897 14147 35931 14181
rect 35965 14147 35999 14181
rect 36033 14147 36067 14181
rect 36101 14147 36135 14181
rect 36169 14147 36203 14181
rect 36237 14147 36271 14181
rect 36305 14147 36339 14181
rect 36373 14147 36407 14181
rect 36441 14147 36475 14181
rect 36509 14147 36543 14181
rect 36577 14147 36611 14181
rect 36645 14147 36679 14181
rect 36713 14147 36747 14181
rect 36781 14147 36815 14181
rect 36849 14147 36883 14181
rect 36917 14147 36951 14181
rect 36985 14147 37019 14181
rect 37053 14147 37087 14181
rect 37121 14147 37155 14181
rect 37189 14147 37223 14181
rect 37257 14147 37291 14181
rect 37325 14147 37359 14181
rect 37393 14147 37427 14181
rect 37461 14147 37495 14181
rect 37529 14147 37579 14181
rect 35579 14136 37579 14147
rect 35579 14025 37579 14036
rect 35579 13991 35591 14025
rect 35625 13991 35659 14025
rect 35693 13991 35727 14025
rect 35761 13991 35795 14025
rect 35829 13991 35863 14025
rect 35897 13991 35931 14025
rect 35965 13991 35999 14025
rect 36033 13991 36067 14025
rect 36101 13991 36135 14025
rect 36169 13991 36203 14025
rect 36237 13991 36271 14025
rect 36305 13991 36339 14025
rect 36373 13991 36407 14025
rect 36441 13991 36475 14025
rect 36509 13991 36543 14025
rect 36577 13991 36611 14025
rect 36645 13991 36679 14025
rect 36713 13991 36747 14025
rect 36781 13991 36815 14025
rect 36849 13991 36883 14025
rect 36917 13991 36951 14025
rect 36985 13991 37019 14025
rect 37053 13991 37087 14025
rect 37121 13991 37155 14025
rect 37189 13991 37223 14025
rect 37257 13991 37291 14025
rect 37325 13991 37359 14025
rect 37393 13991 37427 14025
rect 37461 13991 37495 14025
rect 37529 13991 37579 14025
rect 35579 13980 37579 13991
rect 35579 13869 37579 13880
rect 35579 13835 35591 13869
rect 35625 13835 35659 13869
rect 35693 13835 35727 13869
rect 35761 13835 35795 13869
rect 35829 13835 35863 13869
rect 35897 13835 35931 13869
rect 35965 13835 35999 13869
rect 36033 13835 36067 13869
rect 36101 13835 36135 13869
rect 36169 13835 36203 13869
rect 36237 13835 36271 13869
rect 36305 13835 36339 13869
rect 36373 13835 36407 13869
rect 36441 13835 36475 13869
rect 36509 13835 36543 13869
rect 36577 13835 36611 13869
rect 36645 13835 36679 13869
rect 36713 13835 36747 13869
rect 36781 13835 36815 13869
rect 36849 13835 36883 13869
rect 36917 13835 36951 13869
rect 36985 13835 37019 13869
rect 37053 13835 37087 13869
rect 37121 13835 37155 13869
rect 37189 13835 37223 13869
rect 37257 13835 37291 13869
rect 37325 13835 37359 13869
rect 37393 13835 37427 13869
rect 37461 13835 37495 13869
rect 37529 13835 37579 13869
rect 35579 13824 37579 13835
rect 35579 13713 37579 13724
rect 35579 13679 35591 13713
rect 35625 13679 35659 13713
rect 35693 13679 35727 13713
rect 35761 13679 35795 13713
rect 35829 13679 35863 13713
rect 35897 13679 35931 13713
rect 35965 13679 35999 13713
rect 36033 13679 36067 13713
rect 36101 13679 36135 13713
rect 36169 13679 36203 13713
rect 36237 13679 36271 13713
rect 36305 13679 36339 13713
rect 36373 13679 36407 13713
rect 36441 13679 36475 13713
rect 36509 13679 36543 13713
rect 36577 13679 36611 13713
rect 36645 13679 36679 13713
rect 36713 13679 36747 13713
rect 36781 13679 36815 13713
rect 36849 13679 36883 13713
rect 36917 13679 36951 13713
rect 36985 13679 37019 13713
rect 37053 13679 37087 13713
rect 37121 13679 37155 13713
rect 37189 13679 37223 13713
rect 37257 13679 37291 13713
rect 37325 13679 37359 13713
rect 37393 13679 37427 13713
rect 37461 13679 37495 13713
rect 37529 13679 37579 13713
rect 35579 13668 37579 13679
rect 35579 13557 37579 13568
rect 35579 13523 35591 13557
rect 35625 13523 35659 13557
rect 35693 13523 35727 13557
rect 35761 13523 35795 13557
rect 35829 13523 35863 13557
rect 35897 13523 35931 13557
rect 35965 13523 35999 13557
rect 36033 13523 36067 13557
rect 36101 13523 36135 13557
rect 36169 13523 36203 13557
rect 36237 13523 36271 13557
rect 36305 13523 36339 13557
rect 36373 13523 36407 13557
rect 36441 13523 36475 13557
rect 36509 13523 36543 13557
rect 36577 13523 36611 13557
rect 36645 13523 36679 13557
rect 36713 13523 36747 13557
rect 36781 13523 36815 13557
rect 36849 13523 36883 13557
rect 36917 13523 36951 13557
rect 36985 13523 37019 13557
rect 37053 13523 37087 13557
rect 37121 13523 37155 13557
rect 37189 13523 37223 13557
rect 37257 13523 37291 13557
rect 37325 13523 37359 13557
rect 37393 13523 37427 13557
rect 37461 13523 37495 13557
rect 37529 13523 37579 13557
rect 35579 13512 37579 13523
rect 35579 13401 37579 13412
rect 35579 13367 35591 13401
rect 35625 13367 35659 13401
rect 35693 13367 35727 13401
rect 35761 13367 35795 13401
rect 35829 13367 35863 13401
rect 35897 13367 35931 13401
rect 35965 13367 35999 13401
rect 36033 13367 36067 13401
rect 36101 13367 36135 13401
rect 36169 13367 36203 13401
rect 36237 13367 36271 13401
rect 36305 13367 36339 13401
rect 36373 13367 36407 13401
rect 36441 13367 36475 13401
rect 36509 13367 36543 13401
rect 36577 13367 36611 13401
rect 36645 13367 36679 13401
rect 36713 13367 36747 13401
rect 36781 13367 36815 13401
rect 36849 13367 36883 13401
rect 36917 13367 36951 13401
rect 36985 13367 37019 13401
rect 37053 13367 37087 13401
rect 37121 13367 37155 13401
rect 37189 13367 37223 13401
rect 37257 13367 37291 13401
rect 37325 13367 37359 13401
rect 37393 13367 37427 13401
rect 37461 13367 37495 13401
rect 37529 13367 37579 13401
rect 35579 13356 37579 13367
rect 35579 13245 37579 13256
rect 35579 13211 35591 13245
rect 35625 13211 35659 13245
rect 35693 13211 35727 13245
rect 35761 13211 35795 13245
rect 35829 13211 35863 13245
rect 35897 13211 35931 13245
rect 35965 13211 35999 13245
rect 36033 13211 36067 13245
rect 36101 13211 36135 13245
rect 36169 13211 36203 13245
rect 36237 13211 36271 13245
rect 36305 13211 36339 13245
rect 36373 13211 36407 13245
rect 36441 13211 36475 13245
rect 36509 13211 36543 13245
rect 36577 13211 36611 13245
rect 36645 13211 36679 13245
rect 36713 13211 36747 13245
rect 36781 13211 36815 13245
rect 36849 13211 36883 13245
rect 36917 13211 36951 13245
rect 36985 13211 37019 13245
rect 37053 13211 37087 13245
rect 37121 13211 37155 13245
rect 37189 13211 37223 13245
rect 37257 13211 37291 13245
rect 37325 13211 37359 13245
rect 37393 13211 37427 13245
rect 37461 13211 37495 13245
rect 37529 13211 37579 13245
rect 35579 13203 37579 13211
rect 13170 2353 13223 2431
rect 13170 2319 13178 2353
rect 13212 2319 13223 2353
rect 13170 2285 13223 2319
rect 13170 2251 13178 2285
rect 13212 2251 13223 2285
rect 12415 2183 12468 2221
rect 12415 2149 12423 2183
rect 12457 2149 12468 2183
rect 12415 2137 12468 2149
rect 12668 2183 12724 2221
rect 12668 2149 12679 2183
rect 12713 2149 12724 2183
rect 12668 2137 12724 2149
rect 12924 2183 12977 2221
rect 12924 2149 12935 2183
rect 12969 2149 12977 2183
rect 12924 2137 12977 2149
rect 13170 2217 13223 2251
rect 13170 2183 13178 2217
rect 13212 2183 13223 2217
rect 13170 2149 13223 2183
rect 13170 2115 13178 2149
rect 13212 2115 13223 2149
rect 13170 2081 13223 2115
rect 13170 2047 13178 2081
rect 13212 2047 13223 2081
rect 13170 2013 13223 2047
rect 13170 1979 13178 2013
rect 13212 1979 13223 2013
rect 13170 1945 13223 1979
rect 12033 1928 12086 1940
rect 12033 1894 12041 1928
rect 12075 1894 12086 1928
rect 12033 1856 12086 1894
rect 12486 1928 12542 1940
rect 12486 1894 12497 1928
rect 12531 1894 12542 1928
rect 12486 1856 12542 1894
rect 12942 1928 12995 1940
rect 12942 1894 12953 1928
rect 12987 1894 12995 1928
rect 12942 1856 12995 1894
rect 13170 1911 13178 1945
rect 13212 1911 13223 1945
rect 13170 1877 13223 1911
rect 13170 1843 13178 1877
rect 13212 1843 13223 1877
rect 13170 1831 13223 1843
rect 13323 2353 13379 2431
rect 13323 2319 13334 2353
rect 13368 2319 13379 2353
rect 13323 2285 13379 2319
rect 13323 2251 13334 2285
rect 13368 2251 13379 2285
rect 13323 2217 13379 2251
rect 13323 2183 13334 2217
rect 13368 2183 13379 2217
rect 13323 2149 13379 2183
rect 13323 2115 13334 2149
rect 13368 2115 13379 2149
rect 13323 2081 13379 2115
rect 13323 2047 13334 2081
rect 13368 2047 13379 2081
rect 13323 2013 13379 2047
rect 13323 1979 13334 2013
rect 13368 1979 13379 2013
rect 13323 1945 13379 1979
rect 13323 1911 13334 1945
rect 13368 1911 13379 1945
rect 13323 1877 13379 1911
rect 13323 1843 13334 1877
rect 13368 1843 13379 1877
rect 13323 1831 13379 1843
rect 13479 2353 13535 2431
rect 13479 2319 13490 2353
rect 13524 2319 13535 2353
rect 13479 2285 13535 2319
rect 13479 2251 13490 2285
rect 13524 2251 13535 2285
rect 13479 2217 13535 2251
rect 13479 2183 13490 2217
rect 13524 2183 13535 2217
rect 13479 2149 13535 2183
rect 13479 2115 13490 2149
rect 13524 2115 13535 2149
rect 13479 2081 13535 2115
rect 13479 2047 13490 2081
rect 13524 2047 13535 2081
rect 13479 2013 13535 2047
rect 13479 1979 13490 2013
rect 13524 1979 13535 2013
rect 13479 1945 13535 1979
rect 13479 1911 13490 1945
rect 13524 1911 13535 1945
rect 13479 1877 13535 1911
rect 13479 1843 13490 1877
rect 13524 1843 13535 1877
rect 13479 1831 13535 1843
rect 13635 2353 13691 2431
rect 13635 2319 13646 2353
rect 13680 2319 13691 2353
rect 13635 2285 13691 2319
rect 13635 2251 13646 2285
rect 13680 2251 13691 2285
rect 13635 2217 13691 2251
rect 13635 2183 13646 2217
rect 13680 2183 13691 2217
rect 13635 2149 13691 2183
rect 13635 2115 13646 2149
rect 13680 2115 13691 2149
rect 13635 2081 13691 2115
rect 13635 2047 13646 2081
rect 13680 2047 13691 2081
rect 13635 2013 13691 2047
rect 13635 1979 13646 2013
rect 13680 1979 13691 2013
rect 13635 1945 13691 1979
rect 13635 1911 13646 1945
rect 13680 1911 13691 1945
rect 13635 1877 13691 1911
rect 13635 1843 13646 1877
rect 13680 1843 13691 1877
rect 13635 1831 13691 1843
rect 13791 2353 13847 2431
rect 13791 2319 13802 2353
rect 13836 2319 13847 2353
rect 13791 2285 13847 2319
rect 13791 2251 13802 2285
rect 13836 2251 13847 2285
rect 13791 2217 13847 2251
rect 13791 2183 13802 2217
rect 13836 2183 13847 2217
rect 13791 2149 13847 2183
rect 13791 2115 13802 2149
rect 13836 2115 13847 2149
rect 13791 2081 13847 2115
rect 13791 2047 13802 2081
rect 13836 2047 13847 2081
rect 13791 2013 13847 2047
rect 13791 1979 13802 2013
rect 13836 1979 13847 2013
rect 13791 1945 13847 1979
rect 13791 1911 13802 1945
rect 13836 1911 13847 1945
rect 13791 1877 13847 1911
rect 13791 1843 13802 1877
rect 13836 1843 13847 1877
rect 13791 1831 13847 1843
rect 13947 2353 14003 2431
rect 13947 2319 13958 2353
rect 13992 2319 14003 2353
rect 13947 2285 14003 2319
rect 13947 2251 13958 2285
rect 13992 2251 14003 2285
rect 13947 2217 14003 2251
rect 13947 2183 13958 2217
rect 13992 2183 14003 2217
rect 13947 2149 14003 2183
rect 13947 2115 13958 2149
rect 13992 2115 14003 2149
rect 13947 2081 14003 2115
rect 13947 2047 13958 2081
rect 13992 2047 14003 2081
rect 13947 2013 14003 2047
rect 13947 1979 13958 2013
rect 13992 1979 14003 2013
rect 13947 1945 14003 1979
rect 13947 1911 13958 1945
rect 13992 1911 14003 1945
rect 13947 1877 14003 1911
rect 13947 1843 13958 1877
rect 13992 1843 14003 1877
rect 13947 1831 14003 1843
rect 14103 2353 14159 2431
rect 14103 2319 14114 2353
rect 14148 2319 14159 2353
rect 14103 2285 14159 2319
rect 14103 2251 14114 2285
rect 14148 2251 14159 2285
rect 14103 2217 14159 2251
rect 14103 2183 14114 2217
rect 14148 2183 14159 2217
rect 14103 2149 14159 2183
rect 14103 2115 14114 2149
rect 14148 2115 14159 2149
rect 14103 2081 14159 2115
rect 14103 2047 14114 2081
rect 14148 2047 14159 2081
rect 14103 2013 14159 2047
rect 14103 1979 14114 2013
rect 14148 1979 14159 2013
rect 14103 1945 14159 1979
rect 14103 1911 14114 1945
rect 14148 1911 14159 1945
rect 14103 1877 14159 1911
rect 14103 1843 14114 1877
rect 14148 1843 14159 1877
rect 14103 1831 14159 1843
rect 14259 2353 14315 2431
rect 14259 2319 14270 2353
rect 14304 2319 14315 2353
rect 14259 2285 14315 2319
rect 14259 2251 14270 2285
rect 14304 2251 14315 2285
rect 14259 2217 14315 2251
rect 14259 2183 14270 2217
rect 14304 2183 14315 2217
rect 14259 2149 14315 2183
rect 14259 2115 14270 2149
rect 14304 2115 14315 2149
rect 14259 2081 14315 2115
rect 14259 2047 14270 2081
rect 14304 2047 14315 2081
rect 14259 2013 14315 2047
rect 14259 1979 14270 2013
rect 14304 1979 14315 2013
rect 14259 1945 14315 1979
rect 14259 1911 14270 1945
rect 14304 1911 14315 1945
rect 14259 1877 14315 1911
rect 14259 1843 14270 1877
rect 14304 1843 14315 1877
rect 14259 1831 14315 1843
rect 14415 2353 14471 2431
rect 14415 2319 14426 2353
rect 14460 2319 14471 2353
rect 14415 2285 14471 2319
rect 14415 2251 14426 2285
rect 14460 2251 14471 2285
rect 14415 2217 14471 2251
rect 14415 2183 14426 2217
rect 14460 2183 14471 2217
rect 14415 2149 14471 2183
rect 14415 2115 14426 2149
rect 14460 2115 14471 2149
rect 14415 2081 14471 2115
rect 14415 2047 14426 2081
rect 14460 2047 14471 2081
rect 14415 2013 14471 2047
rect 14415 1979 14426 2013
rect 14460 1979 14471 2013
rect 14415 1945 14471 1979
rect 14415 1911 14426 1945
rect 14460 1911 14471 1945
rect 14415 1877 14471 1911
rect 14415 1843 14426 1877
rect 14460 1843 14471 1877
rect 14415 1831 14471 1843
rect 14571 2353 14627 2431
rect 14571 2319 14582 2353
rect 14616 2319 14627 2353
rect 14571 2285 14627 2319
rect 14571 2251 14582 2285
rect 14616 2251 14627 2285
rect 14571 2217 14627 2251
rect 14571 2183 14582 2217
rect 14616 2183 14627 2217
rect 14571 2149 14627 2183
rect 14571 2115 14582 2149
rect 14616 2115 14627 2149
rect 14571 2081 14627 2115
rect 14571 2047 14582 2081
rect 14616 2047 14627 2081
rect 14571 2013 14627 2047
rect 14571 1979 14582 2013
rect 14616 1979 14627 2013
rect 14571 1945 14627 1979
rect 14571 1911 14582 1945
rect 14616 1911 14627 1945
rect 14571 1877 14627 1911
rect 14571 1843 14582 1877
rect 14616 1843 14627 1877
rect 14571 1831 14627 1843
rect 14727 2353 14783 2431
rect 14727 2319 14738 2353
rect 14772 2319 14783 2353
rect 14727 2285 14783 2319
rect 14727 2251 14738 2285
rect 14772 2251 14783 2285
rect 14727 2217 14783 2251
rect 14727 2183 14738 2217
rect 14772 2183 14783 2217
rect 14727 2149 14783 2183
rect 14727 2115 14738 2149
rect 14772 2115 14783 2149
rect 14727 2081 14783 2115
rect 14727 2047 14738 2081
rect 14772 2047 14783 2081
rect 14727 2013 14783 2047
rect 14727 1979 14738 2013
rect 14772 1979 14783 2013
rect 14727 1945 14783 1979
rect 14727 1911 14738 1945
rect 14772 1911 14783 1945
rect 14727 1877 14783 1911
rect 14727 1843 14738 1877
rect 14772 1843 14783 1877
rect 14727 1831 14783 1843
rect 14883 2353 14939 2431
rect 14883 2319 14894 2353
rect 14928 2319 14939 2353
rect 14883 2285 14939 2319
rect 14883 2251 14894 2285
rect 14928 2251 14939 2285
rect 14883 2217 14939 2251
rect 14883 2183 14894 2217
rect 14928 2183 14939 2217
rect 14883 2149 14939 2183
rect 14883 2115 14894 2149
rect 14928 2115 14939 2149
rect 14883 2081 14939 2115
rect 14883 2047 14894 2081
rect 14928 2047 14939 2081
rect 14883 2013 14939 2047
rect 14883 1979 14894 2013
rect 14928 1979 14939 2013
rect 14883 1945 14939 1979
rect 14883 1911 14894 1945
rect 14928 1911 14939 1945
rect 14883 1877 14939 1911
rect 14883 1843 14894 1877
rect 14928 1843 14939 1877
rect 14883 1831 14939 1843
rect 15039 2353 15092 2431
rect 15039 2319 15050 2353
rect 15084 2319 15092 2353
rect 15039 2285 15092 2319
rect 15039 2251 15050 2285
rect 15084 2251 15092 2285
rect 15039 2217 15092 2251
rect 15039 2183 15050 2217
rect 15084 2183 15092 2217
rect 15039 2149 15092 2183
rect 15039 2115 15050 2149
rect 15084 2115 15092 2149
rect 15039 2081 15092 2115
rect 15039 2047 15050 2081
rect 15084 2047 15092 2081
rect 15039 2013 15092 2047
rect 15039 1979 15050 2013
rect 15084 1979 15092 2013
rect 15039 1945 15092 1979
rect 15039 1911 15050 1945
rect 15084 1911 15092 1945
rect 15039 1877 15092 1911
rect 15039 1843 15050 1877
rect 15084 1843 15092 1877
rect 15039 1831 15092 1843
<< mvndiffc >>
rect 11749 3520 11783 3554
rect 11749 3452 11783 3486
rect 11749 3384 11783 3418
rect 11749 3316 11783 3350
rect 11749 3248 11783 3282
rect 11749 3180 11783 3214
rect 11749 3112 11783 3146
rect 11749 3044 11783 3078
rect 11905 3520 11939 3554
rect 11905 3452 11939 3486
rect 11905 3384 11939 3418
rect 11905 3316 11939 3350
rect 11905 3248 11939 3282
rect 11905 3180 11939 3214
rect 11905 3112 11939 3146
rect 11905 3044 11939 3078
rect 12061 3520 12095 3554
rect 12061 3452 12095 3486
rect 12061 3384 12095 3418
rect 12061 3316 12095 3350
rect 12061 3248 12095 3282
rect 12061 3180 12095 3214
rect 12061 3112 12095 3146
rect 12061 3044 12095 3078
rect 12217 3520 12251 3554
rect 12217 3452 12251 3486
rect 12217 3384 12251 3418
rect 12217 3316 12251 3350
rect 12217 3248 12251 3282
rect 12217 3180 12251 3214
rect 12217 3112 12251 3146
rect 12217 3044 12251 3078
rect 12373 3520 12407 3554
rect 12373 3452 12407 3486
rect 12373 3384 12407 3418
rect 12373 3316 12407 3350
rect 12373 3248 12407 3282
rect 12373 3180 12407 3214
rect 12373 3112 12407 3146
rect 12373 3044 12407 3078
rect 12529 3520 12563 3554
rect 12529 3452 12563 3486
rect 12529 3384 12563 3418
rect 12529 3316 12563 3350
rect 12529 3248 12563 3282
rect 12529 3180 12563 3214
rect 12529 3112 12563 3146
rect 12529 3044 12563 3078
rect 12685 3520 12719 3554
rect 12685 3452 12719 3486
rect 12685 3384 12719 3418
rect 12685 3316 12719 3350
rect 12685 3248 12719 3282
rect 12685 3180 12719 3214
rect 12685 3112 12719 3146
rect 12685 3044 12719 3078
rect 12841 3520 12875 3554
rect 12841 3452 12875 3486
rect 12841 3384 12875 3418
rect 12841 3316 12875 3350
rect 12841 3248 12875 3282
rect 12841 3180 12875 3214
rect 12841 3112 12875 3146
rect 12841 3044 12875 3078
rect 12997 3520 13031 3554
rect 12997 3452 13031 3486
rect 12997 3384 13031 3418
rect 12997 3316 13031 3350
rect 12997 3248 13031 3282
rect 12997 3180 13031 3214
rect 12997 3112 13031 3146
rect 12997 3044 13031 3078
rect 13153 3520 13187 3554
rect 13153 3452 13187 3486
rect 13153 3384 13187 3418
rect 13153 3316 13187 3350
rect 13153 3248 13187 3282
rect 13153 3180 13187 3214
rect 13153 3112 13187 3146
rect 13153 3044 13187 3078
rect 13309 3520 13343 3554
rect 13309 3452 13343 3486
rect 13309 3384 13343 3418
rect 13309 3316 13343 3350
rect 13309 3248 13343 3282
rect 13309 3180 13343 3214
rect 13309 3112 13343 3146
rect 13309 3044 13343 3078
rect 13465 3520 13499 3554
rect 13465 3452 13499 3486
rect 13465 3384 13499 3418
rect 13465 3316 13499 3350
rect 13465 3248 13499 3282
rect 13465 3180 13499 3214
rect 13465 3112 13499 3146
rect 13465 3044 13499 3078
rect 13621 3520 13655 3554
rect 13621 3452 13655 3486
rect 13621 3384 13655 3418
rect 13621 3316 13655 3350
rect 13621 3248 13655 3282
rect 13621 3180 13655 3214
rect 13621 3112 13655 3146
rect 13621 3044 13655 3078
rect 13742 3520 13776 3554
rect 13742 3452 13776 3486
rect 13742 3384 13776 3418
rect 13742 3316 13776 3350
rect 13742 3248 13776 3282
rect 13742 3180 13776 3214
rect 13742 3112 13776 3146
rect 13742 3044 13776 3078
rect 13918 3520 13952 3554
rect 13918 3452 13952 3486
rect 13918 3384 13952 3418
rect 13918 3316 13952 3350
rect 13918 3248 13952 3282
rect 13918 3180 13952 3214
rect 13918 3112 13952 3146
rect 13918 3044 13952 3078
rect 14042 3520 14076 3554
rect 14042 3452 14076 3486
rect 14042 3384 14076 3418
rect 14042 3316 14076 3350
rect 14042 3248 14076 3282
rect 14042 3180 14076 3214
rect 14042 3112 14076 3146
rect 14042 3044 14076 3078
rect 14218 3520 14252 3554
rect 14218 3452 14252 3486
rect 14218 3384 14252 3418
rect 14218 3316 14252 3350
rect 14218 3248 14252 3282
rect 14218 3180 14252 3214
rect 14218 3112 14252 3146
rect 14218 3044 14252 3078
rect 14374 3520 14408 3554
rect 14374 3452 14408 3486
rect 14374 3384 14408 3418
rect 14374 3316 14408 3350
rect 14374 3248 14408 3282
rect 14374 3180 14408 3214
rect 14374 3112 14408 3146
rect 14374 3044 14408 3078
rect 14530 3520 14564 3554
rect 14530 3452 14564 3486
rect 14530 3384 14564 3418
rect 14530 3316 14564 3350
rect 14530 3248 14564 3282
rect 14530 3180 14564 3214
rect 14530 3112 14564 3146
rect 14530 3044 14564 3078
rect 12423 2446 12457 2480
rect 12679 2446 12713 2480
rect 12935 2446 12969 2480
<< mvpdiffc >>
rect 35591 15083 35625 15117
rect 35659 15083 35693 15117
rect 35727 15083 35761 15117
rect 35795 15083 35829 15117
rect 35863 15083 35897 15117
rect 35931 15083 35965 15117
rect 35999 15083 36033 15117
rect 36067 15083 36101 15117
rect 36135 15083 36169 15117
rect 36203 15083 36237 15117
rect 36271 15083 36305 15117
rect 36339 15083 36373 15117
rect 36407 15083 36441 15117
rect 36475 15083 36509 15117
rect 36543 15083 36577 15117
rect 36611 15083 36645 15117
rect 36679 15083 36713 15117
rect 36747 15083 36781 15117
rect 36815 15083 36849 15117
rect 36883 15083 36917 15117
rect 36951 15083 36985 15117
rect 37019 15083 37053 15117
rect 37087 15083 37121 15117
rect 37155 15083 37189 15117
rect 37223 15083 37257 15117
rect 37291 15083 37325 15117
rect 37359 15083 37393 15117
rect 37427 15083 37461 15117
rect 37495 15083 37529 15117
rect 35591 14927 35625 14961
rect 35659 14927 35693 14961
rect 35727 14927 35761 14961
rect 35795 14927 35829 14961
rect 35863 14927 35897 14961
rect 35931 14927 35965 14961
rect 35999 14927 36033 14961
rect 36067 14927 36101 14961
rect 36135 14927 36169 14961
rect 36203 14927 36237 14961
rect 36271 14927 36305 14961
rect 36339 14927 36373 14961
rect 36407 14927 36441 14961
rect 36475 14927 36509 14961
rect 36543 14927 36577 14961
rect 36611 14927 36645 14961
rect 36679 14927 36713 14961
rect 36747 14927 36781 14961
rect 36815 14927 36849 14961
rect 36883 14927 36917 14961
rect 36951 14927 36985 14961
rect 37019 14927 37053 14961
rect 37087 14927 37121 14961
rect 37155 14927 37189 14961
rect 37223 14927 37257 14961
rect 37291 14927 37325 14961
rect 37359 14927 37393 14961
rect 37427 14927 37461 14961
rect 37495 14927 37529 14961
rect 35591 14771 35625 14805
rect 35659 14771 35693 14805
rect 35727 14771 35761 14805
rect 35795 14771 35829 14805
rect 35863 14771 35897 14805
rect 35931 14771 35965 14805
rect 35999 14771 36033 14805
rect 36067 14771 36101 14805
rect 36135 14771 36169 14805
rect 36203 14771 36237 14805
rect 36271 14771 36305 14805
rect 36339 14771 36373 14805
rect 36407 14771 36441 14805
rect 36475 14771 36509 14805
rect 36543 14771 36577 14805
rect 36611 14771 36645 14805
rect 36679 14771 36713 14805
rect 36747 14771 36781 14805
rect 36815 14771 36849 14805
rect 36883 14771 36917 14805
rect 36951 14771 36985 14805
rect 37019 14771 37053 14805
rect 37087 14771 37121 14805
rect 37155 14771 37189 14805
rect 37223 14771 37257 14805
rect 37291 14771 37325 14805
rect 37359 14771 37393 14805
rect 37427 14771 37461 14805
rect 37495 14771 37529 14805
rect 35591 14615 35625 14649
rect 35659 14615 35693 14649
rect 35727 14615 35761 14649
rect 35795 14615 35829 14649
rect 35863 14615 35897 14649
rect 35931 14615 35965 14649
rect 35999 14615 36033 14649
rect 36067 14615 36101 14649
rect 36135 14615 36169 14649
rect 36203 14615 36237 14649
rect 36271 14615 36305 14649
rect 36339 14615 36373 14649
rect 36407 14615 36441 14649
rect 36475 14615 36509 14649
rect 36543 14615 36577 14649
rect 36611 14615 36645 14649
rect 36679 14615 36713 14649
rect 36747 14615 36781 14649
rect 36815 14615 36849 14649
rect 36883 14615 36917 14649
rect 36951 14615 36985 14649
rect 37019 14615 37053 14649
rect 37087 14615 37121 14649
rect 37155 14615 37189 14649
rect 37223 14615 37257 14649
rect 37291 14615 37325 14649
rect 37359 14615 37393 14649
rect 37427 14615 37461 14649
rect 37495 14615 37529 14649
rect 35591 14459 35625 14493
rect 35659 14459 35693 14493
rect 35727 14459 35761 14493
rect 35795 14459 35829 14493
rect 35863 14459 35897 14493
rect 35931 14459 35965 14493
rect 35999 14459 36033 14493
rect 36067 14459 36101 14493
rect 36135 14459 36169 14493
rect 36203 14459 36237 14493
rect 36271 14459 36305 14493
rect 36339 14459 36373 14493
rect 36407 14459 36441 14493
rect 36475 14459 36509 14493
rect 36543 14459 36577 14493
rect 36611 14459 36645 14493
rect 36679 14459 36713 14493
rect 36747 14459 36781 14493
rect 36815 14459 36849 14493
rect 36883 14459 36917 14493
rect 36951 14459 36985 14493
rect 37019 14459 37053 14493
rect 37087 14459 37121 14493
rect 37155 14459 37189 14493
rect 37223 14459 37257 14493
rect 37291 14459 37325 14493
rect 37359 14459 37393 14493
rect 37427 14459 37461 14493
rect 37495 14459 37529 14493
rect 35591 14303 35625 14337
rect 35659 14303 35693 14337
rect 35727 14303 35761 14337
rect 35795 14303 35829 14337
rect 35863 14303 35897 14337
rect 35931 14303 35965 14337
rect 35999 14303 36033 14337
rect 36067 14303 36101 14337
rect 36135 14303 36169 14337
rect 36203 14303 36237 14337
rect 36271 14303 36305 14337
rect 36339 14303 36373 14337
rect 36407 14303 36441 14337
rect 36475 14303 36509 14337
rect 36543 14303 36577 14337
rect 36611 14303 36645 14337
rect 36679 14303 36713 14337
rect 36747 14303 36781 14337
rect 36815 14303 36849 14337
rect 36883 14303 36917 14337
rect 36951 14303 36985 14337
rect 37019 14303 37053 14337
rect 37087 14303 37121 14337
rect 37155 14303 37189 14337
rect 37223 14303 37257 14337
rect 37291 14303 37325 14337
rect 37359 14303 37393 14337
rect 37427 14303 37461 14337
rect 37495 14303 37529 14337
rect 35591 14147 35625 14181
rect 35659 14147 35693 14181
rect 35727 14147 35761 14181
rect 35795 14147 35829 14181
rect 35863 14147 35897 14181
rect 35931 14147 35965 14181
rect 35999 14147 36033 14181
rect 36067 14147 36101 14181
rect 36135 14147 36169 14181
rect 36203 14147 36237 14181
rect 36271 14147 36305 14181
rect 36339 14147 36373 14181
rect 36407 14147 36441 14181
rect 36475 14147 36509 14181
rect 36543 14147 36577 14181
rect 36611 14147 36645 14181
rect 36679 14147 36713 14181
rect 36747 14147 36781 14181
rect 36815 14147 36849 14181
rect 36883 14147 36917 14181
rect 36951 14147 36985 14181
rect 37019 14147 37053 14181
rect 37087 14147 37121 14181
rect 37155 14147 37189 14181
rect 37223 14147 37257 14181
rect 37291 14147 37325 14181
rect 37359 14147 37393 14181
rect 37427 14147 37461 14181
rect 37495 14147 37529 14181
rect 35591 13991 35625 14025
rect 35659 13991 35693 14025
rect 35727 13991 35761 14025
rect 35795 13991 35829 14025
rect 35863 13991 35897 14025
rect 35931 13991 35965 14025
rect 35999 13991 36033 14025
rect 36067 13991 36101 14025
rect 36135 13991 36169 14025
rect 36203 13991 36237 14025
rect 36271 13991 36305 14025
rect 36339 13991 36373 14025
rect 36407 13991 36441 14025
rect 36475 13991 36509 14025
rect 36543 13991 36577 14025
rect 36611 13991 36645 14025
rect 36679 13991 36713 14025
rect 36747 13991 36781 14025
rect 36815 13991 36849 14025
rect 36883 13991 36917 14025
rect 36951 13991 36985 14025
rect 37019 13991 37053 14025
rect 37087 13991 37121 14025
rect 37155 13991 37189 14025
rect 37223 13991 37257 14025
rect 37291 13991 37325 14025
rect 37359 13991 37393 14025
rect 37427 13991 37461 14025
rect 37495 13991 37529 14025
rect 35591 13835 35625 13869
rect 35659 13835 35693 13869
rect 35727 13835 35761 13869
rect 35795 13835 35829 13869
rect 35863 13835 35897 13869
rect 35931 13835 35965 13869
rect 35999 13835 36033 13869
rect 36067 13835 36101 13869
rect 36135 13835 36169 13869
rect 36203 13835 36237 13869
rect 36271 13835 36305 13869
rect 36339 13835 36373 13869
rect 36407 13835 36441 13869
rect 36475 13835 36509 13869
rect 36543 13835 36577 13869
rect 36611 13835 36645 13869
rect 36679 13835 36713 13869
rect 36747 13835 36781 13869
rect 36815 13835 36849 13869
rect 36883 13835 36917 13869
rect 36951 13835 36985 13869
rect 37019 13835 37053 13869
rect 37087 13835 37121 13869
rect 37155 13835 37189 13869
rect 37223 13835 37257 13869
rect 37291 13835 37325 13869
rect 37359 13835 37393 13869
rect 37427 13835 37461 13869
rect 37495 13835 37529 13869
rect 35591 13679 35625 13713
rect 35659 13679 35693 13713
rect 35727 13679 35761 13713
rect 35795 13679 35829 13713
rect 35863 13679 35897 13713
rect 35931 13679 35965 13713
rect 35999 13679 36033 13713
rect 36067 13679 36101 13713
rect 36135 13679 36169 13713
rect 36203 13679 36237 13713
rect 36271 13679 36305 13713
rect 36339 13679 36373 13713
rect 36407 13679 36441 13713
rect 36475 13679 36509 13713
rect 36543 13679 36577 13713
rect 36611 13679 36645 13713
rect 36679 13679 36713 13713
rect 36747 13679 36781 13713
rect 36815 13679 36849 13713
rect 36883 13679 36917 13713
rect 36951 13679 36985 13713
rect 37019 13679 37053 13713
rect 37087 13679 37121 13713
rect 37155 13679 37189 13713
rect 37223 13679 37257 13713
rect 37291 13679 37325 13713
rect 37359 13679 37393 13713
rect 37427 13679 37461 13713
rect 37495 13679 37529 13713
rect 35591 13523 35625 13557
rect 35659 13523 35693 13557
rect 35727 13523 35761 13557
rect 35795 13523 35829 13557
rect 35863 13523 35897 13557
rect 35931 13523 35965 13557
rect 35999 13523 36033 13557
rect 36067 13523 36101 13557
rect 36135 13523 36169 13557
rect 36203 13523 36237 13557
rect 36271 13523 36305 13557
rect 36339 13523 36373 13557
rect 36407 13523 36441 13557
rect 36475 13523 36509 13557
rect 36543 13523 36577 13557
rect 36611 13523 36645 13557
rect 36679 13523 36713 13557
rect 36747 13523 36781 13557
rect 36815 13523 36849 13557
rect 36883 13523 36917 13557
rect 36951 13523 36985 13557
rect 37019 13523 37053 13557
rect 37087 13523 37121 13557
rect 37155 13523 37189 13557
rect 37223 13523 37257 13557
rect 37291 13523 37325 13557
rect 37359 13523 37393 13557
rect 37427 13523 37461 13557
rect 37495 13523 37529 13557
rect 35591 13367 35625 13401
rect 35659 13367 35693 13401
rect 35727 13367 35761 13401
rect 35795 13367 35829 13401
rect 35863 13367 35897 13401
rect 35931 13367 35965 13401
rect 35999 13367 36033 13401
rect 36067 13367 36101 13401
rect 36135 13367 36169 13401
rect 36203 13367 36237 13401
rect 36271 13367 36305 13401
rect 36339 13367 36373 13401
rect 36407 13367 36441 13401
rect 36475 13367 36509 13401
rect 36543 13367 36577 13401
rect 36611 13367 36645 13401
rect 36679 13367 36713 13401
rect 36747 13367 36781 13401
rect 36815 13367 36849 13401
rect 36883 13367 36917 13401
rect 36951 13367 36985 13401
rect 37019 13367 37053 13401
rect 37087 13367 37121 13401
rect 37155 13367 37189 13401
rect 37223 13367 37257 13401
rect 37291 13367 37325 13401
rect 37359 13367 37393 13401
rect 37427 13367 37461 13401
rect 37495 13367 37529 13401
rect 35591 13211 35625 13245
rect 35659 13211 35693 13245
rect 35727 13211 35761 13245
rect 35795 13211 35829 13245
rect 35863 13211 35897 13245
rect 35931 13211 35965 13245
rect 35999 13211 36033 13245
rect 36067 13211 36101 13245
rect 36135 13211 36169 13245
rect 36203 13211 36237 13245
rect 36271 13211 36305 13245
rect 36339 13211 36373 13245
rect 36407 13211 36441 13245
rect 36475 13211 36509 13245
rect 36543 13211 36577 13245
rect 36611 13211 36645 13245
rect 36679 13211 36713 13245
rect 36747 13211 36781 13245
rect 36815 13211 36849 13245
rect 36883 13211 36917 13245
rect 36951 13211 36985 13245
rect 37019 13211 37053 13245
rect 37087 13211 37121 13245
rect 37155 13211 37189 13245
rect 37223 13211 37257 13245
rect 37291 13211 37325 13245
rect 37359 13211 37393 13245
rect 37427 13211 37461 13245
rect 37495 13211 37529 13245
rect 13178 2319 13212 2353
rect 13178 2251 13212 2285
rect 12423 2149 12457 2183
rect 12679 2149 12713 2183
rect 12935 2149 12969 2183
rect 13178 2183 13212 2217
rect 13178 2115 13212 2149
rect 13178 2047 13212 2081
rect 13178 1979 13212 2013
rect 12041 1894 12075 1928
rect 12497 1894 12531 1928
rect 12953 1894 12987 1928
rect 13178 1911 13212 1945
rect 13178 1843 13212 1877
rect 13334 2319 13368 2353
rect 13334 2251 13368 2285
rect 13334 2183 13368 2217
rect 13334 2115 13368 2149
rect 13334 2047 13368 2081
rect 13334 1979 13368 2013
rect 13334 1911 13368 1945
rect 13334 1843 13368 1877
rect 13490 2319 13524 2353
rect 13490 2251 13524 2285
rect 13490 2183 13524 2217
rect 13490 2115 13524 2149
rect 13490 2047 13524 2081
rect 13490 1979 13524 2013
rect 13490 1911 13524 1945
rect 13490 1843 13524 1877
rect 13646 2319 13680 2353
rect 13646 2251 13680 2285
rect 13646 2183 13680 2217
rect 13646 2115 13680 2149
rect 13646 2047 13680 2081
rect 13646 1979 13680 2013
rect 13646 1911 13680 1945
rect 13646 1843 13680 1877
rect 13802 2319 13836 2353
rect 13802 2251 13836 2285
rect 13802 2183 13836 2217
rect 13802 2115 13836 2149
rect 13802 2047 13836 2081
rect 13802 1979 13836 2013
rect 13802 1911 13836 1945
rect 13802 1843 13836 1877
rect 13958 2319 13992 2353
rect 13958 2251 13992 2285
rect 13958 2183 13992 2217
rect 13958 2115 13992 2149
rect 13958 2047 13992 2081
rect 13958 1979 13992 2013
rect 13958 1911 13992 1945
rect 13958 1843 13992 1877
rect 14114 2319 14148 2353
rect 14114 2251 14148 2285
rect 14114 2183 14148 2217
rect 14114 2115 14148 2149
rect 14114 2047 14148 2081
rect 14114 1979 14148 2013
rect 14114 1911 14148 1945
rect 14114 1843 14148 1877
rect 14270 2319 14304 2353
rect 14270 2251 14304 2285
rect 14270 2183 14304 2217
rect 14270 2115 14304 2149
rect 14270 2047 14304 2081
rect 14270 1979 14304 2013
rect 14270 1911 14304 1945
rect 14270 1843 14304 1877
rect 14426 2319 14460 2353
rect 14426 2251 14460 2285
rect 14426 2183 14460 2217
rect 14426 2115 14460 2149
rect 14426 2047 14460 2081
rect 14426 1979 14460 2013
rect 14426 1911 14460 1945
rect 14426 1843 14460 1877
rect 14582 2319 14616 2353
rect 14582 2251 14616 2285
rect 14582 2183 14616 2217
rect 14582 2115 14616 2149
rect 14582 2047 14616 2081
rect 14582 1979 14616 2013
rect 14582 1911 14616 1945
rect 14582 1843 14616 1877
rect 14738 2319 14772 2353
rect 14738 2251 14772 2285
rect 14738 2183 14772 2217
rect 14738 2115 14772 2149
rect 14738 2047 14772 2081
rect 14738 1979 14772 2013
rect 14738 1911 14772 1945
rect 14738 1843 14772 1877
rect 14894 2319 14928 2353
rect 14894 2251 14928 2285
rect 14894 2183 14928 2217
rect 14894 2115 14928 2149
rect 14894 2047 14928 2081
rect 14894 1979 14928 2013
rect 14894 1911 14928 1945
rect 14894 1843 14928 1877
rect 15050 2319 15084 2353
rect 15050 2251 15084 2285
rect 15050 2183 15084 2217
rect 15050 2115 15084 2149
rect 15050 2047 15084 2081
rect 15050 1979 15084 2013
rect 15050 1911 15084 1945
rect 15050 1843 15084 1877
<< psubdiff >>
rect 20576 1657 20578 1691
rect 20612 1657 20647 1691
rect 20681 1657 20716 1691
rect 20750 1657 20785 1691
rect 20819 1657 20854 1691
rect 20888 1657 20923 1691
rect 20957 1657 20992 1691
rect 21026 1657 21061 1691
rect 21095 1657 21130 1691
rect 21164 1657 21199 1691
rect 21233 1657 21268 1691
rect 21302 1657 21337 1691
rect 21371 1657 21406 1691
rect 21440 1657 21475 1691
rect 21509 1657 21543 1691
rect 21577 1657 21611 1691
rect 21645 1657 21679 1691
rect 21713 1657 21747 1691
rect 21781 1657 21815 1691
rect 21849 1657 21883 1691
rect 21917 1657 21951 1691
rect 21985 1657 22019 1691
rect 22053 1657 22087 1691
rect 22121 1657 22155 1691
rect 22189 1657 22223 1691
rect 22257 1657 22291 1691
rect 22325 1657 22359 1691
rect 22393 1657 22427 1691
rect 22461 1657 22495 1691
rect 22529 1657 22563 1691
rect 22597 1657 22631 1691
rect 22665 1657 22699 1691
rect 22733 1657 22767 1691
rect 22801 1657 22835 1691
rect 22869 1657 22903 1691
rect 22937 1657 22971 1691
rect 23005 1657 23039 1691
rect 23073 1657 23107 1691
rect 23141 1657 23175 1691
rect 23209 1657 23243 1691
rect 23277 1657 23311 1691
rect 23345 1657 23379 1691
rect 23413 1657 23447 1691
rect 23481 1657 23515 1691
rect 23549 1657 23583 1691
rect 23617 1657 23641 1691
<< mvpsubdiff >>
rect 11721 3640 11745 3674
rect 11779 3640 11815 3674
rect 11849 3640 11885 3674
rect 11919 3640 11955 3674
rect 11989 3640 12025 3674
rect 12059 3640 12095 3674
rect 12129 3640 12165 3674
rect 12199 3640 12235 3674
rect 12269 3640 12305 3674
rect 12339 3640 12375 3674
rect 12409 3640 12445 3674
rect 12479 3640 12515 3674
rect 12549 3640 12585 3674
rect 12619 3640 12655 3674
rect 12689 3640 12725 3674
rect 12759 3640 12795 3674
rect 12829 3640 12864 3674
rect 12898 3640 12933 3674
rect 12967 3640 13002 3674
rect 13036 3640 13071 3674
rect 13105 3640 13140 3674
rect 13174 3640 13209 3674
rect 13243 3640 13278 3674
rect 13312 3640 13347 3674
rect 13381 3640 13416 3674
rect 13450 3640 13485 3674
rect 13519 3640 13554 3674
rect 13588 3640 13623 3674
rect 13657 3640 13692 3674
rect 13726 3640 13761 3674
rect 13795 3640 13830 3674
rect 13864 3640 13899 3674
rect 13933 3640 13968 3674
rect 14002 3640 14037 3674
rect 14071 3640 14106 3674
rect 14140 3640 14175 3674
rect 14209 3640 14244 3674
rect 14278 3640 14313 3674
rect 14347 3640 14382 3674
rect 14416 3640 14451 3674
rect 14485 3640 14520 3674
rect 14554 3640 14589 3674
rect 14623 3640 14647 3674
rect 12520 2566 12544 2600
rect 12578 2566 12614 2600
rect 12648 2566 12684 2600
rect 12718 2566 12753 2600
rect 12787 2566 12822 2600
rect 12856 2566 12880 2600
rect 18139 1657 18163 1691
rect 18197 1657 18232 1691
rect 18266 1657 18301 1691
rect 18335 1657 18370 1691
rect 18404 1657 18439 1691
rect 18473 1657 18508 1691
rect 18542 1657 18577 1691
rect 18611 1657 18646 1691
rect 18680 1657 18715 1691
rect 18749 1657 18784 1691
rect 18818 1657 18853 1691
rect 18887 1657 18922 1691
rect 18956 1657 18991 1691
rect 19025 1657 19060 1691
rect 19094 1657 19129 1691
rect 19163 1657 19198 1691
rect 19232 1657 19267 1691
rect 19301 1657 19336 1691
rect 19370 1657 19405 1691
rect 19439 1657 19474 1691
rect 19508 1657 19543 1691
rect 19577 1657 19612 1691
rect 19646 1657 19681 1691
rect 19715 1657 19750 1691
rect 19784 1657 19819 1691
rect 19853 1657 19888 1691
rect 19922 1657 19957 1691
rect 19991 1657 20026 1691
rect 20060 1657 20095 1691
rect 20129 1657 20164 1691
rect 20198 1657 20233 1691
rect 20267 1657 20302 1691
rect 20336 1657 20371 1691
rect 20405 1657 20440 1691
rect 20474 1657 20509 1691
rect 20543 1657 20576 1691
<< mvnsubdiff >>
rect 12063 1723 12087 1757
rect 12121 1723 12156 1757
rect 12190 1723 12225 1757
rect 12259 1723 12294 1757
rect 12328 1723 12363 1757
rect 12397 1723 12432 1757
rect 12466 1723 12501 1757
rect 12535 1723 12570 1757
rect 12604 1723 12639 1757
rect 12673 1723 12708 1757
rect 12742 1723 12777 1757
rect 12811 1723 12846 1757
rect 12880 1723 12915 1757
rect 12949 1723 12984 1757
rect 13018 1723 13053 1757
rect 13087 1723 13122 1757
rect 13156 1723 13191 1757
rect 13225 1723 13260 1757
rect 13294 1723 13329 1757
rect 13363 1723 13398 1757
rect 13432 1723 13467 1757
rect 13501 1723 13536 1757
rect 13570 1723 13605 1757
rect 13639 1723 13674 1757
rect 13708 1723 13743 1757
rect 13777 1723 13812 1757
rect 13846 1723 13881 1757
rect 13915 1723 13950 1757
rect 13984 1723 14019 1757
rect 14053 1723 14088 1757
rect 14122 1723 14157 1757
rect 14191 1723 14226 1757
rect 14260 1723 14295 1757
rect 14329 1723 14364 1757
rect 14398 1723 14433 1757
rect 14467 1723 14502 1757
rect 14536 1723 14571 1757
rect 14605 1723 14640 1757
rect 14674 1723 14709 1757
rect 14743 1723 14778 1757
rect 14812 1723 14847 1757
rect 14881 1723 14916 1757
rect 14950 1723 14985 1757
rect 15019 1723 15054 1757
rect 15088 1723 15123 1757
rect 15157 1723 15192 1757
rect 15226 1723 15261 1757
rect 15295 1723 15329 1757
rect 15363 1723 15397 1757
rect 15431 1723 15465 1757
rect 15499 1723 15533 1757
rect 15567 1723 15601 1757
rect 15635 1723 15669 1757
rect 15703 1723 15737 1757
rect 15771 1723 15795 1757
<< psubdiffcont >>
rect 20578 1657 20612 1691
rect 20647 1657 20681 1691
rect 20716 1657 20750 1691
rect 20785 1657 20819 1691
rect 20854 1657 20888 1691
rect 20923 1657 20957 1691
rect 20992 1657 21026 1691
rect 21061 1657 21095 1691
rect 21130 1657 21164 1691
rect 21199 1657 21233 1691
rect 21268 1657 21302 1691
rect 21337 1657 21371 1691
rect 21406 1657 21440 1691
rect 21475 1657 21509 1691
rect 21543 1657 21577 1691
rect 21611 1657 21645 1691
rect 21679 1657 21713 1691
rect 21747 1657 21781 1691
rect 21815 1657 21849 1691
rect 21883 1657 21917 1691
rect 21951 1657 21985 1691
rect 22019 1657 22053 1691
rect 22087 1657 22121 1691
rect 22155 1657 22189 1691
rect 22223 1657 22257 1691
rect 22291 1657 22325 1691
rect 22359 1657 22393 1691
rect 22427 1657 22461 1691
rect 22495 1657 22529 1691
rect 22563 1657 22597 1691
rect 22631 1657 22665 1691
rect 22699 1657 22733 1691
rect 22767 1657 22801 1691
rect 22835 1657 22869 1691
rect 22903 1657 22937 1691
rect 22971 1657 23005 1691
rect 23039 1657 23073 1691
rect 23107 1657 23141 1691
rect 23175 1657 23209 1691
rect 23243 1657 23277 1691
rect 23311 1657 23345 1691
rect 23379 1657 23413 1691
rect 23447 1657 23481 1691
rect 23515 1657 23549 1691
rect 23583 1657 23617 1691
<< mvpsubdiffcont >>
rect 11745 3640 11779 3674
rect 11815 3640 11849 3674
rect 11885 3640 11919 3674
rect 11955 3640 11989 3674
rect 12025 3640 12059 3674
rect 12095 3640 12129 3674
rect 12165 3640 12199 3674
rect 12235 3640 12269 3674
rect 12305 3640 12339 3674
rect 12375 3640 12409 3674
rect 12445 3640 12479 3674
rect 12515 3640 12549 3674
rect 12585 3640 12619 3674
rect 12655 3640 12689 3674
rect 12725 3640 12759 3674
rect 12795 3640 12829 3674
rect 12864 3640 12898 3674
rect 12933 3640 12967 3674
rect 13002 3640 13036 3674
rect 13071 3640 13105 3674
rect 13140 3640 13174 3674
rect 13209 3640 13243 3674
rect 13278 3640 13312 3674
rect 13347 3640 13381 3674
rect 13416 3640 13450 3674
rect 13485 3640 13519 3674
rect 13554 3640 13588 3674
rect 13623 3640 13657 3674
rect 13692 3640 13726 3674
rect 13761 3640 13795 3674
rect 13830 3640 13864 3674
rect 13899 3640 13933 3674
rect 13968 3640 14002 3674
rect 14037 3640 14071 3674
rect 14106 3640 14140 3674
rect 14175 3640 14209 3674
rect 14244 3640 14278 3674
rect 14313 3640 14347 3674
rect 14382 3640 14416 3674
rect 14451 3640 14485 3674
rect 14520 3640 14554 3674
rect 14589 3640 14623 3674
rect 12544 2566 12578 2600
rect 12614 2566 12648 2600
rect 12684 2566 12718 2600
rect 12753 2566 12787 2600
rect 12822 2566 12856 2600
rect 18163 1657 18197 1691
rect 18232 1657 18266 1691
rect 18301 1657 18335 1691
rect 18370 1657 18404 1691
rect 18439 1657 18473 1691
rect 18508 1657 18542 1691
rect 18577 1657 18611 1691
rect 18646 1657 18680 1691
rect 18715 1657 18749 1691
rect 18784 1657 18818 1691
rect 18853 1657 18887 1691
rect 18922 1657 18956 1691
rect 18991 1657 19025 1691
rect 19060 1657 19094 1691
rect 19129 1657 19163 1691
rect 19198 1657 19232 1691
rect 19267 1657 19301 1691
rect 19336 1657 19370 1691
rect 19405 1657 19439 1691
rect 19474 1657 19508 1691
rect 19543 1657 19577 1691
rect 19612 1657 19646 1691
rect 19681 1657 19715 1691
rect 19750 1657 19784 1691
rect 19819 1657 19853 1691
rect 19888 1657 19922 1691
rect 19957 1657 19991 1691
rect 20026 1657 20060 1691
rect 20095 1657 20129 1691
rect 20164 1657 20198 1691
rect 20233 1657 20267 1691
rect 20302 1657 20336 1691
rect 20371 1657 20405 1691
rect 20440 1657 20474 1691
rect 20509 1657 20543 1691
<< mvnsubdiffcont >>
rect 12087 1723 12121 1757
rect 12156 1723 12190 1757
rect 12225 1723 12259 1757
rect 12294 1723 12328 1757
rect 12363 1723 12397 1757
rect 12432 1723 12466 1757
rect 12501 1723 12535 1757
rect 12570 1723 12604 1757
rect 12639 1723 12673 1757
rect 12708 1723 12742 1757
rect 12777 1723 12811 1757
rect 12846 1723 12880 1757
rect 12915 1723 12949 1757
rect 12984 1723 13018 1757
rect 13053 1723 13087 1757
rect 13122 1723 13156 1757
rect 13191 1723 13225 1757
rect 13260 1723 13294 1757
rect 13329 1723 13363 1757
rect 13398 1723 13432 1757
rect 13467 1723 13501 1757
rect 13536 1723 13570 1757
rect 13605 1723 13639 1757
rect 13674 1723 13708 1757
rect 13743 1723 13777 1757
rect 13812 1723 13846 1757
rect 13881 1723 13915 1757
rect 13950 1723 13984 1757
rect 14019 1723 14053 1757
rect 14088 1723 14122 1757
rect 14157 1723 14191 1757
rect 14226 1723 14260 1757
rect 14295 1723 14329 1757
rect 14364 1723 14398 1757
rect 14433 1723 14467 1757
rect 14502 1723 14536 1757
rect 14571 1723 14605 1757
rect 14640 1723 14674 1757
rect 14709 1723 14743 1757
rect 14778 1723 14812 1757
rect 14847 1723 14881 1757
rect 14916 1723 14950 1757
rect 14985 1723 15019 1757
rect 15054 1723 15088 1757
rect 15123 1723 15157 1757
rect 15192 1723 15226 1757
rect 15261 1723 15295 1757
rect 15329 1723 15363 1757
rect 15397 1723 15431 1757
rect 15465 1723 15499 1757
rect 15533 1723 15567 1757
rect 15601 1723 15635 1757
rect 15669 1723 15703 1757
rect 15737 1723 15771 1757
<< poly >>
rect 35547 14972 35579 15072
rect 37579 15056 37677 15072
rect 37579 15022 37627 15056
rect 37661 15022 37677 15056
rect 37579 14986 37677 15022
rect 37579 14972 37627 14986
rect 37611 14952 37627 14972
rect 37661 14952 37677 14986
rect 37611 14916 37677 14952
rect 35547 14816 35579 14916
rect 37579 14882 37627 14916
rect 37661 14882 37677 14916
rect 37579 14846 37677 14882
rect 37579 14816 37627 14846
rect 37611 14812 37627 14816
rect 37661 14812 37677 14846
rect 37611 14776 37677 14812
rect 37611 14760 37627 14776
rect 35547 14660 35579 14760
rect 37579 14742 37627 14760
rect 37661 14742 37677 14776
rect 37579 14706 37677 14742
rect 37579 14672 37627 14706
rect 37661 14672 37677 14706
rect 37579 14660 37677 14672
rect 37611 14636 37677 14660
rect 37611 14604 37627 14636
rect 35547 14504 35579 14604
rect 37579 14602 37627 14604
rect 37661 14602 37677 14636
rect 37579 14566 37677 14602
rect 37579 14532 37627 14566
rect 37661 14532 37677 14566
rect 37579 14504 37677 14532
rect 37611 14496 37677 14504
rect 37611 14462 37627 14496
rect 37661 14462 37677 14496
rect 37611 14448 37677 14462
rect 35547 14348 35579 14448
rect 37579 14426 37677 14448
rect 37579 14392 37627 14426
rect 37661 14392 37677 14426
rect 37579 14356 37677 14392
rect 37579 14348 37627 14356
rect 37611 14322 37627 14348
rect 37661 14322 37677 14356
rect 37611 14292 37677 14322
rect 35547 14192 35579 14292
rect 37579 14286 37677 14292
rect 37579 14252 37627 14286
rect 37661 14252 37677 14286
rect 37579 14216 37677 14252
rect 37579 14192 37627 14216
rect 37611 14182 37627 14192
rect 37661 14182 37677 14216
rect 37611 14146 37677 14182
rect 37611 14136 37627 14146
rect 35547 14036 35579 14136
rect 37579 14112 37627 14136
rect 37661 14112 37677 14146
rect 37579 14076 37677 14112
rect 37579 14042 37627 14076
rect 37661 14042 37677 14076
rect 37579 14036 37677 14042
rect 37611 14006 37677 14036
rect 37611 13980 37627 14006
rect 35547 13880 35579 13980
rect 37579 13972 37627 13980
rect 37661 13972 37677 14006
rect 37579 13936 37677 13972
rect 37579 13902 37627 13936
rect 37661 13902 37677 13936
rect 37579 13880 37677 13902
rect 37611 13866 37677 13880
rect 37611 13832 37627 13866
rect 37661 13832 37677 13866
rect 37611 13824 37677 13832
rect 35547 13724 35579 13824
rect 37579 13796 37677 13824
rect 37579 13762 37627 13796
rect 37661 13762 37677 13796
rect 37579 13726 37677 13762
rect 37579 13724 37627 13726
rect 37611 13692 37627 13724
rect 37661 13692 37677 13726
rect 37611 13668 37677 13692
rect 35547 13568 35579 13668
rect 37579 13656 37677 13668
rect 37579 13622 37627 13656
rect 37661 13622 37677 13656
rect 37579 13586 37677 13622
rect 37579 13568 37627 13586
rect 37611 13552 37627 13568
rect 37661 13552 37677 13586
rect 37611 13516 37677 13552
rect 37611 13512 37627 13516
rect 35547 13412 35579 13512
rect 37579 13482 37627 13512
rect 37661 13482 37677 13516
rect 37579 13446 37677 13482
rect 37579 13412 37627 13446
rect 37661 13412 37677 13446
rect 37611 13376 37677 13412
rect 37611 13356 37627 13376
rect 35547 13256 35579 13356
rect 37579 13342 37627 13356
rect 37661 13342 37677 13376
rect 37579 13306 37677 13342
rect 37579 13272 37627 13306
rect 37661 13272 37677 13306
rect 37579 13256 37677 13272
rect 11794 3566 11894 3598
rect 11950 3566 12050 3598
rect 12106 3566 12206 3598
rect 12262 3566 12362 3598
rect 12418 3566 12518 3598
rect 12574 3566 12674 3598
rect 12730 3566 12830 3598
rect 12886 3566 12986 3598
rect 13042 3566 13142 3598
rect 13198 3566 13298 3598
rect 13354 3566 13454 3598
rect 13510 3566 13610 3598
rect 13787 3566 13907 3598
rect 14087 3566 14207 3598
rect 14263 3566 14363 3598
rect 14419 3566 14519 3598
rect 11794 2934 11894 2966
rect 11950 2934 12050 2966
rect 12106 2934 12206 2966
rect 12262 2934 12362 2966
rect 12418 2934 12518 2966
rect 12574 2934 12674 2966
rect 12730 2934 12830 2966
rect 12886 2934 12986 2966
rect 11794 2918 12361 2934
rect 11794 2884 11810 2918
rect 11844 2884 11882 2918
rect 11916 2884 11954 2918
rect 11988 2884 12026 2918
rect 12060 2884 12098 2918
rect 12132 2884 12169 2918
rect 12203 2884 12240 2918
rect 12274 2884 12311 2918
rect 12345 2884 12361 2918
rect 11794 2868 12361 2884
rect 12418 2918 12986 2934
rect 12418 2884 12434 2918
rect 12468 2884 12505 2918
rect 12539 2884 12576 2918
rect 12610 2884 12648 2918
rect 12682 2884 12720 2918
rect 12754 2884 12792 2918
rect 12826 2884 12864 2918
rect 12898 2884 12936 2918
rect 12970 2884 12986 2918
rect 12418 2868 12986 2884
rect 13042 2910 13142 2966
rect 13198 2934 13298 2966
rect 13354 2934 13454 2966
rect 13042 2876 13076 2910
rect 13110 2876 13142 2910
rect 13042 2842 13142 2876
rect 13199 2918 13454 2934
rect 13199 2884 13215 2918
rect 13249 2884 13309 2918
rect 13343 2884 13404 2918
rect 13438 2884 13454 2918
rect 13199 2868 13454 2884
rect 13510 2910 13610 2966
rect 13510 2876 13543 2910
rect 13577 2876 13610 2910
rect 13042 2808 13076 2842
rect 13110 2808 13142 2842
rect 13042 2792 13142 2808
rect 13510 2842 13610 2876
rect 13510 2808 13543 2842
rect 13577 2808 13610 2842
rect 13510 2792 13610 2808
rect 13787 2910 13907 2966
rect 13787 2876 13832 2910
rect 13866 2876 13907 2910
rect 13787 2842 13907 2876
rect 13787 2808 13832 2842
rect 13866 2808 13907 2842
rect 13787 2792 13907 2808
rect 14087 2901 14207 2966
rect 14087 2867 14122 2901
rect 14156 2867 14207 2901
rect 14087 2833 14207 2867
rect 14087 2799 14122 2833
rect 14156 2799 14207 2833
rect 14087 2783 14207 2799
rect 14263 2901 14363 2966
rect 14263 2867 14299 2901
rect 14333 2867 14363 2901
rect 14263 2833 14363 2867
rect 14263 2799 14299 2833
rect 14333 2799 14363 2833
rect 14263 2783 14363 2799
rect 14419 2901 14519 2966
rect 14419 2867 14453 2901
rect 14487 2867 14519 2901
rect 14419 2833 14519 2867
rect 14419 2799 14453 2833
rect 14487 2799 14519 2833
rect 14419 2783 14519 2799
rect 13223 2525 13479 2541
rect 12468 2492 12668 2524
rect 12724 2492 12924 2524
rect 13223 2491 13239 2525
rect 13273 2491 13334 2525
rect 13368 2491 13429 2525
rect 13463 2491 13479 2525
rect 13223 2475 13479 2491
rect 13223 2431 13323 2475
rect 13379 2431 13479 2475
rect 13535 2513 13791 2529
rect 13535 2479 13551 2513
rect 13585 2479 13646 2513
rect 13680 2479 13741 2513
rect 13775 2479 13791 2513
rect 13535 2463 13791 2479
rect 13535 2431 13635 2463
rect 13691 2431 13791 2463
rect 13847 2513 14415 2529
rect 13847 2479 13863 2513
rect 13897 2479 13935 2513
rect 13969 2479 14007 2513
rect 14041 2479 14079 2513
rect 14113 2479 14151 2513
rect 14185 2479 14223 2513
rect 14257 2479 14294 2513
rect 14328 2479 14365 2513
rect 14399 2479 14415 2513
rect 13847 2463 14415 2479
rect 13847 2431 13947 2463
rect 14003 2431 14103 2463
rect 14159 2431 14259 2463
rect 14315 2431 14415 2463
rect 14471 2513 15039 2529
rect 14471 2479 14487 2513
rect 14521 2479 14558 2513
rect 14592 2479 14629 2513
rect 14663 2479 14701 2513
rect 14735 2479 14773 2513
rect 14807 2479 14845 2513
rect 14879 2479 14917 2513
rect 14951 2479 14989 2513
rect 15023 2479 15039 2513
rect 14471 2463 15039 2479
rect 14471 2431 14571 2463
rect 14627 2431 14727 2463
rect 14783 2431 14883 2463
rect 14939 2431 15039 2463
rect 12468 2352 12668 2408
rect 12468 2318 12519 2352
rect 12553 2318 12587 2352
rect 12621 2318 12668 2352
rect 12468 2221 12668 2318
rect 12724 2323 12924 2408
rect 12724 2289 12774 2323
rect 12808 2289 12842 2323
rect 12876 2289 12924 2323
rect 12724 2221 12924 2289
rect 12468 2105 12668 2137
rect 12724 2105 12924 2137
rect 12086 2022 12942 2038
rect 12086 1988 12132 2022
rect 12166 1988 12205 2022
rect 12239 1988 12278 2022
rect 12312 1988 12351 2022
rect 12385 1988 12424 2022
rect 12458 1988 12497 2022
rect 12531 1988 12570 2022
rect 12604 1988 12642 2022
rect 12676 1988 12714 2022
rect 12748 1988 12786 2022
rect 12820 1988 12858 2022
rect 12892 1988 12942 2022
rect 12086 1972 12942 1988
rect 12086 1940 12486 1972
rect 12542 1940 12942 1972
rect 12086 1824 12486 1856
rect 12542 1824 12942 1856
rect 13223 1799 13323 1831
rect 13379 1799 13479 1831
rect 13535 1799 13635 1831
rect 13691 1799 13791 1831
rect 13847 1799 13947 1831
rect 14003 1799 14103 1831
rect 14159 1799 14259 1831
rect 14315 1799 14415 1831
rect 14471 1799 14571 1831
rect 14627 1799 14727 1831
rect 14783 1799 14883 1831
rect 14939 1799 15039 1831
<< polycont >>
rect 37627 15022 37661 15056
rect 37627 14952 37661 14986
rect 37627 14882 37661 14916
rect 37627 14812 37661 14846
rect 37627 14742 37661 14776
rect 37627 14672 37661 14706
rect 37627 14602 37661 14636
rect 37627 14532 37661 14566
rect 37627 14462 37661 14496
rect 37627 14392 37661 14426
rect 37627 14322 37661 14356
rect 37627 14252 37661 14286
rect 37627 14182 37661 14216
rect 37627 14112 37661 14146
rect 37627 14042 37661 14076
rect 37627 13972 37661 14006
rect 37627 13902 37661 13936
rect 37627 13832 37661 13866
rect 37627 13762 37661 13796
rect 37627 13692 37661 13726
rect 37627 13622 37661 13656
rect 37627 13552 37661 13586
rect 37627 13482 37661 13516
rect 37627 13412 37661 13446
rect 37627 13342 37661 13376
rect 37627 13272 37661 13306
rect 11810 2884 11844 2918
rect 11882 2884 11916 2918
rect 11954 2884 11988 2918
rect 12026 2884 12060 2918
rect 12098 2884 12132 2918
rect 12169 2884 12203 2918
rect 12240 2884 12274 2918
rect 12311 2884 12345 2918
rect 12434 2884 12468 2918
rect 12505 2884 12539 2918
rect 12576 2884 12610 2918
rect 12648 2884 12682 2918
rect 12720 2884 12754 2918
rect 12792 2884 12826 2918
rect 12864 2884 12898 2918
rect 12936 2884 12970 2918
rect 13076 2876 13110 2910
rect 13215 2884 13249 2918
rect 13309 2884 13343 2918
rect 13404 2884 13438 2918
rect 13543 2876 13577 2910
rect 13076 2808 13110 2842
rect 13543 2808 13577 2842
rect 13832 2876 13866 2910
rect 13832 2808 13866 2842
rect 14122 2867 14156 2901
rect 14122 2799 14156 2833
rect 14299 2867 14333 2901
rect 14299 2799 14333 2833
rect 14453 2867 14487 2901
rect 14453 2799 14487 2833
rect 13239 2491 13273 2525
rect 13334 2491 13368 2525
rect 13429 2491 13463 2525
rect 13551 2479 13585 2513
rect 13646 2479 13680 2513
rect 13741 2479 13775 2513
rect 13863 2479 13897 2513
rect 13935 2479 13969 2513
rect 14007 2479 14041 2513
rect 14079 2479 14113 2513
rect 14151 2479 14185 2513
rect 14223 2479 14257 2513
rect 14294 2479 14328 2513
rect 14365 2479 14399 2513
rect 14487 2479 14521 2513
rect 14558 2479 14592 2513
rect 14629 2479 14663 2513
rect 14701 2479 14735 2513
rect 14773 2479 14807 2513
rect 14845 2479 14879 2513
rect 14917 2479 14951 2513
rect 14989 2479 15023 2513
rect 12519 2318 12553 2352
rect 12587 2318 12621 2352
rect 12774 2289 12808 2323
rect 12842 2289 12876 2323
rect 12132 1988 12166 2022
rect 12205 1988 12239 2022
rect 12278 1988 12312 2022
rect 12351 1988 12385 2022
rect 12424 1988 12458 2022
rect 12497 1988 12531 2022
rect 12570 1988 12604 2022
rect 12642 1988 12676 2022
rect 12714 1988 12748 2022
rect 12786 1988 12820 2022
rect 12858 1988 12892 2022
<< locali >>
rect 35625 15083 35647 15117
rect 35693 15083 35719 15117
rect 35761 15083 35791 15117
rect 35829 15083 35863 15117
rect 35897 15083 35931 15117
rect 35969 15083 35999 15117
rect 36041 15083 36067 15117
rect 36113 15083 36135 15117
rect 36185 15083 36203 15117
rect 36257 15083 36271 15117
rect 36329 15083 36339 15117
rect 36401 15083 36407 15117
rect 36473 15083 36475 15117
rect 36509 15083 36511 15117
rect 36577 15083 36583 15117
rect 36645 15083 36655 15117
rect 36713 15083 36727 15117
rect 36781 15083 36799 15117
rect 36849 15083 36871 15117
rect 36917 15083 36943 15117
rect 36985 15083 37015 15117
rect 37053 15083 37087 15117
rect 37121 15083 37155 15117
rect 37193 15083 37223 15117
rect 37265 15083 37291 15117
rect 37337 15083 37359 15117
rect 37409 15083 37427 15117
rect 37481 15083 37495 15117
rect 37627 15060 37661 15072
rect 37627 14987 37661 15022
rect 35625 14927 35647 14961
rect 35693 14927 35719 14961
rect 35761 14927 35791 14961
rect 35829 14927 35863 14961
rect 35897 14927 35931 14961
rect 35969 14927 35999 14961
rect 36041 14927 36067 14961
rect 36113 14927 36135 14961
rect 36185 14927 36203 14961
rect 36257 14927 36271 14961
rect 36329 14927 36339 14961
rect 36401 14927 36407 14961
rect 36473 14927 36475 14961
rect 36509 14927 36511 14961
rect 36577 14927 36583 14961
rect 36645 14927 36655 14961
rect 36713 14927 36727 14961
rect 36781 14927 36799 14961
rect 36849 14927 36871 14961
rect 36917 14927 36943 14961
rect 36985 14927 37015 14961
rect 37053 14927 37087 14961
rect 37121 14927 37155 14961
rect 37193 14927 37223 14961
rect 37265 14927 37291 14961
rect 37337 14927 37359 14961
rect 37409 14927 37427 14961
rect 37481 14927 37495 14961
rect 37627 14916 37661 14952
rect 37627 14846 37661 14880
rect 35625 14771 35647 14805
rect 35693 14771 35719 14805
rect 35761 14771 35791 14805
rect 35829 14771 35863 14805
rect 35897 14771 35931 14805
rect 35969 14771 35999 14805
rect 36041 14771 36067 14805
rect 36113 14771 36135 14805
rect 36185 14771 36203 14805
rect 36257 14771 36271 14805
rect 36329 14771 36339 14805
rect 36401 14771 36407 14805
rect 36473 14771 36475 14805
rect 36509 14771 36511 14805
rect 36577 14771 36583 14805
rect 36645 14771 36655 14805
rect 36713 14771 36727 14805
rect 36781 14771 36799 14805
rect 36849 14771 36871 14805
rect 36917 14771 36943 14805
rect 36985 14771 37015 14805
rect 37053 14771 37087 14805
rect 37121 14771 37155 14805
rect 37193 14771 37223 14805
rect 37265 14771 37291 14805
rect 37337 14771 37359 14805
rect 37409 14771 37427 14805
rect 37481 14771 37495 14805
rect 37627 14776 37661 14807
rect 37627 14706 37661 14734
rect 35625 14615 35647 14649
rect 35693 14615 35719 14649
rect 35761 14615 35791 14649
rect 35829 14615 35863 14649
rect 35897 14615 35931 14649
rect 35969 14615 35999 14649
rect 36041 14615 36067 14649
rect 36113 14615 36135 14649
rect 36185 14615 36203 14649
rect 36257 14615 36271 14649
rect 36329 14615 36339 14649
rect 36401 14615 36407 14649
rect 36473 14615 36475 14649
rect 36509 14615 36511 14649
rect 36577 14615 36583 14649
rect 36645 14615 36655 14649
rect 36713 14615 36727 14649
rect 36781 14615 36799 14649
rect 36849 14615 36871 14649
rect 36917 14615 36943 14649
rect 36985 14615 37015 14649
rect 37053 14615 37087 14649
rect 37121 14615 37155 14649
rect 37193 14615 37223 14649
rect 37265 14615 37291 14649
rect 37337 14615 37359 14649
rect 37409 14615 37427 14649
rect 37481 14615 37495 14649
rect 37627 14636 37661 14661
rect 37627 14566 37661 14588
rect 37627 14496 37661 14515
rect 35625 14459 35647 14493
rect 35693 14459 35719 14493
rect 35761 14459 35791 14493
rect 35829 14459 35863 14493
rect 35897 14459 35931 14493
rect 35969 14459 35999 14493
rect 36041 14459 36067 14493
rect 36113 14459 36135 14493
rect 36185 14459 36203 14493
rect 36257 14459 36271 14493
rect 36329 14459 36339 14493
rect 36401 14459 36407 14493
rect 36473 14459 36475 14493
rect 36509 14459 36511 14493
rect 36577 14459 36583 14493
rect 36645 14459 36655 14493
rect 36713 14459 36727 14493
rect 36781 14459 36799 14493
rect 36849 14459 36871 14493
rect 36917 14459 36943 14493
rect 36985 14459 37015 14493
rect 37053 14459 37087 14493
rect 37121 14459 37155 14493
rect 37193 14459 37223 14493
rect 37265 14459 37291 14493
rect 37337 14459 37359 14493
rect 37409 14459 37427 14493
rect 37481 14459 37495 14493
rect 37627 14426 37661 14442
rect 37627 14356 37661 14369
rect 35625 14303 35647 14337
rect 35693 14303 35719 14337
rect 35761 14303 35791 14337
rect 35829 14303 35863 14337
rect 35897 14303 35931 14337
rect 35969 14303 35999 14337
rect 36041 14303 36067 14337
rect 36113 14303 36135 14337
rect 36185 14303 36203 14337
rect 36257 14303 36271 14337
rect 36329 14303 36339 14337
rect 36401 14303 36407 14337
rect 36473 14303 36475 14337
rect 36509 14303 36511 14337
rect 36577 14303 36583 14337
rect 36645 14303 36655 14337
rect 36713 14303 36727 14337
rect 36781 14303 36799 14337
rect 36849 14303 36871 14337
rect 36917 14303 36943 14337
rect 36985 14303 37015 14337
rect 37053 14303 37087 14337
rect 37121 14303 37155 14337
rect 37193 14303 37223 14337
rect 37265 14303 37291 14337
rect 37337 14303 37359 14337
rect 37409 14303 37427 14337
rect 37481 14303 37495 14337
rect 37627 14286 37661 14296
rect 37627 14216 37661 14223
rect 35625 14147 35647 14181
rect 35693 14147 35719 14181
rect 35761 14147 35791 14181
rect 35829 14147 35863 14181
rect 35897 14147 35931 14181
rect 35969 14147 35999 14181
rect 36041 14147 36067 14181
rect 36113 14147 36135 14181
rect 36185 14147 36203 14181
rect 36257 14147 36271 14181
rect 36329 14147 36339 14181
rect 36401 14147 36407 14181
rect 36473 14147 36475 14181
rect 36509 14147 36511 14181
rect 36577 14147 36583 14181
rect 36645 14147 36655 14181
rect 36713 14147 36727 14181
rect 36781 14147 36799 14181
rect 36849 14147 36871 14181
rect 36917 14147 36943 14181
rect 36985 14147 37015 14181
rect 37053 14147 37087 14181
rect 37121 14147 37155 14181
rect 37193 14147 37223 14181
rect 37265 14147 37291 14181
rect 37337 14147 37359 14181
rect 37409 14147 37427 14181
rect 37481 14147 37495 14181
rect 37627 14146 37661 14150
rect 37627 14111 37661 14112
rect 37627 14076 37661 14077
rect 37627 14038 37661 14042
rect 35625 13991 35647 14025
rect 35693 13991 35719 14025
rect 35761 13991 35791 14025
rect 35829 13991 35863 14025
rect 35897 13991 35931 14025
rect 35969 13991 35999 14025
rect 36041 13991 36067 14025
rect 36113 13991 36135 14025
rect 36185 13991 36203 14025
rect 36257 13991 36271 14025
rect 36329 13991 36339 14025
rect 36401 13991 36407 14025
rect 36473 13991 36475 14025
rect 36509 13991 36511 14025
rect 36577 13991 36583 14025
rect 36645 13991 36655 14025
rect 36713 13991 36727 14025
rect 36781 13991 36799 14025
rect 36849 13991 36871 14025
rect 36917 13991 36943 14025
rect 36985 13991 37015 14025
rect 37053 13991 37087 14025
rect 37121 13991 37155 14025
rect 37193 13991 37223 14025
rect 37265 13991 37291 14025
rect 37337 13991 37359 14025
rect 37409 13991 37427 14025
rect 37481 13991 37495 14025
rect 37627 13965 37661 13972
rect 37627 13892 37661 13902
rect 35625 13835 35647 13869
rect 35693 13835 35719 13869
rect 35761 13835 35791 13869
rect 35829 13835 35863 13869
rect 35897 13835 35931 13869
rect 35969 13835 35999 13869
rect 36041 13835 36067 13869
rect 36113 13835 36135 13869
rect 36185 13835 36203 13869
rect 36257 13835 36271 13869
rect 36329 13835 36339 13869
rect 36401 13835 36407 13869
rect 36473 13835 36475 13869
rect 36509 13835 36511 13869
rect 36577 13835 36583 13869
rect 36645 13835 36655 13869
rect 36713 13835 36727 13869
rect 36781 13835 36799 13869
rect 36849 13835 36871 13869
rect 36917 13835 36943 13869
rect 36985 13835 37015 13869
rect 37053 13835 37087 13869
rect 37121 13835 37155 13869
rect 37193 13835 37223 13869
rect 37265 13835 37291 13869
rect 37337 13835 37359 13869
rect 37409 13835 37427 13869
rect 37481 13835 37495 13869
rect 37627 13819 37661 13832
rect 37627 13746 37661 13762
rect 35625 13679 35647 13713
rect 35693 13679 35719 13713
rect 35761 13679 35791 13713
rect 35829 13679 35863 13713
rect 35897 13679 35931 13713
rect 35969 13679 35999 13713
rect 36041 13679 36067 13713
rect 36113 13679 36135 13713
rect 36185 13679 36203 13713
rect 36257 13679 36271 13713
rect 36329 13679 36339 13713
rect 36401 13679 36407 13713
rect 36473 13679 36475 13713
rect 36509 13679 36511 13713
rect 36577 13679 36583 13713
rect 36645 13679 36655 13713
rect 36713 13679 36727 13713
rect 36781 13679 36799 13713
rect 36849 13679 36871 13713
rect 36917 13679 36943 13713
rect 36985 13679 37015 13713
rect 37053 13679 37087 13713
rect 37121 13679 37155 13713
rect 37193 13679 37223 13713
rect 37265 13679 37291 13713
rect 37337 13679 37359 13713
rect 37409 13679 37427 13713
rect 37481 13679 37495 13713
rect 37627 13672 37661 13692
rect 37627 13598 37661 13622
rect 35625 13523 35647 13557
rect 35693 13523 35719 13557
rect 35761 13523 35791 13557
rect 35829 13523 35863 13557
rect 35897 13523 35931 13557
rect 35969 13523 35999 13557
rect 36041 13523 36067 13557
rect 36113 13523 36135 13557
rect 36185 13523 36203 13557
rect 36257 13523 36271 13557
rect 36329 13523 36339 13557
rect 36401 13523 36407 13557
rect 36473 13523 36475 13557
rect 36509 13523 36511 13557
rect 36577 13523 36583 13557
rect 36645 13523 36655 13557
rect 36713 13523 36727 13557
rect 36781 13523 36799 13557
rect 36849 13523 36871 13557
rect 36917 13523 36943 13557
rect 36985 13523 37015 13557
rect 37053 13523 37087 13557
rect 37121 13523 37155 13557
rect 37193 13523 37223 13557
rect 37265 13523 37291 13557
rect 37337 13523 37359 13557
rect 37409 13523 37427 13557
rect 37481 13523 37495 13557
rect 37627 13524 37661 13552
rect 37627 13450 37661 13482
rect 35625 13367 35647 13401
rect 35693 13367 35719 13401
rect 35761 13367 35791 13401
rect 35829 13367 35863 13401
rect 35897 13367 35931 13401
rect 35969 13367 35999 13401
rect 36041 13367 36067 13401
rect 36113 13367 36135 13401
rect 36185 13367 36203 13401
rect 36257 13367 36271 13401
rect 36329 13367 36339 13401
rect 36401 13367 36407 13401
rect 36473 13367 36475 13401
rect 36509 13367 36511 13401
rect 36577 13367 36583 13401
rect 36645 13367 36655 13401
rect 36713 13367 36727 13401
rect 36781 13367 36799 13401
rect 36849 13367 36871 13401
rect 36917 13367 36943 13401
rect 36985 13367 37015 13401
rect 37053 13367 37087 13401
rect 37121 13367 37155 13401
rect 37193 13367 37223 13401
rect 37265 13367 37291 13401
rect 37337 13367 37359 13401
rect 37409 13367 37427 13401
rect 37481 13367 37495 13401
rect 37627 13376 37661 13412
rect 37627 13306 37661 13342
rect 37627 13256 37661 13268
rect 35625 13211 35647 13245
rect 35693 13211 35719 13245
rect 35761 13211 35791 13245
rect 35829 13211 35863 13245
rect 35897 13211 35931 13245
rect 35969 13211 35999 13245
rect 36041 13211 36067 13245
rect 36113 13211 36135 13245
rect 36185 13211 36203 13245
rect 36257 13211 36271 13245
rect 36329 13211 36339 13245
rect 36401 13211 36407 13245
rect 36473 13211 36475 13245
rect 36509 13211 36511 13245
rect 36577 13211 36583 13245
rect 36645 13211 36655 13245
rect 36713 13211 36727 13245
rect 36781 13211 36799 13245
rect 36849 13211 36871 13245
rect 36917 13211 36943 13245
rect 36985 13211 37015 13245
rect 37053 13211 37087 13245
rect 37121 13211 37155 13245
rect 37193 13211 37223 13245
rect 37265 13211 37291 13245
rect 37337 13211 37359 13245
rect 37409 13211 37427 13245
rect 37481 13211 37495 13245
rect 11721 3640 11745 3674
rect 11786 3640 11815 3674
rect 11860 3640 11885 3674
rect 11934 3640 11955 3674
rect 12008 3640 12025 3674
rect 12082 3640 12095 3674
rect 12156 3640 12165 3674
rect 12230 3640 12235 3674
rect 12269 3640 12270 3674
rect 12304 3640 12305 3674
rect 12339 3640 12344 3674
rect 12409 3640 12418 3674
rect 12479 3640 12492 3674
rect 12549 3640 12566 3674
rect 12619 3640 12640 3674
rect 12689 3640 12714 3674
rect 12759 3640 12788 3674
rect 12829 3640 12862 3674
rect 12898 3640 12933 3674
rect 12970 3640 13002 3674
rect 13044 3640 13071 3674
rect 13118 3640 13140 3674
rect 13192 3640 13209 3674
rect 13266 3640 13278 3674
rect 13340 3640 13347 3674
rect 13414 3640 13416 3674
rect 13450 3640 13454 3674
rect 13519 3640 13528 3674
rect 13588 3640 13602 3674
rect 13657 3640 13676 3674
rect 13726 3640 13750 3674
rect 13795 3640 13824 3674
rect 13864 3640 13898 3674
rect 13933 3640 13968 3674
rect 14005 3640 14037 3674
rect 14078 3640 14106 3674
rect 14151 3640 14175 3674
rect 14224 3640 14244 3674
rect 14297 3640 14313 3674
rect 14370 3640 14382 3674
rect 14443 3640 14451 3674
rect 14516 3640 14520 3674
rect 14554 3640 14555 3674
rect 14623 3640 14647 3674
rect 11749 3567 11783 3570
rect 11749 3494 11783 3520
rect 11749 3422 11783 3452
rect 11749 3350 11783 3384
rect 11749 3282 11783 3316
rect 11749 3214 11783 3244
rect 11749 3146 11783 3180
rect 11749 3078 11783 3112
rect 11749 3028 11783 3044
rect 11905 3567 11939 3570
rect 11905 3486 11939 3520
rect 11905 3418 11939 3445
rect 11905 3350 11939 3357
rect 11905 3303 11939 3316
rect 11905 3215 11939 3248
rect 11905 3146 11939 3180
rect 11905 3078 11939 3112
rect 11905 3028 11939 3044
rect 12061 3567 12095 3570
rect 12061 3486 12095 3520
rect 12061 3418 12095 3445
rect 12061 3350 12095 3357
rect 12061 3303 12095 3316
rect 12061 3215 12095 3248
rect 12061 3146 12095 3180
rect 12061 3078 12095 3112
rect 12061 3028 12095 3044
rect 12217 3554 12251 3570
rect 12217 3486 12251 3520
rect 12217 3418 12251 3452
rect 12217 3350 12251 3357
rect 12217 3313 12251 3316
rect 12217 3235 12251 3248
rect 12217 3157 12251 3180
rect 12217 3078 12251 3112
rect 12217 3028 12251 3044
rect 12373 3567 12407 3570
rect 12373 3486 12407 3520
rect 12373 3418 12407 3450
rect 12373 3350 12407 3368
rect 12373 3282 12407 3286
rect 12373 3214 12407 3248
rect 12373 3146 12407 3180
rect 12373 3078 12407 3112
rect 12373 3028 12407 3044
rect 12529 3567 12563 3570
rect 12529 3486 12563 3520
rect 12529 3418 12563 3450
rect 12529 3350 12563 3368
rect 12529 3282 12563 3286
rect 12529 3214 12563 3248
rect 12529 3146 12563 3180
rect 12529 3078 12563 3112
rect 12529 3028 12563 3044
rect 12685 3567 12719 3570
rect 12685 3486 12719 3520
rect 12685 3418 12719 3450
rect 12685 3350 12719 3368
rect 12685 3282 12719 3286
rect 12685 3214 12719 3248
rect 12841 3554 12875 3570
rect 12841 3486 12875 3520
rect 12841 3418 12875 3452
rect 12841 3350 12875 3384
rect 12841 3282 12875 3316
rect 12841 3214 12875 3248
rect 12997 3567 13031 3570
rect 12997 3491 13031 3520
rect 12997 3418 13031 3452
rect 12997 3350 13031 3382
rect 12997 3282 13031 3307
rect 13153 3554 13187 3570
rect 13153 3486 13187 3520
rect 13153 3418 13187 3452
rect 13153 3350 13187 3384
rect 13153 3282 13187 3316
rect 12997 3214 13031 3248
rect 12685 3146 12719 3180
rect 12875 3180 12891 3211
rect 12853 3177 12891 3180
rect 12685 3078 12719 3112
rect 12685 3028 12719 3044
rect 12841 3146 12875 3177
rect 12841 3078 12875 3112
rect 12841 3028 12875 3044
rect 12997 3146 13031 3180
rect 12997 3078 13031 3112
rect 12997 3028 13031 3044
rect 13065 3220 13075 3249
rect 13109 3220 13119 3249
rect 13065 3182 13119 3220
rect 13065 3148 13075 3182
rect 13109 3148 13119 3182
rect 11794 2884 11810 2918
rect 11872 2884 11882 2918
rect 11916 2884 11924 2918
rect 11988 2884 12010 2918
rect 12060 2884 12096 2918
rect 12132 2884 12169 2918
rect 12216 2884 12240 2918
rect 12301 2884 12311 2918
rect 12345 2884 12361 2918
rect 12418 2884 12434 2918
rect 12468 2884 12476 2918
rect 12539 2884 12559 2918
rect 12610 2884 12642 2918
rect 12682 2884 12720 2918
rect 12759 2884 12792 2918
rect 12842 2884 12864 2918
rect 12925 2884 12936 2918
rect 12970 2884 12986 2918
rect 13065 2910 13119 3148
rect 13153 3214 13187 3248
rect 13153 3146 13187 3180
rect 13153 3078 13187 3112
rect 13153 3028 13187 3044
rect 13277 3554 13383 3570
rect 13277 3520 13309 3554
rect 13343 3520 13383 3554
rect 13277 3486 13383 3520
rect 13277 3452 13309 3486
rect 13343 3452 13383 3486
rect 13277 3418 13383 3452
rect 13277 3384 13309 3418
rect 13343 3384 13383 3418
rect 13277 3350 13383 3384
rect 13277 3316 13309 3350
rect 13343 3316 13383 3350
rect 13277 3282 13383 3316
rect 13277 3248 13309 3282
rect 13343 3248 13383 3282
rect 13277 3214 13383 3248
rect 13277 3180 13309 3214
rect 13343 3180 13383 3214
rect 13277 3146 13383 3180
rect 13277 3112 13309 3146
rect 13343 3112 13383 3146
rect 13277 3078 13383 3112
rect 13277 3044 13309 3078
rect 13343 3044 13383 3078
rect 13277 3002 13383 3044
rect 13465 3554 13499 3570
rect 13465 3486 13499 3520
rect 13465 3418 13499 3452
rect 13465 3350 13499 3384
rect 13465 3282 13499 3316
rect 13621 3554 13655 3570
rect 13621 3486 13655 3520
rect 13621 3418 13655 3452
rect 13621 3350 13655 3384
rect 13621 3282 13655 3316
rect 13465 3214 13499 3248
rect 13465 3146 13499 3180
rect 13465 3078 13499 3112
rect 13465 3028 13499 3044
rect 13533 3254 13587 3257
rect 13533 3220 13544 3254
rect 13578 3220 13587 3254
rect 13533 3182 13587 3220
rect 13533 3148 13544 3182
rect 13578 3148 13587 3182
rect 13311 2968 13349 3002
rect 13065 2876 13076 2910
rect 13110 2876 13119 2910
rect 13199 2884 13215 2918
rect 13251 2884 13309 2918
rect 13345 2884 13404 2918
rect 13439 2884 13454 2918
rect 13533 2910 13587 3148
rect 13621 3214 13655 3248
rect 13621 3154 13655 3180
rect 13742 3554 13776 3570
rect 13742 3486 13776 3520
rect 13742 3418 13776 3452
rect 13742 3350 13776 3384
rect 13742 3282 13776 3316
rect 13742 3214 13776 3248
rect 13742 3156 13776 3180
rect 13621 3146 13625 3154
rect 13655 3112 13659 3120
rect 13621 3082 13659 3112
rect 13621 3078 13625 3082
rect 13742 3078 13776 3112
rect 13621 3028 13655 3044
rect 13742 3015 13776 3044
rect 13918 3554 13952 3570
rect 13918 3486 13952 3520
rect 13918 3418 13952 3452
rect 13918 3381 13952 3384
rect 13918 3299 13952 3316
rect 14042 3554 14076 3570
rect 14042 3486 14076 3520
rect 14042 3418 14076 3452
rect 14042 3350 14076 3384
rect 14042 3312 14076 3316
rect 14218 3554 14252 3570
rect 14218 3486 14252 3520
rect 14218 3418 14252 3452
rect 14218 3350 14252 3384
rect 14047 3282 14085 3312
rect 14076 3278 14085 3282
rect 14218 3282 14252 3316
rect 13918 3214 13952 3248
rect 13918 3146 13952 3180
rect 13918 3078 13952 3112
rect 13918 3028 13952 3044
rect 14042 3214 14076 3248
rect 14042 3146 14076 3180
rect 14042 3078 14076 3112
rect 14042 3028 14076 3044
rect 14218 3227 14252 3248
rect 14218 3154 14252 3180
rect 14218 3082 14252 3112
rect 14218 3028 14252 3044
rect 14374 3554 14408 3570
rect 14374 3486 14408 3520
rect 14374 3418 14408 3452
rect 14374 3350 14408 3384
rect 14374 3282 14408 3316
rect 14374 3214 14408 3248
rect 14374 3146 14408 3180
rect 14374 3078 14408 3112
rect 14374 3028 14408 3044
rect 14530 3554 14621 3570
rect 14564 3520 14621 3554
rect 14530 3486 14621 3520
rect 14564 3452 14621 3486
rect 14530 3418 14621 3452
rect 14564 3384 14621 3418
rect 14530 3350 14621 3384
rect 14564 3316 14621 3350
rect 14530 3282 14621 3316
rect 14564 3248 14621 3282
rect 14530 3214 14621 3248
rect 14564 3180 14621 3214
rect 14530 3146 14621 3180
rect 14564 3112 14621 3146
rect 14530 3078 14621 3112
rect 14564 3044 14621 3078
rect 14530 3028 14621 3044
rect 14931 3028 15037 3570
rect 15104 3028 15177 3570
rect 15227 3028 15333 3570
rect 15384 3028 15490 3570
rect 15538 3028 15644 3570
rect 15691 3028 15797 3570
rect 15848 3028 15954 3570
rect 16008 3028 16114 3570
rect 16159 3028 16265 3570
rect 16318 3028 16424 3570
rect 16467 3028 16573 3570
rect 16618 3028 16724 3570
rect 16775 3028 16881 3570
rect 16918 3028 17024 3570
rect 17089 3028 17195 3570
rect 17236 3028 17342 3570
rect 17383 3028 17489 3570
rect 17526 3028 17632 3570
rect 17669 3028 17775 3570
rect 14442 2994 14496 3012
rect 14441 2960 14479 2994
rect 13065 2842 13119 2876
rect 13065 2808 13076 2842
rect 13110 2808 13119 2842
rect 13065 2792 13119 2808
rect 13533 2876 13543 2910
rect 13577 2876 13587 2910
rect 13533 2842 13587 2876
rect 13533 2808 13543 2842
rect 13577 2808 13587 2842
rect 13533 2792 13587 2808
rect 13621 2919 13774 2925
rect 13621 2885 13636 2919
rect 13670 2885 13708 2919
rect 13742 2885 13774 2919
rect 12304 2743 12574 2749
rect 12304 2709 12317 2743
rect 12351 2709 12423 2743
rect 12457 2709 12528 2743
rect 12562 2709 12574 2743
rect 13621 2743 13774 2885
rect 13621 2709 13636 2743
rect 13670 2709 13708 2743
rect 13742 2709 13774 2743
rect 13808 2910 14013 2928
rect 13808 2876 13832 2910
rect 13866 2876 14013 2910
rect 13808 2842 14013 2876
rect 13808 2808 13832 2842
rect 13866 2808 14013 2842
rect 12304 2648 12574 2709
rect 12935 2661 13033 2675
rect 12116 2596 12270 2602
rect 12116 2562 12131 2596
rect 12165 2562 12224 2596
rect 12258 2562 12270 2596
rect 12116 2514 12270 2562
rect 12116 2480 12131 2514
rect 12165 2480 12224 2514
rect 12258 2480 12270 2514
rect 11954 2237 12075 2257
rect 11954 2203 12001 2237
rect 12035 2203 12075 2237
rect 11954 2160 12075 2203
rect 11954 2126 12001 2160
rect 12035 2126 12075 2160
rect 11954 2083 12075 2126
rect 11954 2049 12001 2083
rect 12035 2049 12075 2083
rect 11954 1928 12075 2049
rect 12116 2022 12270 2480
rect 12304 2480 12457 2648
rect 12935 2627 12981 2661
rect 13015 2627 13033 2661
rect 12520 2566 12544 2600
rect 12578 2596 12614 2600
rect 12648 2596 12684 2600
rect 12718 2596 12753 2600
rect 12787 2596 12822 2600
rect 12578 2566 12583 2596
rect 12648 2566 12656 2596
rect 12718 2566 12729 2596
rect 12787 2566 12801 2596
rect 12856 2566 12880 2600
rect 12935 2568 13033 2627
rect 13808 2667 14013 2808
rect 14089 2919 14209 2925
rect 14089 2885 14095 2919
rect 14129 2901 14167 2919
rect 14156 2885 14167 2901
rect 14201 2885 14209 2919
rect 14089 2867 14122 2885
rect 14156 2867 14209 2885
rect 14299 2901 14333 2917
rect 14442 2901 14496 2960
rect 14089 2833 14209 2867
rect 14333 2867 14347 2883
rect 14309 2849 14347 2867
rect 14442 2867 14453 2901
rect 14487 2867 14496 2901
rect 14089 2799 14122 2833
rect 14156 2799 14209 2833
rect 14089 2778 14209 2799
rect 14299 2833 14333 2849
rect 14299 2783 14333 2799
rect 14442 2833 14496 2867
rect 14442 2799 14453 2833
rect 14487 2799 14496 2833
rect 14442 2772 14496 2799
rect 14547 2696 14621 3028
rect 14547 2670 14553 2696
rect 13808 2633 13820 2667
rect 13854 2633 13894 2667
rect 13928 2633 13967 2667
rect 14001 2633 14013 2667
rect 14587 2662 14625 2696
rect 13808 2620 14013 2633
rect 18493 2623 18536 2657
rect 18570 2623 18613 2657
rect 18647 2623 18689 2657
rect 18723 2623 18765 2657
rect 18799 2623 18841 2657
rect 18875 2623 18917 2657
rect 18951 2623 18993 2657
rect 19027 2623 19069 2657
rect 19103 2623 19145 2657
rect 19179 2623 19221 2657
rect 19255 2623 19297 2657
rect 19331 2623 19373 2657
rect 19407 2623 19449 2657
rect 19483 2623 19525 2657
rect 19559 2623 19601 2657
rect 19635 2623 19677 2657
rect 12304 2446 12423 2480
rect 12304 2284 12457 2446
rect 12617 2562 12656 2566
rect 12690 2562 12729 2566
rect 12763 2562 12801 2566
rect 12583 2514 12835 2562
rect 12617 2480 12656 2514
rect 12690 2480 12729 2514
rect 12763 2480 12801 2514
rect 12583 2446 12679 2480
rect 12713 2446 12835 2480
rect 12583 2430 12835 2446
rect 12935 2534 12981 2568
rect 13015 2534 13033 2568
rect 12935 2480 13033 2534
rect 13223 2491 13239 2525
rect 13273 2491 13334 2525
rect 13368 2491 13429 2525
rect 13463 2491 13479 2525
rect 12969 2475 13033 2480
rect 12969 2446 12981 2475
rect 12935 2441 12981 2446
rect 13015 2441 13033 2475
rect 12935 2396 13033 2441
rect 12503 2382 13033 2396
rect 12503 2357 12981 2382
rect 12503 2352 12637 2357
rect 12503 2318 12519 2352
rect 12553 2318 12587 2352
rect 12621 2318 12637 2352
rect 12935 2348 12981 2357
rect 13015 2348 13033 2382
rect 12758 2302 12774 2323
rect 12808 2302 12842 2323
rect 12758 2284 12761 2302
rect 12808 2289 12833 2302
rect 12876 2289 12892 2323
rect 12304 2268 12761 2284
rect 12795 2268 12833 2289
rect 12867 2268 12892 2289
rect 12304 2237 12892 2268
rect 12304 2183 12457 2237
rect 12304 2149 12423 2183
rect 12304 2130 12457 2149
rect 12640 2183 12766 2203
rect 12640 2149 12679 2183
rect 12713 2149 12766 2183
rect 12640 2124 12766 2149
rect 12935 2183 13033 2348
rect 12969 2149 13033 2183
rect 12935 2133 13033 2149
rect 13178 2353 13212 2369
rect 13178 2285 13212 2319
rect 13178 2217 13212 2251
rect 13178 2149 13212 2183
rect 12640 2090 12645 2124
rect 12679 2090 12717 2124
rect 12751 2090 12766 2124
rect 12640 2079 12766 2090
rect 13178 2081 13212 2115
rect 12953 2070 13073 2079
rect 12953 2036 12962 2070
rect 12996 2036 13034 2070
rect 13068 2036 13073 2070
rect 12116 1988 12132 2022
rect 12166 1988 12205 2022
rect 12239 1988 12278 2022
rect 12312 1988 12351 2022
rect 12385 1988 12424 2022
rect 12458 1988 12497 2022
rect 12531 1988 12570 2022
rect 12604 1988 12642 2022
rect 12676 1988 12714 2022
rect 12748 1988 12786 2022
rect 12820 1988 12858 2022
rect 12892 1988 12908 2022
rect 11954 1894 12041 1928
rect 12497 1928 12531 1944
rect 11954 1863 12075 1894
rect 12529 1883 12531 1894
rect 12495 1878 12531 1883
rect 12953 1928 13073 2036
rect 12987 1894 13073 1928
rect 12495 1845 12529 1878
rect 12953 1860 13073 1894
rect 13246 2222 13300 2491
rect 13246 2188 13254 2222
rect 13288 2188 13300 2222
rect 13246 2150 13300 2188
rect 13246 2116 13254 2150
rect 13288 2116 13300 2150
rect 13246 2061 13300 2116
rect 13334 2385 13368 2423
rect 13334 2285 13368 2319
rect 13334 2217 13368 2251
rect 13334 2149 13368 2183
rect 13334 2081 13368 2115
rect 13178 2013 13212 2047
rect 13178 1945 13212 1953
rect 13178 1877 13212 1879
rect 13178 1840 13212 1843
rect 13402 2222 13456 2491
rect 13535 2479 13551 2513
rect 13585 2488 13638 2522
rect 13672 2513 13725 2522
rect 13894 2513 13942 2516
rect 13976 2513 14024 2516
rect 14058 2513 14106 2516
rect 14140 2513 14189 2516
rect 13680 2488 13725 2513
rect 13585 2479 13646 2488
rect 13680 2479 13741 2488
rect 13775 2479 13791 2513
rect 13847 2482 13860 2513
rect 13847 2479 13863 2482
rect 13897 2479 13935 2513
rect 13976 2482 14007 2513
rect 14058 2482 14079 2513
rect 14140 2482 14151 2513
rect 13969 2479 14007 2482
rect 14041 2479 14079 2482
rect 14113 2479 14151 2482
rect 14185 2482 14189 2513
rect 14223 2513 14272 2516
rect 14306 2513 14355 2516
rect 14539 2513 14586 2514
rect 14620 2513 14667 2514
rect 14185 2479 14223 2482
rect 14257 2482 14272 2513
rect 14328 2482 14355 2513
rect 14257 2479 14294 2482
rect 14328 2479 14365 2482
rect 14399 2479 14415 2513
rect 14471 2479 14487 2513
rect 14539 2480 14558 2513
rect 14620 2480 14629 2513
rect 14521 2479 14558 2480
rect 14592 2479 14629 2480
rect 14663 2480 14667 2513
rect 14701 2513 14748 2514
rect 14782 2513 14829 2514
rect 14863 2513 14910 2514
rect 14944 2513 14992 2514
rect 14663 2479 14701 2480
rect 14735 2480 14748 2513
rect 14807 2480 14829 2513
rect 14879 2480 14910 2513
rect 14735 2479 14773 2480
rect 14807 2479 14845 2480
rect 14879 2479 14917 2480
rect 14951 2479 14989 2513
rect 15026 2480 15039 2513
rect 15023 2479 15039 2480
rect 13402 2188 13412 2222
rect 13446 2188 13456 2222
rect 13402 2150 13456 2188
rect 13402 2116 13412 2150
rect 13446 2116 13456 2150
rect 13402 2061 13456 2116
rect 13490 2353 13524 2369
rect 13490 2285 13524 2319
rect 13490 2217 13524 2251
rect 13490 2149 13524 2183
rect 13490 2081 13524 2115
rect 13334 2013 13368 2047
rect 13334 1945 13368 1979
rect 13334 1877 13368 1911
rect 13334 1827 13368 1843
rect 13490 2013 13524 2047
rect 13558 2147 13612 2479
rect 13558 2113 13567 2147
rect 13601 2113 13612 2147
rect 13558 2075 13612 2113
rect 13558 2041 13567 2075
rect 13601 2041 13612 2075
rect 13646 2353 13680 2369
rect 13646 2296 13680 2319
rect 13646 2224 13680 2251
rect 13646 2149 13680 2183
rect 13646 2081 13680 2115
rect 13490 1945 13524 1953
rect 13490 1877 13524 1879
rect 13490 1840 13524 1843
rect 13646 2013 13680 2047
rect 13714 2147 13768 2479
rect 15350 2455 15384 2493
rect 13714 2113 13727 2147
rect 13761 2113 13768 2147
rect 13714 2075 13768 2113
rect 13714 2041 13727 2075
rect 13761 2041 13768 2075
rect 13802 2353 13836 2369
rect 13802 2285 13836 2319
rect 13802 2217 13836 2251
rect 13802 2149 13836 2183
rect 13802 2100 13836 2115
rect 13646 1945 13680 1979
rect 13646 1877 13680 1911
rect 13646 1827 13680 1843
rect 13802 2013 13836 2047
rect 13802 1945 13836 1979
rect 13802 1877 13836 1892
rect 13802 1840 13836 1843
rect 13958 2355 13959 2369
rect 13958 2353 13993 2355
rect 13992 2319 13993 2353
rect 13958 2313 13993 2319
rect 13958 2285 13959 2313
rect 13992 2251 13993 2279
rect 13958 2237 13993 2251
rect 13958 2217 13959 2237
rect 14114 2353 14148 2369
rect 14114 2285 14148 2319
rect 14114 2217 14148 2251
rect 13958 2149 13992 2183
rect 13958 2081 13992 2115
rect 13958 2013 13992 2047
rect 13958 1945 13992 1979
rect 13958 1877 13992 1911
rect 13958 1827 13992 1843
rect 14114 2149 14148 2183
rect 14114 2081 14148 2115
rect 14114 2013 14148 2022
rect 14114 1945 14148 1950
rect 14114 1877 14148 1878
rect 14114 1840 14148 1843
rect 14270 2353 14304 2355
rect 14270 2313 14304 2319
rect 14270 2237 14304 2251
rect 14270 2149 14304 2183
rect 14270 2081 14304 2115
rect 14270 2013 14304 2047
rect 14270 1945 14304 1979
rect 14270 1877 14304 1911
rect 14270 1827 14304 1843
rect 14426 2353 14460 2369
rect 14426 2285 14460 2319
rect 14426 2217 14460 2251
rect 14426 2149 14460 2183
rect 14426 2081 14460 2115
rect 14426 2013 14460 2022
rect 14426 1945 14460 1950
rect 14426 1877 14460 1878
rect 14426 1840 14460 1843
rect 14582 2355 14583 2369
rect 14582 2353 14617 2355
rect 14616 2319 14617 2353
rect 14582 2313 14617 2319
rect 14582 2285 14583 2313
rect 14616 2251 14617 2279
rect 14582 2237 14617 2251
rect 14582 2217 14583 2237
rect 14738 2353 14772 2369
rect 14738 2285 14772 2319
rect 14738 2217 14772 2251
rect 14582 2149 14616 2183
rect 14582 2081 14616 2115
rect 14582 2013 14616 2047
rect 14582 1945 14616 1979
rect 14582 1877 14616 1911
rect 14582 1827 14616 1843
rect 14738 2149 14772 2183
rect 14738 2081 14772 2115
rect 14738 2013 14772 2022
rect 14738 1945 14772 1950
rect 14738 1877 14772 1878
rect 14738 1840 14772 1843
rect 14894 2353 14928 2355
rect 14894 2313 14928 2319
rect 14894 2237 14928 2251
rect 14894 2149 14928 2183
rect 14894 2081 14928 2115
rect 14894 2013 14928 2047
rect 14894 1945 14928 1979
rect 14894 1877 14928 1911
rect 14894 1827 14928 1843
rect 15050 2353 15084 2369
rect 15050 2285 15084 2319
rect 15385 2298 15454 2498
rect 15457 2454 15491 2492
rect 16410 2455 16444 2493
rect 17651 2439 17689 2473
rect 16410 2412 16444 2421
rect 16656 2333 16694 2367
rect 16960 2263 17006 2297
rect 17252 2263 17298 2297
rect 18476 2260 18515 2294
rect 18549 2260 18588 2294
rect 18622 2260 18661 2294
rect 18695 2260 18734 2294
rect 18768 2260 18807 2294
rect 18841 2260 18880 2294
rect 18914 2260 18953 2294
rect 18987 2260 19026 2294
rect 19060 2260 19099 2294
rect 19133 2260 19172 2294
rect 19206 2260 19245 2294
rect 19279 2260 19318 2294
rect 19352 2260 19391 2294
rect 19425 2260 19464 2294
rect 19498 2260 19537 2294
rect 19571 2260 19610 2294
rect 19644 2260 19682 2294
rect 19716 2260 19754 2294
rect 15050 2217 15084 2251
rect 16240 2196 16278 2230
rect 15050 2149 15084 2183
rect 16832 2182 16870 2216
rect 15050 2081 15084 2115
rect 15927 2109 15966 2143
rect 16246 2109 16285 2143
rect 20468 2114 20507 2148
rect 20541 2114 20580 2148
rect 20614 2114 20653 2148
rect 20687 2114 20726 2148
rect 20760 2114 20799 2148
rect 20833 2114 20872 2148
rect 20906 2114 20945 2148
rect 20979 2114 21018 2148
rect 21052 2114 21091 2148
rect 21125 2114 21164 2148
rect 21198 2114 21237 2148
rect 21271 2114 21310 2148
rect 21344 2114 21383 2148
rect 21417 2114 21456 2148
rect 21490 2114 21529 2148
rect 21563 2114 21602 2148
rect 21636 2114 21675 2148
rect 21709 2114 21748 2148
rect 21782 2114 21821 2148
rect 21855 2114 21894 2148
rect 21928 2114 21967 2148
rect 22001 2114 22040 2148
rect 22074 2114 22113 2148
rect 22147 2114 22185 2148
rect 22219 2114 22257 2148
rect 22291 2114 22329 2148
rect 22363 2114 22401 2148
rect 22435 2114 22473 2148
rect 22507 2114 22545 2148
rect 22579 2114 22617 2148
rect 22651 2114 22689 2148
rect 22723 2114 22761 2148
rect 22795 2114 22833 2148
rect 22867 2114 22905 2148
rect 22939 2114 22977 2148
rect 23011 2114 23049 2148
rect 23083 2114 23121 2148
rect 23155 2114 23193 2148
rect 23227 2114 23265 2148
rect 23299 2114 23337 2148
rect 23371 2114 23409 2148
rect 23443 2114 23481 2148
rect 23515 2114 23553 2148
rect 16098 2033 16137 2067
rect 15050 2013 15084 2022
rect 15050 1945 15084 1950
rect 15050 1877 15084 1878
rect 15050 1840 15084 1843
rect 15404 1959 15465 1993
rect 15499 1959 15559 1993
rect 15370 1873 15593 1959
rect 16411 1915 16445 1953
rect 18493 1941 18537 1975
rect 18571 1941 18615 1975
rect 18649 1941 18693 1975
rect 18727 1941 18771 1975
rect 18805 1941 18848 1975
rect 18882 1941 18925 1975
rect 18959 1941 19002 1975
rect 19036 1941 19079 1975
rect 19113 1941 19156 1975
rect 19190 1941 19233 1975
rect 19267 1941 19310 1975
rect 15404 1839 15465 1873
rect 15499 1839 15559 1873
rect 12063 1723 12087 1757
rect 12121 1723 12141 1757
rect 12190 1723 12214 1757
rect 12259 1723 12287 1757
rect 12328 1723 12360 1757
rect 12397 1723 12432 1757
rect 12467 1723 12501 1757
rect 12540 1723 12570 1757
rect 12613 1723 12639 1757
rect 12686 1723 12708 1757
rect 12759 1723 12777 1757
rect 12832 1723 12846 1757
rect 12905 1723 12915 1757
rect 12978 1723 12984 1757
rect 13051 1723 13053 1757
rect 13087 1723 13090 1757
rect 13156 1723 13163 1757
rect 13225 1723 13236 1757
rect 13294 1723 13309 1757
rect 13363 1723 13382 1757
rect 13432 1723 13455 1757
rect 13501 1723 13528 1757
rect 13570 1723 13601 1757
rect 13639 1723 13674 1757
rect 13708 1723 13743 1757
rect 13781 1723 13812 1757
rect 13854 1723 13881 1757
rect 13927 1723 13950 1757
rect 14000 1723 14019 1757
rect 14073 1723 14088 1757
rect 14146 1723 14157 1757
rect 14219 1723 14226 1757
rect 14292 1723 14295 1757
rect 14329 1723 14331 1757
rect 14398 1723 14404 1757
rect 14467 1723 14477 1757
rect 14536 1723 14550 1757
rect 14605 1723 14623 1757
rect 14674 1723 14696 1757
rect 14743 1723 14769 1757
rect 14812 1723 14842 1757
rect 14881 1723 14915 1757
rect 14950 1723 14985 1757
rect 15022 1723 15054 1757
rect 15095 1723 15123 1757
rect 15168 1723 15192 1757
rect 15241 1723 15261 1757
rect 15314 1723 15329 1757
rect 15387 1723 15397 1757
rect 15460 1723 15465 1757
rect 15532 1723 15533 1757
rect 15567 1723 15570 1757
rect 15635 1723 15642 1757
rect 15703 1723 15714 1757
rect 15771 1723 15786 1757
rect 21011 1691 21051 1692
rect 21085 1691 21125 1692
rect 21159 1691 21199 1692
rect 21233 1691 21273 1692
rect 21307 1691 21347 1692
rect 21381 1691 21421 1692
rect 21455 1691 21495 1692
rect 21529 1691 21569 1692
rect 21603 1691 21643 1692
rect 21677 1691 21717 1692
rect 21751 1691 21791 1692
rect 21825 1691 21865 1692
rect 21899 1691 21939 1692
rect 21973 1691 22013 1692
rect 22047 1691 22087 1692
rect 22121 1691 22161 1692
rect 22195 1691 22235 1692
rect 22269 1691 22309 1692
rect 22343 1691 22383 1692
rect 22417 1691 22457 1692
rect 22491 1691 22531 1692
rect 22565 1691 22605 1692
rect 22639 1691 22679 1692
rect 22713 1691 22753 1692
rect 22787 1691 22827 1692
rect 22861 1691 22901 1692
rect 22935 1691 22975 1692
rect 23009 1691 23049 1692
rect 23083 1691 23123 1692
rect 23157 1691 23196 1692
rect 23230 1691 23269 1692
rect 23303 1691 23342 1692
rect 23376 1691 23415 1692
rect 23449 1691 23488 1692
rect 23522 1691 23561 1692
rect 18139 1657 18160 1691
rect 18197 1657 18232 1691
rect 18266 1657 18301 1691
rect 18338 1657 18370 1691
rect 18410 1657 18439 1691
rect 18482 1657 18508 1691
rect 18554 1657 18577 1691
rect 18626 1657 18646 1691
rect 18698 1657 18715 1691
rect 18770 1657 18784 1691
rect 18842 1657 18853 1691
rect 18914 1657 18922 1691
rect 18986 1657 18991 1691
rect 19058 1657 19060 1691
rect 19094 1657 19096 1691
rect 19163 1657 19168 1691
rect 19232 1657 19240 1691
rect 19301 1657 19312 1691
rect 19370 1657 19384 1691
rect 19439 1657 19456 1691
rect 19508 1657 19528 1691
rect 19577 1657 19600 1691
rect 19646 1657 19672 1691
rect 19715 1657 19744 1691
rect 19784 1657 19816 1691
rect 19853 1657 19888 1691
rect 19922 1657 19957 1691
rect 19994 1657 20026 1691
rect 20066 1657 20095 1691
rect 20138 1657 20164 1691
rect 20210 1657 20233 1691
rect 20282 1657 20302 1691
rect 20354 1657 20371 1691
rect 20426 1657 20440 1691
rect 20498 1657 20509 1691
rect 20570 1657 20578 1691
rect 20642 1657 20647 1691
rect 20714 1657 20716 1691
rect 20750 1657 20785 1691
rect 20819 1657 20854 1691
rect 20888 1657 20923 1691
rect 20957 1658 20977 1691
rect 21026 1658 21051 1691
rect 21095 1658 21125 1691
rect 20957 1657 20992 1658
rect 21026 1657 21061 1658
rect 21095 1657 21130 1658
rect 21164 1657 21199 1691
rect 21233 1657 21268 1691
rect 21307 1658 21337 1691
rect 21381 1658 21406 1691
rect 21455 1658 21475 1691
rect 21529 1658 21543 1691
rect 21603 1658 21611 1691
rect 21677 1658 21679 1691
rect 21302 1657 21337 1658
rect 21371 1657 21406 1658
rect 21440 1657 21475 1658
rect 21509 1657 21543 1658
rect 21577 1657 21611 1658
rect 21645 1657 21679 1658
rect 21713 1658 21717 1691
rect 21781 1658 21791 1691
rect 21849 1658 21865 1691
rect 21917 1658 21939 1691
rect 21985 1658 22013 1691
rect 21713 1657 21747 1658
rect 21781 1657 21815 1658
rect 21849 1657 21883 1658
rect 21917 1657 21951 1658
rect 21985 1657 22019 1658
rect 22053 1657 22087 1691
rect 22121 1657 22155 1691
rect 22195 1658 22223 1691
rect 22269 1658 22291 1691
rect 22343 1658 22359 1691
rect 22417 1658 22427 1691
rect 22491 1658 22495 1691
rect 22189 1657 22223 1658
rect 22257 1657 22291 1658
rect 22325 1657 22359 1658
rect 22393 1657 22427 1658
rect 22461 1657 22495 1658
rect 22529 1658 22531 1691
rect 22597 1658 22605 1691
rect 22665 1658 22679 1691
rect 22733 1658 22753 1691
rect 22801 1658 22827 1691
rect 22869 1658 22901 1691
rect 22529 1657 22563 1658
rect 22597 1657 22631 1658
rect 22665 1657 22699 1658
rect 22733 1657 22767 1658
rect 22801 1657 22835 1658
rect 22869 1657 22903 1658
rect 22937 1657 22971 1691
rect 23009 1658 23039 1691
rect 23083 1658 23107 1691
rect 23157 1658 23175 1691
rect 23230 1658 23243 1691
rect 23303 1658 23311 1691
rect 23376 1658 23379 1691
rect 23005 1657 23039 1658
rect 23073 1657 23107 1658
rect 23141 1657 23175 1658
rect 23209 1657 23243 1658
rect 23277 1657 23311 1658
rect 23345 1657 23379 1658
rect 23413 1658 23415 1691
rect 23481 1658 23488 1691
rect 23549 1658 23561 1691
rect 23413 1657 23447 1658
rect 23481 1657 23515 1658
rect 23549 1657 23583 1658
rect 23617 1657 23641 1691
<< viali >>
rect 35575 15083 35591 15117
rect 35591 15083 35609 15117
rect 35647 15083 35659 15117
rect 35659 15083 35681 15117
rect 35719 15083 35727 15117
rect 35727 15083 35753 15117
rect 35791 15083 35795 15117
rect 35795 15083 35825 15117
rect 35863 15083 35897 15117
rect 35935 15083 35965 15117
rect 35965 15083 35969 15117
rect 36007 15083 36033 15117
rect 36033 15083 36041 15117
rect 36079 15083 36101 15117
rect 36101 15083 36113 15117
rect 36151 15083 36169 15117
rect 36169 15083 36185 15117
rect 36223 15083 36237 15117
rect 36237 15083 36257 15117
rect 36295 15083 36305 15117
rect 36305 15083 36329 15117
rect 36367 15083 36373 15117
rect 36373 15083 36401 15117
rect 36439 15083 36441 15117
rect 36441 15083 36473 15117
rect 36511 15083 36543 15117
rect 36543 15083 36545 15117
rect 36583 15083 36611 15117
rect 36611 15083 36617 15117
rect 36655 15083 36679 15117
rect 36679 15083 36689 15117
rect 36727 15083 36747 15117
rect 36747 15083 36761 15117
rect 36799 15083 36815 15117
rect 36815 15083 36833 15117
rect 36871 15083 36883 15117
rect 36883 15083 36905 15117
rect 36943 15083 36951 15117
rect 36951 15083 36977 15117
rect 37015 15083 37019 15117
rect 37019 15083 37049 15117
rect 37087 15083 37121 15117
rect 37159 15083 37189 15117
rect 37189 15083 37193 15117
rect 37231 15083 37257 15117
rect 37257 15083 37265 15117
rect 37303 15083 37325 15117
rect 37325 15083 37337 15117
rect 37375 15083 37393 15117
rect 37393 15083 37409 15117
rect 37447 15083 37461 15117
rect 37461 15083 37481 15117
rect 37519 15083 37529 15117
rect 37529 15083 37553 15117
rect 37627 15056 37661 15060
rect 37627 15026 37661 15056
rect 37627 14986 37661 14987
rect 35575 14927 35591 14961
rect 35591 14927 35609 14961
rect 35647 14927 35659 14961
rect 35659 14927 35681 14961
rect 35719 14927 35727 14961
rect 35727 14927 35753 14961
rect 35791 14927 35795 14961
rect 35795 14927 35825 14961
rect 35863 14927 35897 14961
rect 35935 14927 35965 14961
rect 35965 14927 35969 14961
rect 36007 14927 36033 14961
rect 36033 14927 36041 14961
rect 36079 14927 36101 14961
rect 36101 14927 36113 14961
rect 36151 14927 36169 14961
rect 36169 14927 36185 14961
rect 36223 14927 36237 14961
rect 36237 14927 36257 14961
rect 36295 14927 36305 14961
rect 36305 14927 36329 14961
rect 36367 14927 36373 14961
rect 36373 14927 36401 14961
rect 36439 14927 36441 14961
rect 36441 14927 36473 14961
rect 36511 14927 36543 14961
rect 36543 14927 36545 14961
rect 36583 14927 36611 14961
rect 36611 14927 36617 14961
rect 36655 14927 36679 14961
rect 36679 14927 36689 14961
rect 36727 14927 36747 14961
rect 36747 14927 36761 14961
rect 36799 14927 36815 14961
rect 36815 14927 36833 14961
rect 36871 14927 36883 14961
rect 36883 14927 36905 14961
rect 36943 14927 36951 14961
rect 36951 14927 36977 14961
rect 37015 14927 37019 14961
rect 37019 14927 37049 14961
rect 37087 14927 37121 14961
rect 37159 14927 37189 14961
rect 37189 14927 37193 14961
rect 37231 14927 37257 14961
rect 37257 14927 37265 14961
rect 37303 14927 37325 14961
rect 37325 14927 37337 14961
rect 37375 14927 37393 14961
rect 37393 14927 37409 14961
rect 37447 14927 37461 14961
rect 37461 14927 37481 14961
rect 37519 14927 37529 14961
rect 37529 14927 37553 14961
rect 37627 14953 37661 14986
rect 37627 14882 37661 14914
rect 37627 14880 37661 14882
rect 37627 14812 37661 14841
rect 37627 14807 37661 14812
rect 35575 14771 35591 14805
rect 35591 14771 35609 14805
rect 35647 14771 35659 14805
rect 35659 14771 35681 14805
rect 35719 14771 35727 14805
rect 35727 14771 35753 14805
rect 35791 14771 35795 14805
rect 35795 14771 35825 14805
rect 35863 14771 35897 14805
rect 35935 14771 35965 14805
rect 35965 14771 35969 14805
rect 36007 14771 36033 14805
rect 36033 14771 36041 14805
rect 36079 14771 36101 14805
rect 36101 14771 36113 14805
rect 36151 14771 36169 14805
rect 36169 14771 36185 14805
rect 36223 14771 36237 14805
rect 36237 14771 36257 14805
rect 36295 14771 36305 14805
rect 36305 14771 36329 14805
rect 36367 14771 36373 14805
rect 36373 14771 36401 14805
rect 36439 14771 36441 14805
rect 36441 14771 36473 14805
rect 36511 14771 36543 14805
rect 36543 14771 36545 14805
rect 36583 14771 36611 14805
rect 36611 14771 36617 14805
rect 36655 14771 36679 14805
rect 36679 14771 36689 14805
rect 36727 14771 36747 14805
rect 36747 14771 36761 14805
rect 36799 14771 36815 14805
rect 36815 14771 36833 14805
rect 36871 14771 36883 14805
rect 36883 14771 36905 14805
rect 36943 14771 36951 14805
rect 36951 14771 36977 14805
rect 37015 14771 37019 14805
rect 37019 14771 37049 14805
rect 37087 14771 37121 14805
rect 37159 14771 37189 14805
rect 37189 14771 37193 14805
rect 37231 14771 37257 14805
rect 37257 14771 37265 14805
rect 37303 14771 37325 14805
rect 37325 14771 37337 14805
rect 37375 14771 37393 14805
rect 37393 14771 37409 14805
rect 37447 14771 37461 14805
rect 37461 14771 37481 14805
rect 37519 14771 37529 14805
rect 37529 14771 37553 14805
rect 37627 14742 37661 14768
rect 37627 14734 37661 14742
rect 37627 14672 37661 14695
rect 37627 14661 37661 14672
rect 35575 14615 35591 14649
rect 35591 14615 35609 14649
rect 35647 14615 35659 14649
rect 35659 14615 35681 14649
rect 35719 14615 35727 14649
rect 35727 14615 35753 14649
rect 35791 14615 35795 14649
rect 35795 14615 35825 14649
rect 35863 14615 35897 14649
rect 35935 14615 35965 14649
rect 35965 14615 35969 14649
rect 36007 14615 36033 14649
rect 36033 14615 36041 14649
rect 36079 14615 36101 14649
rect 36101 14615 36113 14649
rect 36151 14615 36169 14649
rect 36169 14615 36185 14649
rect 36223 14615 36237 14649
rect 36237 14615 36257 14649
rect 36295 14615 36305 14649
rect 36305 14615 36329 14649
rect 36367 14615 36373 14649
rect 36373 14615 36401 14649
rect 36439 14615 36441 14649
rect 36441 14615 36473 14649
rect 36511 14615 36543 14649
rect 36543 14615 36545 14649
rect 36583 14615 36611 14649
rect 36611 14615 36617 14649
rect 36655 14615 36679 14649
rect 36679 14615 36689 14649
rect 36727 14615 36747 14649
rect 36747 14615 36761 14649
rect 36799 14615 36815 14649
rect 36815 14615 36833 14649
rect 36871 14615 36883 14649
rect 36883 14615 36905 14649
rect 36943 14615 36951 14649
rect 36951 14615 36977 14649
rect 37015 14615 37019 14649
rect 37019 14615 37049 14649
rect 37087 14615 37121 14649
rect 37159 14615 37189 14649
rect 37189 14615 37193 14649
rect 37231 14615 37257 14649
rect 37257 14615 37265 14649
rect 37303 14615 37325 14649
rect 37325 14615 37337 14649
rect 37375 14615 37393 14649
rect 37393 14615 37409 14649
rect 37447 14615 37461 14649
rect 37461 14615 37481 14649
rect 37519 14615 37529 14649
rect 37529 14615 37553 14649
rect 37627 14602 37661 14622
rect 37627 14588 37661 14602
rect 37627 14532 37661 14549
rect 37627 14515 37661 14532
rect 35575 14459 35591 14493
rect 35591 14459 35609 14493
rect 35647 14459 35659 14493
rect 35659 14459 35681 14493
rect 35719 14459 35727 14493
rect 35727 14459 35753 14493
rect 35791 14459 35795 14493
rect 35795 14459 35825 14493
rect 35863 14459 35897 14493
rect 35935 14459 35965 14493
rect 35965 14459 35969 14493
rect 36007 14459 36033 14493
rect 36033 14459 36041 14493
rect 36079 14459 36101 14493
rect 36101 14459 36113 14493
rect 36151 14459 36169 14493
rect 36169 14459 36185 14493
rect 36223 14459 36237 14493
rect 36237 14459 36257 14493
rect 36295 14459 36305 14493
rect 36305 14459 36329 14493
rect 36367 14459 36373 14493
rect 36373 14459 36401 14493
rect 36439 14459 36441 14493
rect 36441 14459 36473 14493
rect 36511 14459 36543 14493
rect 36543 14459 36545 14493
rect 36583 14459 36611 14493
rect 36611 14459 36617 14493
rect 36655 14459 36679 14493
rect 36679 14459 36689 14493
rect 36727 14459 36747 14493
rect 36747 14459 36761 14493
rect 36799 14459 36815 14493
rect 36815 14459 36833 14493
rect 36871 14459 36883 14493
rect 36883 14459 36905 14493
rect 36943 14459 36951 14493
rect 36951 14459 36977 14493
rect 37015 14459 37019 14493
rect 37019 14459 37049 14493
rect 37087 14459 37121 14493
rect 37159 14459 37189 14493
rect 37189 14459 37193 14493
rect 37231 14459 37257 14493
rect 37257 14459 37265 14493
rect 37303 14459 37325 14493
rect 37325 14459 37337 14493
rect 37375 14459 37393 14493
rect 37393 14459 37409 14493
rect 37447 14459 37461 14493
rect 37461 14459 37481 14493
rect 37519 14459 37529 14493
rect 37529 14459 37553 14493
rect 37627 14462 37661 14476
rect 37627 14442 37661 14462
rect 37627 14392 37661 14403
rect 37627 14369 37661 14392
rect 35575 14303 35591 14337
rect 35591 14303 35609 14337
rect 35647 14303 35659 14337
rect 35659 14303 35681 14337
rect 35719 14303 35727 14337
rect 35727 14303 35753 14337
rect 35791 14303 35795 14337
rect 35795 14303 35825 14337
rect 35863 14303 35897 14337
rect 35935 14303 35965 14337
rect 35965 14303 35969 14337
rect 36007 14303 36033 14337
rect 36033 14303 36041 14337
rect 36079 14303 36101 14337
rect 36101 14303 36113 14337
rect 36151 14303 36169 14337
rect 36169 14303 36185 14337
rect 36223 14303 36237 14337
rect 36237 14303 36257 14337
rect 36295 14303 36305 14337
rect 36305 14303 36329 14337
rect 36367 14303 36373 14337
rect 36373 14303 36401 14337
rect 36439 14303 36441 14337
rect 36441 14303 36473 14337
rect 36511 14303 36543 14337
rect 36543 14303 36545 14337
rect 36583 14303 36611 14337
rect 36611 14303 36617 14337
rect 36655 14303 36679 14337
rect 36679 14303 36689 14337
rect 36727 14303 36747 14337
rect 36747 14303 36761 14337
rect 36799 14303 36815 14337
rect 36815 14303 36833 14337
rect 36871 14303 36883 14337
rect 36883 14303 36905 14337
rect 36943 14303 36951 14337
rect 36951 14303 36977 14337
rect 37015 14303 37019 14337
rect 37019 14303 37049 14337
rect 37087 14303 37121 14337
rect 37159 14303 37189 14337
rect 37189 14303 37193 14337
rect 37231 14303 37257 14337
rect 37257 14303 37265 14337
rect 37303 14303 37325 14337
rect 37325 14303 37337 14337
rect 37375 14303 37393 14337
rect 37393 14303 37409 14337
rect 37447 14303 37461 14337
rect 37461 14303 37481 14337
rect 37519 14303 37529 14337
rect 37529 14303 37553 14337
rect 37627 14322 37661 14330
rect 37627 14296 37661 14322
rect 37627 14252 37661 14257
rect 37627 14223 37661 14252
rect 37627 14182 37661 14184
rect 35575 14147 35591 14181
rect 35591 14147 35609 14181
rect 35647 14147 35659 14181
rect 35659 14147 35681 14181
rect 35719 14147 35727 14181
rect 35727 14147 35753 14181
rect 35791 14147 35795 14181
rect 35795 14147 35825 14181
rect 35863 14147 35897 14181
rect 35935 14147 35965 14181
rect 35965 14147 35969 14181
rect 36007 14147 36033 14181
rect 36033 14147 36041 14181
rect 36079 14147 36101 14181
rect 36101 14147 36113 14181
rect 36151 14147 36169 14181
rect 36169 14147 36185 14181
rect 36223 14147 36237 14181
rect 36237 14147 36257 14181
rect 36295 14147 36305 14181
rect 36305 14147 36329 14181
rect 36367 14147 36373 14181
rect 36373 14147 36401 14181
rect 36439 14147 36441 14181
rect 36441 14147 36473 14181
rect 36511 14147 36543 14181
rect 36543 14147 36545 14181
rect 36583 14147 36611 14181
rect 36611 14147 36617 14181
rect 36655 14147 36679 14181
rect 36679 14147 36689 14181
rect 36727 14147 36747 14181
rect 36747 14147 36761 14181
rect 36799 14147 36815 14181
rect 36815 14147 36833 14181
rect 36871 14147 36883 14181
rect 36883 14147 36905 14181
rect 36943 14147 36951 14181
rect 36951 14147 36977 14181
rect 37015 14147 37019 14181
rect 37019 14147 37049 14181
rect 37087 14147 37121 14181
rect 37159 14147 37189 14181
rect 37189 14147 37193 14181
rect 37231 14147 37257 14181
rect 37257 14147 37265 14181
rect 37303 14147 37325 14181
rect 37325 14147 37337 14181
rect 37375 14147 37393 14181
rect 37393 14147 37409 14181
rect 37447 14147 37461 14181
rect 37461 14147 37481 14181
rect 37519 14147 37529 14181
rect 37529 14147 37553 14181
rect 37627 14150 37661 14182
rect 37627 14077 37661 14111
rect 35575 13991 35591 14025
rect 35591 13991 35609 14025
rect 35647 13991 35659 14025
rect 35659 13991 35681 14025
rect 35719 13991 35727 14025
rect 35727 13991 35753 14025
rect 35791 13991 35795 14025
rect 35795 13991 35825 14025
rect 35863 13991 35897 14025
rect 35935 13991 35965 14025
rect 35965 13991 35969 14025
rect 36007 13991 36033 14025
rect 36033 13991 36041 14025
rect 36079 13991 36101 14025
rect 36101 13991 36113 14025
rect 36151 13991 36169 14025
rect 36169 13991 36185 14025
rect 36223 13991 36237 14025
rect 36237 13991 36257 14025
rect 36295 13991 36305 14025
rect 36305 13991 36329 14025
rect 36367 13991 36373 14025
rect 36373 13991 36401 14025
rect 36439 13991 36441 14025
rect 36441 13991 36473 14025
rect 36511 13991 36543 14025
rect 36543 13991 36545 14025
rect 36583 13991 36611 14025
rect 36611 13991 36617 14025
rect 36655 13991 36679 14025
rect 36679 13991 36689 14025
rect 36727 13991 36747 14025
rect 36747 13991 36761 14025
rect 36799 13991 36815 14025
rect 36815 13991 36833 14025
rect 36871 13991 36883 14025
rect 36883 13991 36905 14025
rect 36943 13991 36951 14025
rect 36951 13991 36977 14025
rect 37015 13991 37019 14025
rect 37019 13991 37049 14025
rect 37087 13991 37121 14025
rect 37159 13991 37189 14025
rect 37189 13991 37193 14025
rect 37231 13991 37257 14025
rect 37257 13991 37265 14025
rect 37303 13991 37325 14025
rect 37325 13991 37337 14025
rect 37375 13991 37393 14025
rect 37393 13991 37409 14025
rect 37447 13991 37461 14025
rect 37461 13991 37481 14025
rect 37519 13991 37529 14025
rect 37529 13991 37553 14025
rect 37627 14006 37661 14038
rect 37627 14004 37661 14006
rect 37627 13936 37661 13965
rect 37627 13931 37661 13936
rect 35575 13835 35591 13869
rect 35591 13835 35609 13869
rect 35647 13835 35659 13869
rect 35659 13835 35681 13869
rect 35719 13835 35727 13869
rect 35727 13835 35753 13869
rect 35791 13835 35795 13869
rect 35795 13835 35825 13869
rect 35863 13835 35897 13869
rect 35935 13835 35965 13869
rect 35965 13835 35969 13869
rect 36007 13835 36033 13869
rect 36033 13835 36041 13869
rect 36079 13835 36101 13869
rect 36101 13835 36113 13869
rect 36151 13835 36169 13869
rect 36169 13835 36185 13869
rect 36223 13835 36237 13869
rect 36237 13835 36257 13869
rect 36295 13835 36305 13869
rect 36305 13835 36329 13869
rect 36367 13835 36373 13869
rect 36373 13835 36401 13869
rect 36439 13835 36441 13869
rect 36441 13835 36473 13869
rect 36511 13835 36543 13869
rect 36543 13835 36545 13869
rect 36583 13835 36611 13869
rect 36611 13835 36617 13869
rect 36655 13835 36679 13869
rect 36679 13835 36689 13869
rect 36727 13835 36747 13869
rect 36747 13835 36761 13869
rect 36799 13835 36815 13869
rect 36815 13835 36833 13869
rect 36871 13835 36883 13869
rect 36883 13835 36905 13869
rect 36943 13835 36951 13869
rect 36951 13835 36977 13869
rect 37015 13835 37019 13869
rect 37019 13835 37049 13869
rect 37087 13835 37121 13869
rect 37159 13835 37189 13869
rect 37189 13835 37193 13869
rect 37231 13835 37257 13869
rect 37257 13835 37265 13869
rect 37303 13835 37325 13869
rect 37325 13835 37337 13869
rect 37375 13835 37393 13869
rect 37393 13835 37409 13869
rect 37447 13835 37461 13869
rect 37461 13835 37481 13869
rect 37519 13835 37529 13869
rect 37529 13835 37553 13869
rect 37627 13866 37661 13892
rect 37627 13858 37661 13866
rect 37627 13796 37661 13819
rect 37627 13785 37661 13796
rect 37627 13726 37661 13746
rect 35575 13679 35591 13713
rect 35591 13679 35609 13713
rect 35647 13679 35659 13713
rect 35659 13679 35681 13713
rect 35719 13679 35727 13713
rect 35727 13679 35753 13713
rect 35791 13679 35795 13713
rect 35795 13679 35825 13713
rect 35863 13679 35897 13713
rect 35935 13679 35965 13713
rect 35965 13679 35969 13713
rect 36007 13679 36033 13713
rect 36033 13679 36041 13713
rect 36079 13679 36101 13713
rect 36101 13679 36113 13713
rect 36151 13679 36169 13713
rect 36169 13679 36185 13713
rect 36223 13679 36237 13713
rect 36237 13679 36257 13713
rect 36295 13679 36305 13713
rect 36305 13679 36329 13713
rect 36367 13679 36373 13713
rect 36373 13679 36401 13713
rect 36439 13679 36441 13713
rect 36441 13679 36473 13713
rect 36511 13679 36543 13713
rect 36543 13679 36545 13713
rect 36583 13679 36611 13713
rect 36611 13679 36617 13713
rect 36655 13679 36679 13713
rect 36679 13679 36689 13713
rect 36727 13679 36747 13713
rect 36747 13679 36761 13713
rect 36799 13679 36815 13713
rect 36815 13679 36833 13713
rect 36871 13679 36883 13713
rect 36883 13679 36905 13713
rect 36943 13679 36951 13713
rect 36951 13679 36977 13713
rect 37015 13679 37019 13713
rect 37019 13679 37049 13713
rect 37087 13679 37121 13713
rect 37159 13679 37189 13713
rect 37189 13679 37193 13713
rect 37231 13679 37257 13713
rect 37257 13679 37265 13713
rect 37303 13679 37325 13713
rect 37325 13679 37337 13713
rect 37375 13679 37393 13713
rect 37393 13679 37409 13713
rect 37447 13679 37461 13713
rect 37461 13679 37481 13713
rect 37519 13679 37529 13713
rect 37529 13679 37553 13713
rect 37627 13712 37661 13726
rect 37627 13656 37661 13672
rect 37627 13638 37661 13656
rect 37627 13586 37661 13598
rect 37627 13564 37661 13586
rect 35575 13523 35591 13557
rect 35591 13523 35609 13557
rect 35647 13523 35659 13557
rect 35659 13523 35681 13557
rect 35719 13523 35727 13557
rect 35727 13523 35753 13557
rect 35791 13523 35795 13557
rect 35795 13523 35825 13557
rect 35863 13523 35897 13557
rect 35935 13523 35965 13557
rect 35965 13523 35969 13557
rect 36007 13523 36033 13557
rect 36033 13523 36041 13557
rect 36079 13523 36101 13557
rect 36101 13523 36113 13557
rect 36151 13523 36169 13557
rect 36169 13523 36185 13557
rect 36223 13523 36237 13557
rect 36237 13523 36257 13557
rect 36295 13523 36305 13557
rect 36305 13523 36329 13557
rect 36367 13523 36373 13557
rect 36373 13523 36401 13557
rect 36439 13523 36441 13557
rect 36441 13523 36473 13557
rect 36511 13523 36543 13557
rect 36543 13523 36545 13557
rect 36583 13523 36611 13557
rect 36611 13523 36617 13557
rect 36655 13523 36679 13557
rect 36679 13523 36689 13557
rect 36727 13523 36747 13557
rect 36747 13523 36761 13557
rect 36799 13523 36815 13557
rect 36815 13523 36833 13557
rect 36871 13523 36883 13557
rect 36883 13523 36905 13557
rect 36943 13523 36951 13557
rect 36951 13523 36977 13557
rect 37015 13523 37019 13557
rect 37019 13523 37049 13557
rect 37087 13523 37121 13557
rect 37159 13523 37189 13557
rect 37189 13523 37193 13557
rect 37231 13523 37257 13557
rect 37257 13523 37265 13557
rect 37303 13523 37325 13557
rect 37325 13523 37337 13557
rect 37375 13523 37393 13557
rect 37393 13523 37409 13557
rect 37447 13523 37461 13557
rect 37461 13523 37481 13557
rect 37519 13523 37529 13557
rect 37529 13523 37553 13557
rect 37627 13516 37661 13524
rect 37627 13490 37661 13516
rect 37627 13446 37661 13450
rect 37627 13416 37661 13446
rect 35575 13367 35591 13401
rect 35591 13367 35609 13401
rect 35647 13367 35659 13401
rect 35659 13367 35681 13401
rect 35719 13367 35727 13401
rect 35727 13367 35753 13401
rect 35791 13367 35795 13401
rect 35795 13367 35825 13401
rect 35863 13367 35897 13401
rect 35935 13367 35965 13401
rect 35965 13367 35969 13401
rect 36007 13367 36033 13401
rect 36033 13367 36041 13401
rect 36079 13367 36101 13401
rect 36101 13367 36113 13401
rect 36151 13367 36169 13401
rect 36169 13367 36185 13401
rect 36223 13367 36237 13401
rect 36237 13367 36257 13401
rect 36295 13367 36305 13401
rect 36305 13367 36329 13401
rect 36367 13367 36373 13401
rect 36373 13367 36401 13401
rect 36439 13367 36441 13401
rect 36441 13367 36473 13401
rect 36511 13367 36543 13401
rect 36543 13367 36545 13401
rect 36583 13367 36611 13401
rect 36611 13367 36617 13401
rect 36655 13367 36679 13401
rect 36679 13367 36689 13401
rect 36727 13367 36747 13401
rect 36747 13367 36761 13401
rect 36799 13367 36815 13401
rect 36815 13367 36833 13401
rect 36871 13367 36883 13401
rect 36883 13367 36905 13401
rect 36943 13367 36951 13401
rect 36951 13367 36977 13401
rect 37015 13367 37019 13401
rect 37019 13367 37049 13401
rect 37087 13367 37121 13401
rect 37159 13367 37189 13401
rect 37189 13367 37193 13401
rect 37231 13367 37257 13401
rect 37257 13367 37265 13401
rect 37303 13367 37325 13401
rect 37325 13367 37337 13401
rect 37375 13367 37393 13401
rect 37393 13367 37409 13401
rect 37447 13367 37461 13401
rect 37461 13367 37481 13401
rect 37519 13367 37529 13401
rect 37529 13367 37553 13401
rect 37627 13342 37661 13376
rect 37627 13272 37661 13302
rect 37627 13268 37661 13272
rect 35575 13211 35591 13245
rect 35591 13211 35609 13245
rect 35647 13211 35659 13245
rect 35659 13211 35681 13245
rect 35719 13211 35727 13245
rect 35727 13211 35753 13245
rect 35791 13211 35795 13245
rect 35795 13211 35825 13245
rect 35863 13211 35897 13245
rect 35935 13211 35965 13245
rect 35965 13211 35969 13245
rect 36007 13211 36033 13245
rect 36033 13211 36041 13245
rect 36079 13211 36101 13245
rect 36101 13211 36113 13245
rect 36151 13211 36169 13245
rect 36169 13211 36185 13245
rect 36223 13211 36237 13245
rect 36237 13211 36257 13245
rect 36295 13211 36305 13245
rect 36305 13211 36329 13245
rect 36367 13211 36373 13245
rect 36373 13211 36401 13245
rect 36439 13211 36441 13245
rect 36441 13211 36473 13245
rect 36511 13211 36543 13245
rect 36543 13211 36545 13245
rect 36583 13211 36611 13245
rect 36611 13211 36617 13245
rect 36655 13211 36679 13245
rect 36679 13211 36689 13245
rect 36727 13211 36747 13245
rect 36747 13211 36761 13245
rect 36799 13211 36815 13245
rect 36815 13211 36833 13245
rect 36871 13211 36883 13245
rect 36883 13211 36905 13245
rect 36943 13211 36951 13245
rect 36951 13211 36977 13245
rect 37015 13211 37019 13245
rect 37019 13211 37049 13245
rect 37087 13211 37121 13245
rect 37159 13211 37189 13245
rect 37189 13211 37193 13245
rect 37231 13211 37257 13245
rect 37257 13211 37265 13245
rect 37303 13211 37325 13245
rect 37325 13211 37337 13245
rect 37375 13211 37393 13245
rect 37393 13211 37409 13245
rect 37447 13211 37461 13245
rect 37461 13211 37481 13245
rect 37519 13211 37529 13245
rect 37529 13211 37553 13245
rect 11752 3640 11779 3674
rect 11779 3640 11786 3674
rect 11826 3640 11849 3674
rect 11849 3640 11860 3674
rect 11900 3640 11919 3674
rect 11919 3640 11934 3674
rect 11974 3640 11989 3674
rect 11989 3640 12008 3674
rect 12048 3640 12059 3674
rect 12059 3640 12082 3674
rect 12122 3640 12129 3674
rect 12129 3640 12156 3674
rect 12196 3640 12199 3674
rect 12199 3640 12230 3674
rect 12270 3640 12304 3674
rect 12344 3640 12375 3674
rect 12375 3640 12378 3674
rect 12418 3640 12445 3674
rect 12445 3640 12452 3674
rect 12492 3640 12515 3674
rect 12515 3640 12526 3674
rect 12566 3640 12585 3674
rect 12585 3640 12600 3674
rect 12640 3640 12655 3674
rect 12655 3640 12674 3674
rect 12714 3640 12725 3674
rect 12725 3640 12748 3674
rect 12788 3640 12795 3674
rect 12795 3640 12822 3674
rect 12862 3640 12864 3674
rect 12864 3640 12896 3674
rect 12936 3640 12967 3674
rect 12967 3640 12970 3674
rect 13010 3640 13036 3674
rect 13036 3640 13044 3674
rect 13084 3640 13105 3674
rect 13105 3640 13118 3674
rect 13158 3640 13174 3674
rect 13174 3640 13192 3674
rect 13232 3640 13243 3674
rect 13243 3640 13266 3674
rect 13306 3640 13312 3674
rect 13312 3640 13340 3674
rect 13380 3640 13381 3674
rect 13381 3640 13414 3674
rect 13454 3640 13485 3674
rect 13485 3640 13488 3674
rect 13528 3640 13554 3674
rect 13554 3640 13562 3674
rect 13602 3640 13623 3674
rect 13623 3640 13636 3674
rect 13676 3640 13692 3674
rect 13692 3640 13710 3674
rect 13750 3640 13761 3674
rect 13761 3640 13784 3674
rect 13824 3640 13830 3674
rect 13830 3640 13858 3674
rect 13898 3640 13899 3674
rect 13899 3640 13932 3674
rect 13971 3640 14002 3674
rect 14002 3640 14005 3674
rect 14044 3640 14071 3674
rect 14071 3640 14078 3674
rect 14117 3640 14140 3674
rect 14140 3640 14151 3674
rect 14190 3640 14209 3674
rect 14209 3640 14224 3674
rect 14263 3640 14278 3674
rect 14278 3640 14297 3674
rect 14336 3640 14347 3674
rect 14347 3640 14370 3674
rect 14409 3640 14416 3674
rect 14416 3640 14443 3674
rect 14482 3640 14485 3674
rect 14485 3640 14516 3674
rect 14555 3640 14589 3674
rect 11749 3554 11783 3567
rect 11749 3533 11783 3554
rect 11749 3486 11783 3494
rect 11749 3460 11783 3486
rect 11749 3418 11783 3422
rect 11749 3388 11783 3418
rect 11749 3316 11783 3350
rect 11749 3248 11783 3278
rect 11749 3244 11783 3248
rect 11905 3554 11939 3567
rect 11905 3533 11939 3554
rect 11905 3452 11939 3479
rect 11905 3445 11939 3452
rect 11905 3384 11939 3391
rect 11905 3357 11939 3384
rect 11905 3282 11939 3303
rect 11905 3269 11939 3282
rect 11905 3214 11939 3215
rect 11905 3181 11939 3214
rect 12061 3554 12095 3567
rect 12061 3533 12095 3554
rect 12061 3452 12095 3479
rect 12061 3445 12095 3452
rect 12061 3384 12095 3391
rect 12061 3357 12095 3384
rect 12061 3282 12095 3303
rect 12061 3269 12095 3282
rect 12061 3214 12095 3215
rect 12061 3181 12095 3214
rect 12217 3384 12251 3391
rect 12217 3357 12251 3384
rect 12217 3282 12251 3313
rect 12217 3279 12251 3282
rect 12217 3214 12251 3235
rect 12217 3201 12251 3214
rect 12217 3146 12251 3157
rect 12217 3123 12251 3146
rect 12373 3554 12407 3567
rect 12373 3533 12407 3554
rect 12373 3452 12407 3484
rect 12373 3450 12407 3452
rect 12373 3384 12407 3402
rect 12373 3368 12407 3384
rect 12373 3316 12407 3320
rect 12373 3286 12407 3316
rect 12529 3554 12563 3567
rect 12529 3533 12563 3554
rect 12529 3452 12563 3484
rect 12529 3450 12563 3452
rect 12529 3384 12563 3402
rect 12529 3368 12563 3384
rect 12529 3316 12563 3320
rect 12529 3286 12563 3316
rect 12685 3554 12719 3567
rect 12685 3533 12719 3554
rect 12685 3452 12719 3484
rect 12685 3450 12719 3452
rect 12685 3384 12719 3402
rect 12685 3368 12719 3384
rect 12685 3316 12719 3320
rect 12685 3286 12719 3316
rect 12997 3554 13031 3567
rect 12997 3533 13031 3554
rect 12997 3486 13031 3491
rect 12997 3457 13031 3486
rect 12997 3384 13031 3416
rect 12997 3382 13031 3384
rect 12997 3316 13031 3341
rect 12997 3307 13031 3316
rect 12819 3180 12841 3211
rect 12841 3180 12853 3211
rect 12819 3177 12853 3180
rect 12891 3177 12925 3211
rect 13075 3220 13109 3254
rect 13075 3148 13109 3182
rect 11838 2884 11844 2918
rect 11844 2884 11872 2918
rect 11924 2884 11954 2918
rect 11954 2884 11958 2918
rect 12010 2884 12026 2918
rect 12026 2884 12044 2918
rect 12096 2884 12098 2918
rect 12098 2884 12130 2918
rect 12182 2884 12203 2918
rect 12203 2884 12216 2918
rect 12267 2884 12274 2918
rect 12274 2884 12301 2918
rect 12476 2884 12505 2918
rect 12505 2884 12510 2918
rect 12559 2884 12576 2918
rect 12576 2884 12593 2918
rect 12642 2884 12648 2918
rect 12648 2884 12676 2918
rect 12725 2884 12754 2918
rect 12754 2884 12759 2918
rect 12808 2884 12826 2918
rect 12826 2884 12842 2918
rect 12891 2884 12898 2918
rect 12898 2884 12925 2918
rect 13544 3220 13578 3254
rect 13544 3148 13578 3182
rect 13277 2968 13311 3002
rect 13349 2968 13383 3002
rect 13217 2884 13249 2918
rect 13249 2884 13251 2918
rect 13311 2884 13343 2918
rect 13343 2884 13345 2918
rect 13405 2884 13438 2918
rect 13438 2884 13439 2918
rect 13625 3146 13659 3154
rect 13625 3120 13655 3146
rect 13655 3120 13659 3146
rect 13625 3078 13659 3082
rect 13625 3048 13655 3078
rect 13655 3048 13659 3078
rect 13742 3146 13776 3156
rect 13742 3122 13776 3146
rect 13918 3350 13952 3381
rect 13918 3347 13952 3350
rect 13918 3282 13952 3299
rect 13918 3265 13952 3282
rect 14013 3282 14047 3312
rect 14013 3278 14042 3282
rect 14042 3278 14047 3282
rect 14085 3278 14119 3312
rect 14218 3214 14252 3227
rect 14218 3193 14252 3214
rect 14218 3146 14252 3154
rect 14218 3120 14252 3146
rect 14218 3078 14252 3082
rect 14218 3048 14252 3078
rect 13742 2981 13776 3015
rect 14407 2960 14441 2994
rect 14479 2960 14513 2994
rect 13636 2885 13670 2919
rect 13708 2885 13742 2919
rect 12317 2709 12351 2743
rect 12423 2709 12457 2743
rect 12528 2709 12562 2743
rect 13636 2709 13670 2743
rect 13708 2709 13742 2743
rect 12131 2562 12165 2596
rect 12224 2562 12258 2596
rect 12131 2480 12165 2514
rect 12224 2480 12258 2514
rect 12001 2203 12035 2237
rect 12001 2126 12035 2160
rect 12001 2049 12035 2083
rect 12981 2627 13015 2661
rect 12583 2566 12614 2596
rect 12614 2566 12617 2596
rect 12656 2566 12684 2596
rect 12684 2566 12690 2596
rect 12729 2566 12753 2596
rect 12753 2566 12763 2596
rect 12801 2566 12822 2596
rect 12822 2566 12835 2596
rect 14095 2901 14129 2919
rect 14095 2885 14122 2901
rect 14122 2885 14129 2901
rect 14167 2885 14201 2919
rect 14275 2867 14299 2883
rect 14299 2867 14309 2883
rect 14275 2849 14309 2867
rect 14347 2849 14381 2883
rect 13820 2633 13854 2667
rect 13894 2633 13928 2667
rect 13967 2633 14001 2667
rect 14553 2662 14587 2696
rect 14625 2662 14659 2696
rect 18459 2623 18493 2657
rect 18536 2623 18570 2657
rect 18613 2623 18647 2657
rect 18689 2623 18723 2657
rect 18765 2623 18799 2657
rect 18841 2623 18875 2657
rect 18917 2623 18951 2657
rect 18993 2623 19027 2657
rect 19069 2623 19103 2657
rect 19145 2623 19179 2657
rect 19221 2623 19255 2657
rect 19297 2623 19331 2657
rect 19373 2623 19407 2657
rect 19449 2623 19483 2657
rect 19525 2623 19559 2657
rect 19601 2623 19635 2657
rect 19677 2623 19711 2657
rect 12583 2562 12617 2566
rect 12656 2562 12690 2566
rect 12729 2562 12763 2566
rect 12801 2562 12835 2566
rect 12583 2480 12617 2514
rect 12656 2480 12690 2514
rect 12729 2480 12763 2514
rect 12801 2480 12835 2514
rect 12981 2534 13015 2568
rect 13551 2513 13585 2522
rect 12981 2441 13015 2475
rect 12981 2348 13015 2382
rect 12761 2289 12774 2302
rect 12774 2289 12795 2302
rect 12833 2289 12842 2302
rect 12842 2289 12867 2302
rect 12761 2268 12795 2289
rect 12833 2268 12867 2289
rect 12645 2090 12679 2124
rect 12717 2090 12751 2124
rect 12962 2036 12996 2070
rect 13034 2036 13068 2070
rect 12495 1894 12497 1917
rect 12497 1894 12529 1917
rect 12495 1883 12529 1894
rect 13254 2188 13288 2222
rect 13254 2116 13288 2150
rect 13334 2423 13368 2457
rect 13334 2353 13368 2385
rect 13334 2351 13368 2353
rect 13178 1979 13212 1987
rect 13178 1953 13212 1979
rect 13178 1911 13212 1913
rect 13178 1879 13212 1911
rect 12495 1811 12529 1845
rect 13178 1806 13212 1840
rect 13551 2488 13585 2513
rect 13638 2513 13672 2522
rect 13725 2513 13759 2522
rect 13860 2513 13894 2516
rect 13942 2513 13976 2516
rect 14024 2513 14058 2516
rect 14106 2513 14140 2516
rect 13638 2488 13646 2513
rect 13646 2488 13672 2513
rect 13725 2488 13741 2513
rect 13741 2488 13759 2513
rect 13860 2482 13863 2513
rect 13863 2482 13894 2513
rect 13942 2482 13969 2513
rect 13969 2482 13976 2513
rect 14024 2482 14041 2513
rect 14041 2482 14058 2513
rect 14106 2482 14113 2513
rect 14113 2482 14140 2513
rect 14189 2482 14223 2516
rect 14272 2513 14306 2516
rect 14355 2513 14389 2516
rect 14505 2513 14539 2514
rect 14586 2513 14620 2514
rect 14272 2482 14294 2513
rect 14294 2482 14306 2513
rect 14355 2482 14365 2513
rect 14365 2482 14389 2513
rect 14505 2480 14521 2513
rect 14521 2480 14539 2513
rect 14586 2480 14592 2513
rect 14592 2480 14620 2513
rect 14667 2480 14701 2514
rect 14748 2513 14782 2514
rect 14829 2513 14863 2514
rect 14910 2513 14944 2514
rect 14992 2513 15026 2514
rect 14748 2480 14773 2513
rect 14773 2480 14782 2513
rect 14829 2480 14845 2513
rect 14845 2480 14863 2513
rect 14910 2480 14917 2513
rect 14917 2480 14944 2513
rect 14992 2480 15023 2513
rect 15023 2480 15026 2513
rect 15350 2493 15384 2527
rect 13412 2188 13446 2222
rect 13412 2116 13446 2150
rect 13567 2113 13601 2147
rect 13567 2041 13601 2075
rect 13646 2285 13680 2296
rect 13646 2262 13680 2285
rect 13646 2217 13680 2224
rect 13646 2190 13680 2217
rect 13490 1979 13524 1987
rect 13490 1953 13524 1979
rect 13490 1911 13524 1913
rect 13490 1879 13524 1911
rect 13490 1806 13524 1840
rect 15350 2421 15384 2455
rect 13727 2113 13761 2147
rect 13727 2041 13761 2075
rect 13802 2081 13836 2100
rect 13802 2066 13836 2081
rect 13802 1979 13836 2013
rect 13802 1911 13836 1926
rect 13802 1892 13836 1911
rect 13802 1806 13836 1840
rect 13959 2355 13993 2389
rect 13959 2285 13993 2313
rect 13959 2279 13992 2285
rect 13992 2279 13993 2285
rect 13959 2217 13993 2237
rect 13959 2203 13992 2217
rect 13992 2203 13993 2217
rect 14114 2047 14148 2056
rect 14114 2022 14148 2047
rect 14114 1979 14148 1984
rect 14114 1950 14148 1979
rect 14114 1911 14148 1912
rect 14114 1878 14148 1911
rect 14114 1806 14148 1840
rect 14270 2355 14304 2389
rect 14270 2285 14304 2313
rect 14270 2279 14304 2285
rect 14270 2217 14304 2237
rect 14270 2203 14304 2217
rect 14426 2047 14460 2056
rect 14426 2022 14460 2047
rect 14426 1979 14460 1984
rect 14426 1950 14460 1979
rect 14426 1911 14460 1912
rect 14426 1878 14460 1911
rect 14426 1806 14460 1840
rect 14583 2355 14617 2389
rect 14583 2285 14617 2313
rect 14583 2279 14616 2285
rect 14616 2279 14617 2285
rect 14583 2217 14617 2237
rect 14583 2203 14616 2217
rect 14616 2203 14617 2217
rect 14738 2047 14772 2056
rect 14738 2022 14772 2047
rect 14738 1979 14772 1984
rect 14738 1950 14772 1979
rect 14738 1911 14772 1912
rect 14738 1878 14772 1911
rect 14738 1806 14772 1840
rect 14894 2355 14928 2389
rect 14894 2285 14928 2313
rect 14894 2279 14928 2285
rect 14894 2217 14928 2237
rect 14894 2203 14928 2217
rect 15457 2492 15491 2526
rect 15457 2420 15491 2454
rect 16410 2493 16444 2527
rect 16410 2421 16444 2455
rect 17617 2439 17651 2473
rect 17689 2439 17723 2473
rect 16622 2333 16656 2367
rect 16694 2333 16728 2367
rect 18442 2260 18476 2294
rect 18515 2260 18549 2294
rect 18588 2260 18622 2294
rect 18661 2260 18695 2294
rect 18734 2260 18768 2294
rect 18807 2260 18841 2294
rect 18880 2260 18914 2294
rect 18953 2260 18987 2294
rect 19026 2260 19060 2294
rect 19099 2260 19133 2294
rect 19172 2260 19206 2294
rect 19245 2260 19279 2294
rect 19318 2260 19352 2294
rect 19391 2260 19425 2294
rect 19464 2260 19498 2294
rect 19537 2260 19571 2294
rect 19610 2260 19644 2294
rect 19682 2260 19716 2294
rect 19754 2260 19788 2294
rect 16206 2196 16240 2230
rect 16278 2196 16312 2230
rect 16798 2182 16832 2216
rect 16870 2182 16904 2216
rect 15893 2109 15927 2143
rect 15966 2109 16000 2143
rect 16212 2109 16246 2143
rect 16285 2109 16319 2143
rect 20434 2114 20468 2148
rect 20507 2114 20541 2148
rect 20580 2114 20614 2148
rect 20653 2114 20687 2148
rect 20726 2114 20760 2148
rect 20799 2114 20833 2148
rect 20872 2114 20906 2148
rect 20945 2114 20979 2148
rect 21018 2114 21052 2148
rect 21091 2114 21125 2148
rect 21164 2114 21198 2148
rect 21237 2114 21271 2148
rect 21310 2114 21344 2148
rect 21383 2114 21417 2148
rect 21456 2114 21490 2148
rect 21529 2114 21563 2148
rect 21602 2114 21636 2148
rect 21675 2114 21709 2148
rect 21748 2114 21782 2148
rect 21821 2114 21855 2148
rect 21894 2114 21928 2148
rect 21967 2114 22001 2148
rect 22040 2114 22074 2148
rect 22113 2114 22147 2148
rect 22185 2114 22219 2148
rect 22257 2114 22291 2148
rect 22329 2114 22363 2148
rect 22401 2114 22435 2148
rect 22473 2114 22507 2148
rect 22545 2114 22579 2148
rect 22617 2114 22651 2148
rect 22689 2114 22723 2148
rect 22761 2114 22795 2148
rect 22833 2114 22867 2148
rect 22905 2114 22939 2148
rect 22977 2114 23011 2148
rect 23049 2114 23083 2148
rect 23121 2114 23155 2148
rect 23193 2114 23227 2148
rect 23265 2114 23299 2148
rect 23337 2114 23371 2148
rect 23409 2114 23443 2148
rect 23481 2114 23515 2148
rect 23553 2114 23587 2148
rect 15050 2047 15084 2056
rect 15050 2022 15084 2047
rect 16064 2033 16098 2067
rect 16137 2033 16171 2067
rect 15050 1979 15084 1984
rect 15050 1950 15084 1979
rect 15050 1911 15084 1912
rect 15050 1878 15084 1911
rect 15050 1806 15084 1840
rect 15370 1959 15404 1993
rect 15465 1959 15499 1993
rect 15559 1959 15593 1993
rect 16411 1953 16445 1987
rect 18459 1941 18493 1975
rect 18537 1941 18571 1975
rect 18615 1941 18649 1975
rect 18693 1941 18727 1975
rect 18771 1941 18805 1975
rect 18848 1941 18882 1975
rect 18925 1941 18959 1975
rect 19002 1941 19036 1975
rect 19079 1941 19113 1975
rect 19156 1941 19190 1975
rect 19233 1941 19267 1975
rect 19310 1941 19344 1975
rect 16411 1881 16445 1915
rect 15370 1839 15404 1873
rect 15465 1839 15499 1873
rect 15559 1839 15593 1873
rect 12141 1723 12156 1757
rect 12156 1723 12175 1757
rect 12214 1723 12225 1757
rect 12225 1723 12248 1757
rect 12287 1723 12294 1757
rect 12294 1723 12321 1757
rect 12360 1723 12363 1757
rect 12363 1723 12394 1757
rect 12433 1723 12466 1757
rect 12466 1723 12467 1757
rect 12506 1723 12535 1757
rect 12535 1723 12540 1757
rect 12579 1723 12604 1757
rect 12604 1723 12613 1757
rect 12652 1723 12673 1757
rect 12673 1723 12686 1757
rect 12725 1723 12742 1757
rect 12742 1723 12759 1757
rect 12798 1723 12811 1757
rect 12811 1723 12832 1757
rect 12871 1723 12880 1757
rect 12880 1723 12905 1757
rect 12944 1723 12949 1757
rect 12949 1723 12978 1757
rect 13017 1723 13018 1757
rect 13018 1723 13051 1757
rect 13090 1723 13122 1757
rect 13122 1723 13124 1757
rect 13163 1723 13191 1757
rect 13191 1723 13197 1757
rect 13236 1723 13260 1757
rect 13260 1723 13270 1757
rect 13309 1723 13329 1757
rect 13329 1723 13343 1757
rect 13382 1723 13398 1757
rect 13398 1723 13416 1757
rect 13455 1723 13467 1757
rect 13467 1723 13489 1757
rect 13528 1723 13536 1757
rect 13536 1723 13562 1757
rect 13601 1723 13605 1757
rect 13605 1723 13635 1757
rect 13674 1723 13708 1757
rect 13747 1723 13777 1757
rect 13777 1723 13781 1757
rect 13820 1723 13846 1757
rect 13846 1723 13854 1757
rect 13893 1723 13915 1757
rect 13915 1723 13927 1757
rect 13966 1723 13984 1757
rect 13984 1723 14000 1757
rect 14039 1723 14053 1757
rect 14053 1723 14073 1757
rect 14112 1723 14122 1757
rect 14122 1723 14146 1757
rect 14185 1723 14191 1757
rect 14191 1723 14219 1757
rect 14258 1723 14260 1757
rect 14260 1723 14292 1757
rect 14331 1723 14364 1757
rect 14364 1723 14365 1757
rect 14404 1723 14433 1757
rect 14433 1723 14438 1757
rect 14477 1723 14502 1757
rect 14502 1723 14511 1757
rect 14550 1723 14571 1757
rect 14571 1723 14584 1757
rect 14623 1723 14640 1757
rect 14640 1723 14657 1757
rect 14696 1723 14709 1757
rect 14709 1723 14730 1757
rect 14769 1723 14778 1757
rect 14778 1723 14803 1757
rect 14842 1723 14847 1757
rect 14847 1723 14876 1757
rect 14915 1723 14916 1757
rect 14916 1723 14949 1757
rect 14988 1723 15019 1757
rect 15019 1723 15022 1757
rect 15061 1723 15088 1757
rect 15088 1723 15095 1757
rect 15134 1723 15157 1757
rect 15157 1723 15168 1757
rect 15207 1723 15226 1757
rect 15226 1723 15241 1757
rect 15280 1723 15295 1757
rect 15295 1723 15314 1757
rect 15353 1723 15363 1757
rect 15363 1723 15387 1757
rect 15426 1723 15431 1757
rect 15431 1723 15460 1757
rect 15498 1723 15499 1757
rect 15499 1723 15532 1757
rect 15570 1723 15601 1757
rect 15601 1723 15604 1757
rect 15642 1723 15669 1757
rect 15669 1723 15676 1757
rect 15714 1723 15737 1757
rect 15737 1723 15748 1757
rect 15786 1723 15820 1757
rect 20977 1691 21011 1692
rect 21051 1691 21085 1692
rect 21125 1691 21159 1692
rect 21199 1691 21233 1692
rect 21273 1691 21307 1692
rect 21347 1691 21381 1692
rect 21421 1691 21455 1692
rect 21495 1691 21529 1692
rect 21569 1691 21603 1692
rect 21643 1691 21677 1692
rect 21717 1691 21751 1692
rect 21791 1691 21825 1692
rect 21865 1691 21899 1692
rect 21939 1691 21973 1692
rect 22013 1691 22047 1692
rect 22087 1691 22121 1692
rect 22161 1691 22195 1692
rect 22235 1691 22269 1692
rect 22309 1691 22343 1692
rect 22383 1691 22417 1692
rect 22457 1691 22491 1692
rect 22531 1691 22565 1692
rect 22605 1691 22639 1692
rect 22679 1691 22713 1692
rect 22753 1691 22787 1692
rect 22827 1691 22861 1692
rect 22901 1691 22935 1692
rect 22975 1691 23009 1692
rect 23049 1691 23083 1692
rect 23123 1691 23157 1692
rect 23196 1691 23230 1692
rect 23269 1691 23303 1692
rect 23342 1691 23376 1692
rect 23415 1691 23449 1692
rect 23488 1691 23522 1692
rect 23561 1691 23595 1692
rect 18160 1657 18163 1691
rect 18163 1657 18194 1691
rect 18232 1657 18266 1691
rect 18304 1657 18335 1691
rect 18335 1657 18338 1691
rect 18376 1657 18404 1691
rect 18404 1657 18410 1691
rect 18448 1657 18473 1691
rect 18473 1657 18482 1691
rect 18520 1657 18542 1691
rect 18542 1657 18554 1691
rect 18592 1657 18611 1691
rect 18611 1657 18626 1691
rect 18664 1657 18680 1691
rect 18680 1657 18698 1691
rect 18736 1657 18749 1691
rect 18749 1657 18770 1691
rect 18808 1657 18818 1691
rect 18818 1657 18842 1691
rect 18880 1657 18887 1691
rect 18887 1657 18914 1691
rect 18952 1657 18956 1691
rect 18956 1657 18986 1691
rect 19024 1657 19025 1691
rect 19025 1657 19058 1691
rect 19096 1657 19129 1691
rect 19129 1657 19130 1691
rect 19168 1657 19198 1691
rect 19198 1657 19202 1691
rect 19240 1657 19267 1691
rect 19267 1657 19274 1691
rect 19312 1657 19336 1691
rect 19336 1657 19346 1691
rect 19384 1657 19405 1691
rect 19405 1657 19418 1691
rect 19456 1657 19474 1691
rect 19474 1657 19490 1691
rect 19528 1657 19543 1691
rect 19543 1657 19562 1691
rect 19600 1657 19612 1691
rect 19612 1657 19634 1691
rect 19672 1657 19681 1691
rect 19681 1657 19706 1691
rect 19744 1657 19750 1691
rect 19750 1657 19778 1691
rect 19816 1657 19819 1691
rect 19819 1657 19850 1691
rect 19888 1657 19922 1691
rect 19960 1657 19991 1691
rect 19991 1657 19994 1691
rect 20032 1657 20060 1691
rect 20060 1657 20066 1691
rect 20104 1657 20129 1691
rect 20129 1657 20138 1691
rect 20176 1657 20198 1691
rect 20198 1657 20210 1691
rect 20248 1657 20267 1691
rect 20267 1657 20282 1691
rect 20320 1657 20336 1691
rect 20336 1657 20354 1691
rect 20392 1657 20405 1691
rect 20405 1657 20426 1691
rect 20464 1657 20474 1691
rect 20474 1657 20498 1691
rect 20536 1657 20543 1691
rect 20543 1657 20570 1691
rect 20608 1657 20612 1691
rect 20612 1657 20642 1691
rect 20680 1657 20681 1691
rect 20681 1657 20714 1691
rect 20977 1658 20992 1691
rect 20992 1658 21011 1691
rect 21051 1658 21061 1691
rect 21061 1658 21085 1691
rect 21125 1658 21130 1691
rect 21130 1658 21159 1691
rect 21199 1658 21233 1691
rect 21273 1658 21302 1691
rect 21302 1658 21307 1691
rect 21347 1658 21371 1691
rect 21371 1658 21381 1691
rect 21421 1658 21440 1691
rect 21440 1658 21455 1691
rect 21495 1658 21509 1691
rect 21509 1658 21529 1691
rect 21569 1658 21577 1691
rect 21577 1658 21603 1691
rect 21643 1658 21645 1691
rect 21645 1658 21677 1691
rect 21717 1658 21747 1691
rect 21747 1658 21751 1691
rect 21791 1658 21815 1691
rect 21815 1658 21825 1691
rect 21865 1658 21883 1691
rect 21883 1658 21899 1691
rect 21939 1658 21951 1691
rect 21951 1658 21973 1691
rect 22013 1658 22019 1691
rect 22019 1658 22047 1691
rect 22087 1658 22121 1691
rect 22161 1658 22189 1691
rect 22189 1658 22195 1691
rect 22235 1658 22257 1691
rect 22257 1658 22269 1691
rect 22309 1658 22325 1691
rect 22325 1658 22343 1691
rect 22383 1658 22393 1691
rect 22393 1658 22417 1691
rect 22457 1658 22461 1691
rect 22461 1658 22491 1691
rect 22531 1658 22563 1691
rect 22563 1658 22565 1691
rect 22605 1658 22631 1691
rect 22631 1658 22639 1691
rect 22679 1658 22699 1691
rect 22699 1658 22713 1691
rect 22753 1658 22767 1691
rect 22767 1658 22787 1691
rect 22827 1658 22835 1691
rect 22835 1658 22861 1691
rect 22901 1658 22903 1691
rect 22903 1658 22935 1691
rect 22975 1658 23005 1691
rect 23005 1658 23009 1691
rect 23049 1658 23073 1691
rect 23073 1658 23083 1691
rect 23123 1658 23141 1691
rect 23141 1658 23157 1691
rect 23196 1658 23209 1691
rect 23209 1658 23230 1691
rect 23269 1658 23277 1691
rect 23277 1658 23303 1691
rect 23342 1658 23345 1691
rect 23345 1658 23376 1691
rect 23415 1658 23447 1691
rect 23447 1658 23449 1691
rect 23488 1658 23515 1691
rect 23515 1658 23522 1691
rect 23561 1658 23583 1691
rect 23583 1658 23595 1691
<< metal1 >>
rect 37686 16157 37770 16163
rect 37686 16105 37702 16157
rect 37754 16105 37770 16157
rect 37686 16093 37770 16105
rect 37686 16041 37702 16093
rect 37754 16041 37770 16093
rect 37686 16029 37770 16041
rect 37686 15977 37702 16029
rect 37754 15977 37770 16029
rect 37686 15971 37770 15977
tri 35666 15123 35669 15126 se
rect 35669 15123 35675 15126
rect 35563 15117 35675 15123
rect 35727 15117 35742 15126
rect 35794 15117 35809 15126
rect 35861 15117 35877 15126
rect 35929 15117 35945 15126
rect 35997 15117 36013 15126
rect 36065 15117 36081 15126
rect 35563 15083 35575 15117
rect 35609 15083 35647 15117
rect 35861 15083 35863 15117
rect 35929 15083 35935 15117
rect 35997 15083 36007 15117
rect 36065 15083 36079 15117
rect 35563 15077 35675 15083
tri 35666 15074 35669 15077 ne
rect 35669 15074 35675 15077
rect 35727 15074 35742 15083
rect 35794 15074 35809 15083
rect 35861 15074 35877 15083
rect 35929 15074 35945 15083
rect 35997 15074 36013 15083
rect 36065 15074 36081 15083
rect 36133 15074 36149 15126
rect 36201 15074 36217 15126
rect 36269 15074 36285 15126
rect 36337 15074 36353 15126
rect 36405 15074 36421 15126
rect 36473 15074 36489 15126
rect 36541 15123 36547 15126
tri 36547 15123 36550 15126 sw
rect 36541 15117 37565 15123
rect 36545 15083 36583 15117
rect 36617 15083 36655 15117
rect 36689 15083 36727 15117
rect 36761 15083 36799 15117
rect 36833 15083 36871 15117
rect 36905 15083 36943 15117
rect 36977 15083 37015 15117
rect 37049 15083 37087 15117
rect 37121 15083 37159 15117
rect 37193 15083 37231 15117
rect 37265 15083 37303 15117
rect 37337 15083 37375 15117
rect 37409 15083 37447 15117
rect 37481 15083 37519 15117
rect 37553 15083 37565 15117
rect 36541 15077 37565 15083
rect 36541 15074 36547 15077
tri 36547 15074 36550 15077 nw
rect 37618 15066 37670 15072
rect 37618 15002 37670 15014
tri 36658 14967 36661 14970 se
rect 36661 14967 36667 14970
rect 35563 14961 36667 14967
rect 36719 14961 36732 14970
rect 35563 14927 35575 14961
rect 35609 14927 35647 14961
rect 35681 14927 35719 14961
rect 35753 14927 35791 14961
rect 35825 14927 35863 14961
rect 35897 14927 35935 14961
rect 35969 14927 36007 14961
rect 36041 14927 36079 14961
rect 36113 14927 36151 14961
rect 36185 14927 36223 14961
rect 36257 14927 36295 14961
rect 36329 14927 36367 14961
rect 36401 14927 36439 14961
rect 36473 14927 36511 14961
rect 36545 14927 36583 14961
rect 36617 14927 36655 14961
rect 36719 14927 36727 14961
rect 35563 14921 36667 14927
tri 36658 14918 36661 14921 ne
rect 36661 14918 36667 14921
rect 36719 14918 36732 14927
rect 36784 14918 36797 14970
rect 36849 14918 36862 14970
rect 36914 14918 36927 14970
rect 36979 14918 36992 14970
rect 37044 14961 37057 14970
rect 37109 14961 37122 14970
rect 37174 14961 37188 14970
rect 37240 14961 37254 14970
rect 37306 14961 37320 14970
rect 37372 14961 37386 14970
rect 37438 14961 37452 14970
rect 37504 14967 37510 14970
tri 37510 14967 37513 14970 sw
rect 37504 14961 37565 14967
rect 37049 14927 37057 14961
rect 37121 14927 37122 14961
rect 37372 14927 37375 14961
rect 37438 14927 37447 14961
rect 37504 14927 37519 14961
rect 37553 14927 37565 14961
rect 37044 14918 37057 14927
rect 37109 14918 37122 14927
rect 37174 14918 37188 14927
rect 37240 14918 37254 14927
rect 37306 14918 37320 14927
rect 37372 14918 37386 14927
rect 37438 14918 37452 14927
rect 37504 14921 37565 14927
rect 37618 14938 37670 14950
rect 37504 14918 37510 14921
tri 37510 14918 37513 14921 nw
rect 37618 14880 37627 14886
rect 37661 14880 37670 14886
rect 37618 14874 37670 14880
tri 35666 14811 35669 14814 se
rect 35669 14811 35675 14814
rect 35563 14805 35675 14811
rect 35727 14805 35742 14814
rect 35794 14805 35809 14814
rect 35861 14805 35877 14814
rect 35929 14805 35945 14814
rect 35997 14805 36013 14814
rect 36065 14805 36081 14814
rect 35563 14771 35575 14805
rect 35609 14771 35647 14805
rect 35861 14771 35863 14805
rect 35929 14771 35935 14805
rect 35997 14771 36007 14805
rect 36065 14771 36079 14805
rect 35563 14765 35675 14771
tri 35666 14762 35669 14765 ne
rect 35669 14762 35675 14765
rect 35727 14762 35742 14771
rect 35794 14762 35809 14771
rect 35861 14762 35877 14771
rect 35929 14762 35945 14771
rect 35997 14762 36013 14771
rect 36065 14762 36081 14771
rect 36133 14762 36149 14814
rect 36201 14762 36217 14814
rect 36269 14762 36285 14814
rect 36337 14762 36353 14814
rect 36405 14762 36421 14814
rect 36473 14762 36489 14814
rect 36541 14811 36547 14814
tri 36547 14811 36550 14814 sw
rect 36541 14805 37565 14811
rect 36545 14771 36583 14805
rect 36617 14771 36655 14805
rect 36689 14771 36727 14805
rect 36761 14771 36799 14805
rect 36833 14771 36871 14805
rect 36905 14771 36943 14805
rect 36977 14771 37015 14805
rect 37049 14771 37087 14805
rect 37121 14771 37159 14805
rect 37193 14771 37231 14805
rect 37265 14771 37303 14805
rect 37337 14771 37375 14805
rect 37409 14771 37447 14805
rect 37481 14771 37519 14805
rect 37553 14771 37565 14805
rect 36541 14765 37565 14771
rect 37618 14809 37627 14822
rect 37661 14809 37670 14822
rect 36541 14762 36547 14765
tri 36547 14762 36550 14765 nw
rect 37618 14744 37627 14757
rect 37661 14744 37670 14757
rect 37618 14679 37627 14692
rect 37661 14679 37670 14692
tri 36658 14655 36661 14658 se
rect 36661 14655 36667 14658
rect 35563 14649 36667 14655
rect 36719 14649 36732 14658
rect 35563 14615 35575 14649
rect 35609 14615 35647 14649
rect 35681 14615 35719 14649
rect 35753 14615 35791 14649
rect 35825 14615 35863 14649
rect 35897 14615 35935 14649
rect 35969 14615 36007 14649
rect 36041 14615 36079 14649
rect 36113 14615 36151 14649
rect 36185 14615 36223 14649
rect 36257 14615 36295 14649
rect 36329 14615 36367 14649
rect 36401 14615 36439 14649
rect 36473 14615 36511 14649
rect 36545 14615 36583 14649
rect 36617 14615 36655 14649
rect 36719 14615 36727 14649
rect 35563 14609 36667 14615
tri 36658 14606 36661 14609 ne
rect 36661 14606 36667 14609
rect 36719 14606 36732 14615
rect 36784 14606 36797 14658
rect 36849 14606 36862 14658
rect 36914 14606 36927 14658
rect 36979 14606 36992 14658
rect 37044 14649 37057 14658
rect 37109 14649 37122 14658
rect 37174 14649 37188 14658
rect 37240 14649 37254 14658
rect 37306 14649 37320 14658
rect 37372 14649 37386 14658
rect 37438 14649 37452 14658
rect 37504 14655 37510 14658
tri 37510 14655 37513 14658 sw
rect 37504 14649 37565 14655
rect 37049 14615 37057 14649
rect 37121 14615 37122 14649
rect 37372 14615 37375 14649
rect 37438 14615 37447 14649
rect 37504 14615 37519 14649
rect 37553 14615 37565 14649
rect 37044 14606 37057 14615
rect 37109 14606 37122 14615
rect 37174 14606 37188 14615
rect 37240 14606 37254 14615
rect 37306 14606 37320 14615
rect 37372 14606 37386 14615
rect 37438 14606 37452 14615
rect 37504 14609 37565 14615
rect 37618 14622 37670 14627
rect 37618 14614 37627 14622
rect 37661 14614 37670 14622
rect 37504 14606 37510 14609
tri 37510 14606 37513 14609 nw
rect 37618 14549 37670 14562
tri 35666 14499 35669 14502 se
rect 35669 14499 35675 14502
rect 35563 14493 35675 14499
rect 35727 14493 35742 14502
rect 35794 14493 35809 14502
rect 35861 14493 35877 14502
rect 35929 14493 35945 14502
rect 35997 14493 36013 14502
rect 36065 14493 36081 14502
rect 35563 14459 35575 14493
rect 35609 14459 35647 14493
rect 35861 14459 35863 14493
rect 35929 14459 35935 14493
rect 35997 14459 36007 14493
rect 36065 14459 36079 14493
rect 35563 14453 35675 14459
tri 35666 14450 35669 14453 ne
rect 35669 14450 35675 14453
rect 35727 14450 35742 14459
rect 35794 14450 35809 14459
rect 35861 14450 35877 14459
rect 35929 14450 35945 14459
rect 35997 14450 36013 14459
rect 36065 14450 36081 14459
rect 36133 14450 36149 14502
rect 36201 14450 36217 14502
rect 36269 14450 36285 14502
rect 36337 14450 36353 14502
rect 36405 14450 36421 14502
rect 36473 14450 36489 14502
rect 36541 14499 36547 14502
tri 36547 14499 36550 14502 sw
rect 36541 14493 37565 14499
rect 36545 14459 36583 14493
rect 36617 14459 36655 14493
rect 36689 14459 36727 14493
rect 36761 14459 36799 14493
rect 36833 14459 36871 14493
rect 36905 14459 36943 14493
rect 36977 14459 37015 14493
rect 37049 14459 37087 14493
rect 37121 14459 37159 14493
rect 37193 14459 37231 14493
rect 37265 14459 37303 14493
rect 37337 14459 37375 14493
rect 37409 14459 37447 14493
rect 37481 14459 37519 14493
rect 37553 14459 37565 14493
rect 36541 14453 37565 14459
rect 37618 14484 37670 14497
rect 36541 14450 36547 14453
tri 36547 14450 36550 14453 nw
rect 37618 14419 37670 14432
rect 37618 14354 37670 14367
tri 36658 14343 36661 14346 se
rect 36661 14343 36667 14346
rect 35563 14337 36667 14343
rect 36719 14337 36732 14346
rect 35563 14303 35575 14337
rect 35609 14303 35647 14337
rect 35681 14303 35719 14337
rect 35753 14303 35791 14337
rect 35825 14303 35863 14337
rect 35897 14303 35935 14337
rect 35969 14303 36007 14337
rect 36041 14303 36079 14337
rect 36113 14303 36151 14337
rect 36185 14303 36223 14337
rect 36257 14303 36295 14337
rect 36329 14303 36367 14337
rect 36401 14303 36439 14337
rect 36473 14303 36511 14337
rect 36545 14303 36583 14337
rect 36617 14303 36655 14337
rect 36719 14303 36727 14337
rect 35563 14297 36667 14303
tri 36658 14296 36659 14297 ne
rect 36659 14296 36667 14297
tri 36659 14294 36661 14296 ne
rect 36661 14294 36667 14296
rect 36719 14294 36732 14303
rect 36784 14294 36797 14346
rect 36849 14294 36862 14346
rect 36914 14294 36927 14346
rect 36979 14294 36992 14346
rect 37044 14337 37057 14346
rect 37109 14337 37122 14346
rect 37174 14337 37188 14346
rect 37240 14337 37254 14346
rect 37306 14337 37320 14346
rect 37372 14337 37386 14346
rect 37438 14337 37452 14346
rect 37504 14343 37510 14346
tri 37510 14343 37513 14346 sw
rect 37504 14337 37565 14343
rect 37049 14303 37057 14337
rect 37121 14303 37122 14337
rect 37372 14303 37375 14337
rect 37438 14303 37447 14337
rect 37504 14303 37519 14337
rect 37553 14303 37565 14337
rect 37044 14294 37057 14303
rect 37109 14294 37122 14303
rect 37174 14294 37188 14303
rect 37240 14294 37254 14303
rect 37306 14294 37320 14303
rect 37372 14294 37386 14303
rect 37438 14294 37452 14303
rect 37504 14297 37565 14303
rect 37504 14296 37512 14297
tri 37512 14296 37513 14297 nw
rect 37618 14296 37627 14302
rect 37661 14296 37670 14302
rect 37504 14294 37510 14296
tri 37510 14294 37512 14296 nw
rect 37618 14289 37670 14296
rect 37618 14224 37627 14237
rect 37661 14224 37670 14237
tri 35666 14187 35669 14190 se
rect 35669 14187 35675 14190
rect 35563 14181 35675 14187
rect 35727 14181 35742 14190
rect 35794 14181 35809 14190
rect 35861 14181 35877 14190
rect 35929 14181 35945 14190
rect 35997 14181 36013 14190
rect 36065 14181 36081 14190
rect 35563 14147 35575 14181
rect 35609 14147 35647 14181
rect 35861 14147 35863 14181
rect 35929 14147 35935 14181
rect 35997 14147 36007 14181
rect 36065 14147 36079 14181
rect 35563 14141 35675 14147
tri 35666 14138 35669 14141 ne
rect 35669 14138 35675 14141
rect 35727 14138 35742 14147
rect 35794 14138 35809 14147
rect 35861 14138 35877 14147
rect 35929 14138 35945 14147
rect 35997 14138 36013 14147
rect 36065 14138 36081 14147
rect 36133 14138 36149 14190
rect 36201 14138 36217 14190
rect 36269 14138 36285 14190
rect 36337 14138 36353 14190
rect 36405 14138 36421 14190
rect 36473 14138 36489 14190
rect 36541 14187 36547 14190
tri 36547 14187 36550 14190 sw
rect 36541 14181 37565 14187
rect 36545 14147 36583 14181
rect 36617 14147 36655 14181
rect 36689 14147 36727 14181
rect 36761 14147 36799 14181
rect 36833 14147 36871 14181
rect 36905 14147 36943 14181
rect 36977 14147 37015 14181
rect 37049 14147 37087 14181
rect 37121 14147 37159 14181
rect 37193 14147 37231 14181
rect 37265 14147 37303 14181
rect 37337 14147 37375 14181
rect 37409 14147 37447 14181
rect 37481 14147 37519 14181
rect 37553 14147 37565 14181
rect 36541 14141 37565 14147
rect 37618 14159 37627 14172
rect 37661 14159 37670 14172
rect 36541 14138 36547 14141
tri 36547 14138 36550 14141 nw
rect 37618 14094 37627 14107
rect 37661 14094 37670 14107
rect 37618 14038 37670 14042
tri 36658 14031 36661 14034 se
rect 36661 14031 36667 14034
rect 35563 14025 36667 14031
rect 36719 14025 36732 14034
rect 35563 13991 35575 14025
rect 35609 13991 35647 14025
rect 35681 13991 35719 14025
rect 35753 13991 35791 14025
rect 35825 13991 35863 14025
rect 35897 13991 35935 14025
rect 35969 13991 36007 14025
rect 36041 13991 36079 14025
rect 36113 13991 36151 14025
rect 36185 13991 36223 14025
rect 36257 13991 36295 14025
rect 36329 13991 36367 14025
rect 36401 13991 36439 14025
rect 36473 13991 36511 14025
rect 36545 13991 36583 14025
rect 36617 13991 36655 14025
rect 36719 13991 36727 14025
rect 35563 13985 36667 13991
tri 36658 13982 36661 13985 ne
rect 36661 13982 36667 13985
rect 36719 13982 36732 13991
rect 36784 13982 36797 14034
rect 36849 13982 36862 14034
rect 36914 13982 36927 14034
rect 36979 13982 36992 14034
rect 37044 14025 37057 14034
rect 37109 14025 37122 14034
rect 37174 14025 37188 14034
rect 37240 14025 37254 14034
rect 37306 14025 37320 14034
rect 37372 14025 37386 14034
rect 37438 14025 37452 14034
rect 37504 14031 37510 14034
tri 37510 14031 37513 14034 sw
rect 37504 14025 37565 14031
rect 37049 13991 37057 14025
rect 37121 13991 37122 14025
rect 37372 13991 37375 14025
rect 37438 13991 37447 14025
rect 37504 13991 37519 14025
rect 37553 13991 37565 14025
rect 37044 13982 37057 13991
rect 37109 13982 37122 13991
rect 37174 13982 37188 13991
rect 37240 13982 37254 13991
rect 37306 13982 37320 13991
rect 37372 13982 37386 13991
rect 37438 13982 37452 13991
rect 37504 13985 37565 13991
rect 37618 14029 37627 14038
rect 37661 14029 37670 14038
rect 37504 13982 37510 13985
tri 37510 13982 37513 13985 nw
rect 37618 13965 37670 13977
rect 37618 13964 37627 13965
rect 37661 13964 37670 13965
rect 37618 13899 37670 13912
tri 35666 13875 35669 13878 se
rect 35669 13875 35675 13878
rect 35563 13869 35675 13875
rect 35727 13869 35742 13878
rect 35794 13869 35809 13878
rect 35861 13869 35877 13878
rect 35929 13869 35945 13878
rect 35997 13869 36013 13878
rect 36065 13869 36081 13878
rect 35563 13835 35575 13869
rect 35609 13835 35647 13869
rect 35861 13835 35863 13869
rect 35929 13835 35935 13869
rect 35997 13835 36007 13869
rect 36065 13835 36079 13869
rect 35563 13829 35675 13835
tri 35666 13826 35669 13829 ne
rect 35669 13826 35675 13829
rect 35727 13826 35742 13835
rect 35794 13826 35809 13835
rect 35861 13826 35877 13835
rect 35929 13826 35945 13835
rect 35997 13826 36013 13835
rect 36065 13826 36081 13835
rect 36133 13826 36149 13878
rect 36201 13826 36217 13878
rect 36269 13826 36285 13878
rect 36337 13826 36353 13878
rect 36405 13826 36421 13878
rect 36473 13826 36489 13878
rect 36541 13875 36547 13878
tri 36547 13875 36550 13878 sw
rect 36541 13869 37565 13875
rect 36545 13835 36583 13869
rect 36617 13835 36655 13869
rect 36689 13835 36727 13869
rect 36761 13835 36799 13869
rect 36833 13835 36871 13869
rect 36905 13835 36943 13869
rect 36977 13835 37015 13869
rect 37049 13835 37087 13869
rect 37121 13835 37159 13869
rect 37193 13835 37231 13869
rect 37265 13835 37303 13869
rect 37337 13835 37375 13869
rect 37409 13835 37447 13869
rect 37481 13835 37519 13869
rect 37553 13835 37565 13869
rect 36541 13829 37565 13835
rect 37618 13834 37670 13847
rect 36541 13826 36547 13829
tri 36547 13826 36550 13829 nw
rect 37618 13769 37670 13782
tri 36658 13719 36661 13722 se
rect 36661 13719 36667 13722
rect 35563 13713 36667 13719
rect 36719 13713 36732 13722
rect 35563 13679 35575 13713
rect 35609 13679 35647 13713
rect 35681 13679 35719 13713
rect 35753 13679 35791 13713
rect 35825 13679 35863 13713
rect 35897 13679 35935 13713
rect 35969 13679 36007 13713
rect 36041 13679 36079 13713
rect 36113 13679 36151 13713
rect 36185 13679 36223 13713
rect 36257 13679 36295 13713
rect 36329 13679 36367 13713
rect 36401 13679 36439 13713
rect 36473 13679 36511 13713
rect 36545 13679 36583 13713
rect 36617 13679 36655 13713
rect 36719 13679 36727 13713
rect 35563 13673 36667 13679
tri 36658 13672 36659 13673 ne
rect 36659 13672 36667 13673
tri 36659 13670 36661 13672 ne
rect 36661 13670 36667 13672
rect 36719 13670 36732 13679
rect 36784 13670 36797 13722
rect 36849 13670 36862 13722
rect 36914 13670 36927 13722
rect 36979 13670 36992 13722
rect 37044 13713 37057 13722
rect 37109 13713 37122 13722
rect 37174 13713 37188 13722
rect 37240 13713 37254 13722
rect 37306 13713 37320 13722
rect 37372 13713 37386 13722
rect 37438 13713 37452 13722
rect 37504 13719 37510 13722
tri 37510 13719 37513 13722 sw
rect 37504 13713 37565 13719
rect 37049 13679 37057 13713
rect 37121 13679 37122 13713
rect 37372 13679 37375 13713
rect 37438 13679 37447 13713
rect 37504 13679 37519 13713
rect 37553 13679 37565 13713
rect 37044 13670 37057 13679
rect 37109 13670 37122 13679
rect 37174 13670 37188 13679
rect 37240 13670 37254 13679
rect 37306 13670 37320 13679
rect 37372 13670 37386 13679
rect 37438 13670 37452 13679
rect 37504 13673 37565 13679
rect 37618 13712 37627 13717
rect 37661 13712 37670 13717
rect 37618 13704 37670 13712
rect 37504 13672 37512 13673
tri 37512 13672 37513 13673 nw
rect 37504 13670 37510 13672
tri 37510 13670 37512 13672 nw
rect 37618 13639 37627 13652
rect 37661 13639 37670 13652
rect 37618 13574 37627 13587
rect 37661 13574 37670 13587
tri 35667 13564 35669 13566 se
rect 35669 13564 35675 13566
tri 35666 13563 35667 13564 se
rect 35667 13563 35675 13564
rect 35563 13557 35675 13563
rect 35727 13557 35742 13566
rect 35794 13557 35809 13566
rect 35861 13557 35877 13566
rect 35929 13557 35945 13566
rect 35997 13557 36013 13566
rect 36065 13557 36081 13566
rect 35563 13523 35575 13557
rect 35609 13523 35647 13557
rect 35861 13523 35863 13557
rect 35929 13523 35935 13557
rect 35997 13523 36007 13557
rect 36065 13523 36079 13557
rect 35563 13517 35675 13523
tri 35666 13514 35669 13517 ne
rect 35669 13514 35675 13517
rect 35727 13514 35742 13523
rect 35794 13514 35809 13523
rect 35861 13514 35877 13523
rect 35929 13514 35945 13523
rect 35997 13514 36013 13523
rect 36065 13514 36081 13523
rect 36133 13514 36149 13566
rect 36201 13514 36217 13566
rect 36269 13514 36285 13566
rect 36337 13514 36353 13566
rect 36405 13514 36421 13566
rect 36473 13514 36489 13566
rect 36541 13564 36547 13566
tri 36547 13564 36549 13566 sw
rect 36541 13563 36549 13564
tri 36549 13563 36550 13564 sw
rect 36541 13557 37565 13563
rect 36545 13523 36583 13557
rect 36617 13523 36655 13557
rect 36689 13523 36727 13557
rect 36761 13523 36799 13557
rect 36833 13523 36871 13557
rect 36905 13523 36943 13557
rect 36977 13523 37015 13557
rect 37049 13523 37087 13557
rect 37121 13523 37159 13557
rect 37193 13523 37231 13557
rect 37265 13523 37303 13557
rect 37337 13523 37375 13557
rect 37409 13523 37447 13557
rect 37481 13523 37519 13557
rect 37553 13523 37565 13557
rect 36541 13517 37565 13523
rect 36541 13514 36547 13517
tri 36547 13514 36550 13517 nw
rect 37618 13509 37627 13522
rect 37661 13509 37670 13522
rect 37618 13450 37670 13457
rect 37618 13444 37627 13450
rect 37661 13444 37670 13450
rect 35495 13410 37565 13422
rect 35495 13401 36667 13410
rect 36719 13401 36732 13410
rect 35495 13367 35575 13401
rect 35609 13367 35647 13401
rect 35681 13367 35719 13401
rect 35753 13367 35791 13401
rect 35825 13367 35863 13401
rect 35897 13367 35935 13401
rect 35969 13367 36007 13401
rect 36041 13367 36079 13401
rect 36113 13367 36151 13401
rect 36185 13367 36223 13401
rect 36257 13367 36295 13401
rect 36329 13367 36367 13401
rect 36401 13367 36439 13401
rect 36473 13367 36511 13401
rect 36545 13367 36583 13401
rect 36617 13367 36655 13401
rect 36719 13367 36727 13401
rect 35495 13358 36667 13367
rect 36719 13358 36732 13367
rect 36784 13358 36797 13410
rect 36849 13358 36862 13410
rect 36914 13358 36927 13410
rect 36979 13358 36992 13410
rect 37044 13401 37057 13410
rect 37109 13401 37122 13410
rect 37174 13401 37188 13410
rect 37240 13401 37254 13410
rect 37306 13401 37320 13410
rect 37372 13401 37386 13410
rect 37438 13401 37452 13410
rect 37504 13401 37565 13410
rect 37049 13367 37057 13401
rect 37121 13367 37122 13401
rect 37372 13367 37375 13401
rect 37438 13367 37447 13401
rect 37504 13367 37519 13401
rect 37553 13367 37565 13401
rect 37044 13358 37057 13367
rect 37109 13358 37122 13367
rect 37174 13358 37188 13367
rect 37240 13358 37254 13367
rect 37306 13358 37320 13367
rect 37372 13358 37386 13367
rect 37438 13358 37452 13367
rect 37504 13358 37565 13367
rect 35495 13342 37565 13358
rect 37618 13379 37670 13392
rect 37618 13314 37670 13327
rect 37618 13256 37670 13262
tri 35666 13251 35669 13254 se
rect 35669 13251 35675 13254
rect 35563 13245 35675 13251
rect 35727 13245 35742 13254
rect 35794 13245 35809 13254
rect 35861 13245 35877 13254
rect 35929 13245 35945 13254
rect 35997 13245 36013 13254
rect 36065 13245 36081 13254
rect 35563 13211 35575 13245
rect 35609 13211 35647 13245
rect 35861 13211 35863 13245
rect 35929 13211 35935 13245
rect 35997 13211 36007 13245
rect 36065 13211 36079 13245
rect 35563 13205 35675 13211
tri 35666 13202 35669 13205 ne
rect 35669 13202 35675 13205
rect 35727 13202 35742 13211
rect 35794 13202 35809 13211
rect 35861 13202 35877 13211
rect 35929 13202 35945 13211
rect 35997 13202 36013 13211
rect 36065 13202 36081 13211
rect 36133 13202 36149 13254
rect 36201 13202 36217 13254
rect 36269 13202 36285 13254
rect 36337 13202 36353 13254
rect 36405 13202 36421 13254
rect 36473 13202 36489 13254
rect 36541 13251 36547 13254
tri 36547 13251 36550 13254 sw
rect 36541 13245 37565 13251
rect 36545 13211 36583 13245
rect 36617 13211 36655 13245
rect 36689 13211 36727 13245
rect 36761 13211 36799 13245
rect 36833 13211 36871 13245
rect 36905 13211 36943 13245
rect 36977 13211 37015 13245
rect 37049 13211 37087 13245
rect 37121 13211 37159 13245
rect 37193 13211 37231 13245
rect 37265 13211 37303 13245
rect 37337 13211 37375 13245
rect 37409 13211 37447 13245
rect 37481 13211 37519 13245
rect 37553 13211 37565 13245
rect 36541 13205 37565 13211
rect 36541 13202 36547 13205
tri 36547 13202 36550 13205 nw
rect 11740 3679 14601 3680
rect 11727 3678 14601 3679
rect 11727 3677 14641 3678
rect 11727 3674 17778 3677
rect 11727 3640 11752 3674
rect 11786 3640 11826 3674
rect 11860 3640 11900 3674
rect 11934 3640 11974 3674
rect 12008 3640 12048 3674
rect 12082 3640 12122 3674
rect 12156 3640 12196 3674
rect 12230 3640 12270 3674
rect 12304 3640 12344 3674
rect 12378 3640 12418 3674
rect 12452 3640 12492 3674
rect 12526 3640 12566 3674
rect 12600 3640 12640 3674
rect 12674 3640 12714 3674
rect 12748 3640 12788 3674
rect 12822 3640 12862 3674
rect 12896 3640 12936 3674
rect 12970 3640 13010 3674
rect 13044 3640 13084 3674
rect 13118 3640 13158 3674
rect 13192 3640 13232 3674
rect 13266 3640 13306 3674
rect 13340 3640 13380 3674
rect 13414 3640 13454 3674
rect 13488 3640 13528 3674
rect 13562 3640 13602 3674
rect 13636 3640 13676 3674
rect 13710 3640 13750 3674
rect 13784 3640 13824 3674
rect 13858 3640 13898 3674
rect 13932 3640 13971 3674
rect 14005 3640 14044 3674
rect 14078 3640 14117 3674
rect 14151 3640 14190 3674
rect 14224 3640 14263 3674
rect 14297 3640 14336 3674
rect 14370 3640 14409 3674
rect 14443 3640 14482 3674
rect 14516 3640 14555 3674
rect 14589 3640 17778 3674
rect 11727 3629 17778 3640
tri 17778 3629 17826 3677 sw
rect 11727 3567 18056 3629
rect 11727 3533 11749 3567
rect 11783 3533 11905 3567
rect 11939 3533 12061 3567
rect 12095 3533 12373 3567
rect 12407 3533 12529 3567
rect 12563 3533 12685 3567
rect 12719 3533 12997 3567
rect 13031 3533 18056 3567
rect 11727 3494 18056 3533
rect 11727 3460 11749 3494
rect 11783 3491 18056 3494
rect 11783 3484 12997 3491
rect 11783 3479 12373 3484
rect 11783 3460 11905 3479
rect 11727 3445 11905 3460
rect 11939 3445 12061 3479
rect 12095 3450 12373 3479
rect 12407 3450 12529 3484
rect 12563 3450 12685 3484
rect 12719 3457 12997 3484
rect 13031 3457 18056 3491
rect 12719 3450 18056 3457
rect 12095 3445 18056 3450
rect 11727 3440 18056 3445
rect 11743 3422 11789 3440
rect 11743 3388 11749 3422
rect 11783 3388 11789 3422
rect 11743 3350 11789 3388
rect 11743 3316 11749 3350
rect 11783 3316 11789 3350
rect 11743 3278 11789 3316
rect 11743 3244 11749 3278
rect 11783 3244 11789 3278
rect 11743 3232 11789 3244
rect 11899 3391 11945 3440
rect 11899 3357 11905 3391
rect 11939 3357 11945 3391
rect 11899 3303 11945 3357
rect 11899 3269 11905 3303
rect 11939 3269 11945 3303
rect 11899 3215 11945 3269
rect 11899 3181 11905 3215
rect 11939 3181 11945 3215
rect 11899 3169 11945 3181
rect 12055 3391 12101 3440
rect 12055 3357 12061 3391
rect 12095 3357 12101 3391
rect 12055 3303 12101 3357
rect 12055 3269 12061 3303
rect 12095 3269 12101 3303
rect 12055 3215 12101 3269
rect 12055 3181 12061 3215
rect 12095 3181 12101 3215
rect 12055 3169 12101 3181
rect 12211 3391 12257 3403
rect 12211 3357 12217 3391
rect 12251 3357 12257 3391
rect 12211 3313 12257 3357
rect 12211 3279 12217 3313
rect 12251 3279 12257 3313
rect 12211 3235 12257 3279
rect 12367 3402 12413 3440
rect 12367 3368 12373 3402
rect 12407 3368 12413 3402
rect 12367 3320 12413 3368
rect 12367 3286 12373 3320
rect 12407 3286 12413 3320
rect 12367 3274 12413 3286
rect 12523 3402 12569 3440
rect 12523 3368 12529 3402
rect 12563 3368 12569 3402
rect 12523 3320 12569 3368
rect 12523 3286 12529 3320
rect 12563 3286 12569 3320
rect 12523 3274 12569 3286
rect 12679 3402 12725 3440
rect 12679 3368 12685 3402
rect 12719 3368 12725 3402
rect 12679 3320 12725 3368
rect 12679 3286 12685 3320
rect 12719 3286 12725 3320
rect 12991 3416 13037 3440
rect 14607 3439 18056 3440
rect 12991 3382 12997 3416
rect 13031 3382 13037 3416
tri 17483 3394 17492 3403 se
rect 17492 3394 17637 3403
rect 12991 3341 13037 3382
rect 12991 3307 12997 3341
rect 13031 3307 13037 3341
rect 12991 3295 13037 3307
rect 13912 3381 17637 3394
rect 13912 3347 13918 3381
rect 13952 3351 17637 3381
rect 17689 3351 17701 3403
rect 17753 3351 17759 3403
rect 17911 3351 17917 3403
rect 17969 3351 17981 3403
rect 18033 3351 18039 3403
rect 13952 3348 17503 3351
tri 17503 3348 17506 3351 nw
rect 13952 3347 13958 3348
rect 13912 3299 13958 3347
rect 17652 3318 17658 3323
rect 12679 3274 12725 3286
rect 12211 3201 12217 3235
rect 12251 3217 12257 3235
rect 13069 3254 13115 3266
rect 13538 3260 13584 3266
rect 13912 3265 13918 3299
rect 13952 3265 13958 3299
rect 14001 3312 17658 3318
rect 14001 3278 14013 3312
rect 14047 3278 14085 3312
rect 14119 3278 17658 3312
rect 14001 3272 17658 3278
rect 17652 3271 17658 3272
rect 17710 3271 17722 3323
rect 17774 3271 17780 3323
rect 13069 3220 13075 3254
rect 13109 3220 13115 3254
rect 13069 3217 13115 3220
rect 13291 3254 13842 3260
rect 13291 3220 13544 3254
rect 13578 3253 13842 3254
tri 13842 3253 13849 3260 sw
rect 13912 3253 13958 3265
rect 13578 3239 13849 3253
tri 13849 3239 13863 3253 sw
rect 13578 3227 13863 3239
tri 13863 3227 13875 3239 sw
rect 14212 3227 14258 3239
rect 13578 3220 13875 3227
rect 13291 3217 13875 3220
tri 13875 3217 13885 3227 sw
rect 14212 3217 14218 3227
rect 12251 3214 14218 3217
rect 12251 3211 13337 3214
rect 12251 3201 12819 3211
rect 12211 3177 12819 3201
rect 12853 3177 12891 3211
rect 12925 3182 13337 3211
rect 12925 3177 13075 3182
rect 12211 3171 13075 3177
rect 12211 3157 12257 3171
rect 12211 3123 12217 3157
rect 12251 3123 12257 3157
rect 13069 3148 13075 3171
rect 13109 3171 13337 3182
rect 13538 3182 13584 3214
tri 13795 3193 13816 3214 ne
rect 13816 3193 14218 3214
rect 14252 3217 14258 3227
rect 14252 3193 14919 3217
rect 13109 3148 13115 3171
rect 13069 3136 13115 3148
rect 13538 3148 13544 3182
rect 13578 3148 13584 3182
tri 13816 3171 13838 3193 ne
rect 13838 3171 14919 3193
rect 13538 3136 13584 3148
rect 13619 3154 13665 3166
rect 12211 3111 12257 3123
rect 13619 3120 13625 3154
rect 13659 3120 13665 3154
rect 13619 3082 13665 3120
rect 13619 3078 13625 3082
rect 11722 3048 13625 3078
rect 13659 3048 13665 3082
rect 11722 3044 13665 3048
rect 11722 2673 11756 3044
rect 13619 3036 13665 3044
rect 13736 3156 13782 3168
rect 13736 3122 13742 3156
rect 13776 3122 13782 3156
rect 13736 3015 13782 3122
rect 14212 3154 14258 3171
rect 14212 3120 14218 3154
rect 14252 3120 14258 3154
rect 14212 3082 14258 3120
rect 14212 3048 14218 3082
rect 14252 3048 14258 3082
rect 14212 3036 14258 3048
rect 13736 3008 13742 3015
rect 13265 3002 13742 3008
rect 13265 2968 13277 3002
rect 13311 2968 13349 3002
rect 13383 2981 13742 3002
rect 13776 3008 13782 3015
rect 13776 2994 14731 3008
rect 13776 2981 14407 2994
rect 13383 2968 14407 2981
rect 13265 2962 14407 2968
rect 11826 2918 12313 2924
rect 11826 2884 11838 2918
rect 11872 2884 11924 2918
rect 11958 2884 12010 2918
rect 12044 2884 12096 2918
rect 12130 2884 12182 2918
rect 12216 2884 12267 2918
rect 12301 2884 12313 2918
rect 11826 2878 12313 2884
rect 12464 2918 12937 2924
rect 12464 2884 12476 2918
rect 12510 2884 12559 2918
rect 12593 2884 12642 2918
rect 12676 2884 12725 2918
rect 12759 2884 12808 2918
rect 12842 2884 12891 2918
rect 12925 2884 12937 2918
rect 12464 2878 12937 2884
rect 13205 2918 13451 2924
rect 13205 2884 13217 2918
rect 13251 2884 13311 2918
rect 13345 2884 13405 2918
rect 13439 2884 13451 2918
rect 13205 2878 13451 2884
rect 13525 2826 13559 2962
tri 14387 2960 14389 2962 ne
rect 14389 2960 14407 2962
rect 14441 2960 14479 2994
rect 14513 2962 14731 2994
rect 14513 2960 14525 2962
tri 14389 2954 14395 2960 ne
rect 14395 2954 14525 2960
tri 14525 2954 14533 2962 nw
rect 13624 2919 14213 2925
rect 13624 2885 13636 2919
rect 13670 2885 13708 2919
rect 13742 2885 14095 2919
rect 14129 2885 14167 2919
rect 14201 2885 14213 2919
rect 13624 2879 14213 2885
rect 14263 2883 14852 2889
rect 14263 2849 14275 2883
rect 14309 2849 14347 2883
rect 14381 2849 14852 2883
rect 14263 2843 14852 2849
tri 13559 2826 13573 2840 sw
tri 13525 2779 13572 2826 ne
rect 13572 2813 13573 2826
tri 13573 2813 13586 2826 sw
rect 13572 2779 15148 2813
rect 12305 2743 13754 2749
rect 12305 2709 12317 2743
rect 12351 2709 12423 2743
rect 12457 2709 12528 2743
rect 12562 2709 13636 2743
rect 13670 2709 13708 2743
rect 13742 2709 13754 2743
rect 12305 2703 13754 2709
tri 14225 2696 14231 2702 se
rect 14231 2696 14690 2702
tri 14221 2692 14225 2696 se
rect 14225 2692 14553 2696
tri 11756 2673 11775 2692 sw
tri 14202 2673 14221 2692 se
rect 14221 2673 14553 2692
rect 11722 2667 11775 2673
tri 11775 2667 11781 2673 sw
rect 12975 2667 14013 2673
rect 11722 2661 11781 2667
tri 11781 2661 11787 2667 sw
rect 12975 2661 13820 2667
rect 11722 2637 11787 2661
tri 11787 2637 11811 2661 sw
tri 11763 2627 11773 2637 ne
rect 11773 2627 11811 2637
tri 11811 2627 11821 2637 sw
rect 12975 2627 12981 2661
rect 13015 2633 13820 2661
rect 13854 2633 13894 2667
rect 13928 2633 13967 2667
rect 14001 2633 14013 2667
tri 14191 2662 14202 2673 se
rect 14202 2662 14553 2673
rect 14587 2662 14625 2696
rect 14659 2662 14690 2696
tri 14186 2657 14191 2662 se
rect 14191 2657 14690 2662
rect 13015 2627 14013 2633
tri 14156 2627 14186 2657 se
rect 14186 2656 14690 2657
rect 14186 2627 14231 2656
tri 11773 2623 11777 2627 ne
rect 11777 2623 11821 2627
tri 11821 2623 11825 2627 sw
tri 11777 2596 11804 2623 ne
rect 11804 2596 11825 2623
tri 11825 2596 11852 2623 sw
rect 12119 2596 12847 2602
tri 11804 2589 11811 2596 ne
rect 11811 2589 11852 2596
tri 11852 2589 11859 2596 sw
tri 11811 2562 11838 2589 ne
rect 11838 2562 11859 2589
tri 11859 2562 11886 2589 sw
rect 12119 2562 12131 2596
rect 12165 2562 12224 2596
rect 12258 2562 12583 2596
rect 12617 2562 12656 2596
rect 12690 2562 12729 2596
rect 12763 2562 12801 2596
rect 12835 2562 12847 2596
tri 11838 2541 11859 2562 ne
rect 11859 2541 11886 2562
tri 11886 2541 11907 2562 sw
tri 11859 2534 11866 2541 ne
rect 11866 2534 11907 2541
tri 11907 2534 11914 2541 sw
tri 11866 2527 11873 2534 ne
rect 11873 2527 11914 2534
tri 11914 2527 11921 2534 sw
tri 11873 2522 11878 2527 ne
rect 11878 2522 11921 2527
tri 11921 2522 11926 2527 sw
tri 11878 2514 11886 2522 ne
rect 11886 2514 11926 2522
tri 11926 2514 11934 2522 sw
rect 12119 2514 12847 2562
tri 11886 2493 11907 2514 ne
rect 11907 2493 11934 2514
tri 11934 2493 11955 2514 sw
tri 11907 2480 11920 2493 ne
rect 11920 2480 11955 2493
tri 11955 2480 11968 2493 sw
rect 12119 2480 12131 2514
rect 12165 2480 12224 2514
rect 12258 2480 12583 2514
rect 12617 2480 12656 2514
rect 12690 2480 12729 2514
rect 12763 2480 12801 2514
rect 12835 2480 12847 2514
tri 11920 2475 11925 2480 ne
rect 11925 2475 11968 2480
tri 11968 2475 11973 2480 sw
tri 11925 2445 11955 2475 ne
rect 11955 2445 11973 2475
tri 11973 2445 12003 2475 sw
rect 12119 2474 12847 2480
rect 12975 2568 13021 2627
tri 14155 2626 14156 2627 se
rect 14156 2626 14231 2627
tri 14231 2626 14261 2656 nw
tri 14152 2623 14155 2626 se
rect 14155 2623 14228 2626
tri 14228 2623 14231 2626 nw
tri 14118 2589 14152 2623 se
rect 14152 2589 14187 2623
tri 14111 2582 14118 2589 se
rect 14118 2582 14187 2589
tri 14187 2582 14228 2623 nw
rect 12975 2534 12981 2568
rect 13015 2534 13021 2568
rect 12975 2475 13021 2534
rect 13702 2550 14155 2582
tri 14155 2550 14187 2582 nw
rect 13702 2528 13771 2550
rect 13539 2522 13771 2528
rect 13539 2488 13551 2522
rect 13585 2488 13638 2522
rect 13672 2488 13725 2522
rect 13759 2488 13771 2522
rect 13539 2482 13771 2488
rect 13848 2516 14401 2522
rect 13848 2482 13860 2516
rect 13894 2482 13942 2516
rect 13976 2482 14024 2516
rect 14058 2482 14106 2516
rect 14140 2482 14189 2516
rect 14223 2482 14272 2516
rect 14306 2482 14355 2516
rect 14389 2482 14401 2516
rect 13848 2476 14401 2482
rect 14493 2514 15038 2520
rect 14493 2480 14505 2514
rect 14539 2480 14586 2514
rect 14620 2480 14667 2514
rect 14701 2480 14748 2514
rect 14782 2480 14829 2514
rect 14863 2480 14910 2514
rect 14944 2480 14992 2514
rect 15026 2480 15038 2514
tri 11955 2441 11959 2445 ne
rect 11959 2441 12003 2445
tri 12003 2441 12007 2445 sw
rect 12975 2441 12981 2475
rect 13015 2441 13021 2475
rect 14111 2474 14169 2476
rect 14493 2474 15038 2480
tri 11959 2423 11977 2441 ne
rect 11977 2440 12007 2441
tri 12007 2440 12008 2441 sw
rect 11977 2426 12008 2440
tri 12008 2426 12022 2440 sw
rect 11977 2423 12022 2426
tri 12022 2423 12025 2426 sw
tri 11977 2421 11979 2423 ne
rect 11979 2421 12025 2423
tri 12025 2421 12027 2423 sw
tri 11979 2420 11980 2421 ne
rect 11980 2420 12027 2421
tri 12027 2420 12028 2421 sw
tri 11980 2407 11993 2420 ne
rect 11993 2407 12028 2420
tri 12028 2407 12041 2420 sw
tri 11993 2405 11995 2407 ne
rect 11995 2260 12041 2407
rect 12975 2382 13021 2441
rect 13328 2457 13374 2469
rect 13328 2423 13334 2457
rect 13368 2423 13374 2457
tri 15100 2426 15114 2440 se
rect 15114 2426 15148 2779
rect 17978 2761 18030 3351
rect 18157 3317 18209 3323
rect 18157 3253 18209 3265
rect 18157 2803 18209 3201
tri 18030 2761 18052 2783 sw
tri 17978 2745 17994 2761 ne
rect 17994 2745 18052 2761
tri 18052 2745 18068 2761 sw
rect 18157 2745 18239 2803
tri 17994 2687 18052 2745 ne
rect 18052 2708 18068 2745
tri 18068 2708 18105 2745 sw
rect 18052 2687 18105 2708
tri 18105 2687 18126 2708 sw
tri 18052 2657 18082 2687 ne
rect 18082 2657 18126 2687
tri 18126 2657 18156 2687 sw
rect 18447 2657 19723 2663
tri 18082 2642 18097 2657 ne
rect 18097 2656 18156 2657
tri 18156 2656 18157 2657 sw
rect 18097 2642 18157 2656
rect 17102 2590 17180 2642
tri 18097 2634 18105 2642 ne
rect 17102 2563 17154 2590
rect 13328 2385 13374 2423
tri 15095 2421 15100 2426 se
rect 15100 2421 15143 2426
tri 15143 2421 15148 2426 nw
rect 15275 2527 17046 2539
rect 15275 2493 15350 2527
rect 15384 2526 16410 2527
rect 15384 2493 15457 2526
rect 15275 2492 15457 2493
rect 15491 2493 16410 2526
rect 16444 2493 17046 2527
rect 15491 2492 17046 2493
rect 15275 2455 17046 2492
rect 15275 2421 15350 2455
rect 15384 2454 16410 2455
rect 15384 2421 15457 2454
tri 15094 2420 15095 2421 se
rect 15095 2420 15142 2421
tri 15142 2420 15143 2421 nw
rect 15275 2420 15457 2421
rect 15491 2421 16410 2454
rect 16444 2421 17046 2455
rect 15491 2420 17046 2421
tri 15075 2401 15094 2420 se
rect 15094 2401 15104 2420
rect 13328 2382 13334 2385
rect 12952 2348 12981 2382
rect 13015 2351 13334 2382
rect 13368 2382 13374 2385
rect 13953 2389 15104 2401
rect 13368 2355 13718 2382
tri 13718 2355 13745 2382 sw
rect 13953 2355 13959 2389
rect 13993 2355 14270 2389
rect 14304 2355 14583 2389
rect 14617 2355 14894 2389
rect 14928 2382 15104 2389
tri 15104 2382 15142 2420 nw
rect 15275 2408 17046 2420
rect 17102 2511 17387 2563
rect 17388 2512 17389 2562
rect 17425 2512 17426 2562
rect 17427 2511 18062 2563
rect 14928 2378 15100 2382
tri 15100 2378 15104 2382 nw
rect 14928 2367 15089 2378
tri 15089 2367 15100 2378 nw
tri 15313 2367 15319 2373 se
rect 15319 2367 16740 2373
rect 14928 2355 15066 2367
rect 13368 2351 13745 2355
rect 13015 2348 13745 2351
rect 12952 2344 13745 2348
tri 13745 2344 13756 2355 sw
rect 13953 2344 15066 2355
tri 15066 2344 15089 2367 nw
tri 15290 2344 15313 2367 se
rect 15313 2344 16622 2367
rect 12952 2336 13756 2344
tri 13700 2333 13703 2336 ne
rect 13703 2333 13756 2336
tri 13756 2333 13767 2344 sw
rect 13953 2333 15055 2344
tri 15055 2333 15066 2344 nw
tri 15279 2333 15290 2344 se
rect 15290 2333 16622 2344
rect 16656 2333 16694 2367
rect 16728 2333 16740 2367
tri 13703 2313 13723 2333 ne
rect 13723 2313 13767 2333
tri 13767 2313 13787 2333 sw
rect 13953 2313 15016 2333
tri 13723 2308 13728 2313 ne
rect 13728 2308 13787 2313
rect 12749 2302 13686 2308
rect 12749 2268 12761 2302
rect 12795 2268 12833 2302
rect 12867 2296 13686 2302
rect 12867 2268 13646 2296
rect 12749 2262 13646 2268
rect 13680 2262 13686 2296
tri 13728 2280 13756 2308 ne
rect 13756 2280 13787 2308
tri 13787 2280 13820 2313 sw
tri 13756 2279 13757 2280 ne
rect 13757 2279 13820 2280
tri 13820 2279 13821 2280 sw
rect 13953 2279 13959 2313
rect 13993 2279 14270 2313
rect 14304 2279 14583 2313
rect 14617 2279 14894 2313
rect 14928 2294 15016 2313
tri 15016 2294 15055 2333 nw
tri 15273 2327 15279 2333 se
rect 15279 2327 16740 2333
tri 15253 2307 15273 2327 se
rect 15273 2307 15319 2327
tri 15319 2307 15339 2327 nw
tri 15240 2294 15253 2307 se
rect 15253 2294 15306 2307
tri 15306 2294 15319 2307 nw
rect 14928 2280 15002 2294
tri 15002 2280 15016 2294 nw
tri 15226 2280 15240 2294 se
rect 15240 2280 15272 2294
rect 14928 2279 14993 2280
tri 12041 2260 12043 2262 sw
rect 11995 2248 12043 2260
tri 12043 2248 12055 2260 sw
rect 11995 2237 12055 2248
tri 12055 2237 12066 2248 sw
rect 11995 2203 12001 2237
rect 12035 2234 12066 2237
tri 12066 2234 12069 2237 sw
rect 12035 2224 12069 2234
tri 12069 2224 12079 2234 sw
tri 13238 2224 13248 2234 se
rect 13248 2224 13294 2234
tri 13294 2224 13304 2234 sw
tri 13396 2224 13406 2234 se
rect 13406 2224 13452 2234
rect 12035 2222 12079 2224
tri 12079 2222 12081 2224 sw
tri 13236 2222 13238 2224 se
rect 13238 2222 13304 2224
tri 13304 2222 13306 2224 sw
tri 13394 2222 13396 2224 se
rect 13396 2222 13452 2224
rect 12035 2213 12081 2222
tri 12081 2213 12090 2222 sw
tri 13227 2213 13236 2222 se
rect 13236 2213 13254 2222
rect 12035 2203 13254 2213
rect 11995 2188 13254 2203
rect 13288 2216 13306 2222
tri 13306 2216 13312 2222 sw
tri 13388 2216 13394 2222 se
rect 13394 2216 13412 2222
rect 13288 2213 13312 2216
tri 13312 2213 13315 2216 sw
tri 13385 2213 13388 2216 se
rect 13388 2213 13412 2216
rect 13288 2188 13412 2213
rect 13446 2188 13452 2222
rect 11995 2167 13452 2188
rect 13640 2224 13686 2262
tri 13757 2260 13776 2279 ne
rect 13776 2260 13821 2279
tri 13821 2260 13840 2279 sw
rect 13953 2271 14993 2279
tri 14993 2271 15002 2280 nw
tri 15217 2271 15226 2280 se
rect 15226 2271 15272 2280
tri 13776 2237 13799 2260 ne
rect 13799 2237 13840 2260
tri 13840 2237 13863 2260 sw
rect 13953 2237 13999 2271
rect 13640 2190 13646 2224
rect 13680 2190 13686 2224
tri 13799 2216 13820 2237 ne
rect 13820 2216 13863 2237
tri 13863 2216 13884 2237 sw
tri 13820 2203 13833 2216 ne
rect 13833 2203 13884 2216
tri 13884 2203 13897 2216 sw
rect 13953 2203 13959 2237
rect 13993 2203 13999 2237
tri 13833 2196 13840 2203 ne
rect 13840 2196 13897 2203
tri 13897 2196 13904 2203 sw
rect 13640 2178 13686 2190
tri 13840 2182 13854 2196 ne
rect 13854 2182 13904 2196
tri 13904 2182 13918 2196 sw
rect 13953 2191 13999 2203
rect 14264 2237 14310 2271
rect 14264 2203 14270 2237
rect 14304 2203 14310 2237
rect 14264 2191 14310 2203
rect 14577 2237 14623 2271
rect 14577 2203 14583 2237
rect 14617 2203 14623 2237
rect 14577 2191 14623 2203
rect 14888 2237 14934 2271
tri 15206 2260 15217 2271 se
rect 15217 2260 15272 2271
tri 15272 2260 15306 2294 nw
tri 15187 2241 15206 2260 se
rect 15206 2241 15253 2260
tri 15253 2241 15272 2260 nw
rect 14888 2203 14894 2237
rect 14928 2203 14934 2237
tri 15182 2236 15187 2241 se
rect 15187 2236 15248 2241
tri 15248 2236 15253 2241 nw
tri 15176 2230 15182 2236 se
rect 15182 2230 15242 2236
tri 15242 2230 15248 2236 nw
rect 16194 2230 16324 2327
tri 15162 2216 15176 2230 se
rect 15176 2216 15208 2230
rect 14888 2191 14934 2203
tri 15142 2196 15162 2216 se
rect 15162 2196 15208 2216
tri 15208 2196 15242 2230 nw
rect 16194 2196 16206 2230
rect 16240 2196 16278 2230
rect 16312 2196 16324 2230
tri 15137 2191 15142 2196 se
rect 15142 2191 15194 2196
tri 15128 2182 15137 2191 se
rect 15137 2182 15194 2191
tri 15194 2182 15208 2196 nw
rect 16194 2190 16324 2196
rect 16786 2216 16916 2222
rect 16786 2182 16798 2216
rect 16832 2182 16870 2216
rect 16904 2182 16916 2216
tri 13854 2178 13858 2182 ne
rect 13858 2178 13918 2182
rect 11995 2160 12053 2167
rect 11995 2126 12001 2160
rect 12035 2152 12053 2160
tri 12053 2152 12068 2167 nw
tri 13215 2152 13230 2167 ne
rect 13230 2152 13305 2167
tri 13305 2152 13320 2167 nw
tri 13370 2152 13385 2167 ne
rect 13385 2152 13452 2167
tri 13858 2159 13877 2178 ne
rect 13877 2159 13918 2178
rect 12035 2150 12051 2152
tri 12051 2150 12053 2152 nw
tri 13230 2150 13232 2152 ne
rect 13232 2150 13303 2152
tri 13303 2150 13305 2152 nw
tri 13385 2150 13387 2152 ne
rect 13387 2150 13452 2152
rect 12035 2126 12041 2150
tri 12041 2140 12051 2150 nw
tri 13232 2140 13242 2150 ne
rect 13242 2140 13254 2150
tri 13242 2134 13248 2140 ne
rect 11995 2083 12041 2126
rect 11995 2049 12001 2083
rect 12035 2049 12041 2083
rect 11995 2037 12041 2049
rect 12633 2124 12763 2130
rect 12633 2090 12645 2124
rect 12679 2090 12717 2124
rect 12751 2090 12763 2124
rect 13248 2116 13254 2140
rect 13288 2116 13294 2150
tri 13294 2141 13303 2150 nw
tri 13387 2141 13396 2150 ne
rect 13396 2141 13412 2150
tri 13396 2131 13406 2141 ne
rect 13248 2104 13294 2116
rect 13406 2116 13412 2141
rect 13446 2116 13452 2150
rect 13406 2104 13452 2116
rect 13561 2156 13607 2159
tri 13607 2156 13610 2159 sw
rect 13561 2148 13610 2156
tri 13610 2148 13618 2156 sw
tri 13713 2148 13721 2156 se
rect 13721 2148 13767 2159
tri 13877 2152 13884 2159 ne
rect 13884 2152 13918 2159
tri 13918 2152 13948 2182 sw
tri 15121 2175 15128 2182 se
rect 15128 2175 15187 2182
tri 15187 2175 15194 2182 nw
rect 16786 2176 16916 2182
tri 15098 2152 15121 2175 se
rect 15121 2152 15164 2175
tri 15164 2152 15187 2175 nw
tri 13884 2148 13888 2152 ne
rect 13888 2148 15160 2152
tri 15160 2148 15164 2152 nw
rect 13561 2147 13618 2148
tri 13618 2147 13619 2148 sw
tri 13712 2147 13713 2148 se
rect 13713 2147 13767 2148
rect 13561 2113 13567 2147
rect 13601 2143 13619 2147
tri 13619 2143 13623 2147 sw
tri 13708 2143 13712 2147 se
rect 13712 2143 13727 2147
rect 13601 2113 13727 2143
rect 13761 2113 13767 2147
tri 13888 2143 13893 2148 ne
rect 13893 2143 15155 2148
tri 15155 2143 15160 2148 nw
rect 15881 2143 16331 2149
tri 13559 2100 13561 2102 se
rect 13561 2100 13767 2113
tri 13893 2112 13924 2143 ne
rect 13924 2112 15121 2143
rect 12633 1999 12763 2090
tri 13535 2076 13559 2100 se
rect 13559 2076 13767 2100
rect 12950 2075 13767 2076
rect 12950 2070 13567 2075
rect 12950 2036 12962 2070
rect 12996 2036 13034 2070
rect 13068 2041 13567 2070
rect 13601 2041 13727 2075
rect 13761 2041 13767 2075
rect 13068 2036 13767 2041
rect 12950 2030 13767 2036
rect 13561 2029 13607 2030
rect 13721 2029 13767 2030
rect 13796 2100 13842 2112
tri 13924 2109 13927 2112 ne
rect 13927 2109 15121 2112
tri 15121 2109 15155 2143 nw
rect 15881 2109 15893 2143
rect 15927 2109 15966 2143
rect 16000 2109 16212 2143
rect 16246 2109 16285 2143
rect 16319 2109 16331 2143
tri 13927 2106 13930 2109 ne
rect 13930 2106 15118 2109
tri 15118 2106 15121 2109 nw
rect 15881 2103 16331 2109
rect 16971 2104 17001 2408
rect 13796 2066 13802 2100
rect 13836 2066 13842 2100
rect 17102 2075 17154 2511
rect 17927 2479 18062 2511
rect 17605 2473 17787 2479
rect 17789 2478 17825 2479
rect 17268 2104 17298 2456
rect 17605 2439 17617 2473
rect 17651 2439 17689 2473
rect 17723 2439 17787 2473
rect 17605 2433 17787 2439
rect 17788 2434 17826 2478
rect 17789 2433 17825 2434
rect 17827 2433 18062 2479
rect 17920 2394 18062 2433
rect 17920 2382 18050 2394
tri 18050 2382 18062 2394 nw
rect 17920 2378 18046 2382
tri 18046 2378 18050 2382 nw
rect 17920 2373 18041 2378
tri 18041 2373 18046 2378 nw
rect 17920 2368 18036 2373
tri 18036 2368 18041 2373 nw
rect 17920 2348 18016 2368
tri 18016 2348 18036 2368 nw
tri 18085 2348 18105 2368 se
rect 18105 2348 18157 2642
rect 18447 2623 18459 2657
rect 18493 2623 18536 2657
rect 18570 2623 18613 2657
rect 18647 2623 18689 2657
rect 18723 2623 18765 2657
rect 18799 2623 18841 2657
rect 18875 2623 18917 2657
rect 18951 2623 18993 2657
rect 19027 2623 19069 2657
rect 19103 2623 19145 2657
rect 19179 2623 19221 2657
rect 19255 2623 19297 2657
rect 19331 2623 19373 2657
rect 19407 2623 19449 2657
rect 19483 2623 19525 2657
rect 19559 2623 19601 2657
rect 19635 2623 19677 2657
rect 19711 2623 19723 2657
rect 18447 2617 19723 2623
tri 17899 2327 17920 2348 se
rect 17920 2327 17995 2348
tri 17995 2327 18016 2348 nw
tri 18064 2327 18085 2348 se
rect 18085 2346 18157 2348
rect 18085 2327 18111 2346
tri 17866 2294 17899 2327 se
rect 17899 2325 17993 2327
tri 17993 2325 17995 2327 nw
tri 18062 2325 18064 2327 se
rect 18064 2325 18111 2327
rect 17899 2294 17962 2325
tri 17962 2294 17993 2325 nw
tri 18031 2294 18062 2325 se
rect 18062 2300 18111 2325
tri 18111 2300 18157 2346 nw
rect 19672 2300 19678 2303
rect 18062 2294 18105 2300
tri 18105 2294 18111 2300 nw
tri 18203 2294 18209 2300 se
rect 18209 2294 19678 2300
tri 17859 2287 17866 2294 se
rect 17866 2287 17955 2294
tri 17955 2287 17962 2294 nw
tri 18024 2287 18031 2294 se
rect 18031 2287 18071 2294
rect 17859 2260 17928 2287
tri 17928 2260 17955 2287 nw
tri 17997 2260 18024 2287 se
rect 18024 2260 18071 2287
tri 18071 2260 18105 2294 nw
tri 18169 2260 18203 2294 se
rect 18203 2260 18442 2294
rect 18476 2260 18515 2294
rect 18549 2260 18588 2294
rect 18622 2260 18661 2294
rect 18695 2260 18734 2294
rect 18768 2260 18807 2294
rect 18841 2260 18880 2294
rect 18914 2260 18953 2294
rect 18987 2260 19026 2294
rect 19060 2260 19099 2294
rect 19133 2260 19172 2294
rect 19206 2260 19245 2294
rect 19279 2260 19318 2294
rect 19352 2260 19391 2294
rect 19425 2260 19464 2294
rect 19498 2260 19537 2294
rect 19571 2260 19610 2294
rect 19644 2260 19678 2294
rect 13796 2013 13842 2066
rect 13796 1999 13802 2013
rect 11959 1987 13802 1999
rect 11959 1953 13178 1987
rect 13212 1953 13490 1987
rect 13524 1979 13802 1987
rect 13836 1999 13842 2013
rect 14108 2056 14154 2068
rect 14108 2022 14114 2056
rect 14148 2022 14154 2056
rect 14108 1999 14154 2022
rect 14420 2056 14466 2068
rect 14420 2022 14426 2056
rect 14460 2022 14466 2056
rect 14420 1999 14466 2022
rect 14732 2056 14778 2068
rect 14732 2022 14738 2056
rect 14772 2022 14778 2056
rect 14732 1999 14778 2022
rect 15044 2056 15090 2068
rect 15044 2022 15050 2056
rect 15084 2022 15090 2056
rect 16052 2067 16628 2075
rect 16630 2074 16666 2075
rect 16052 2033 16064 2067
rect 16098 2033 16137 2067
rect 16171 2033 16628 2067
rect 16052 2027 16628 2033
rect 16629 2028 16667 2074
rect 16630 2027 16666 2028
rect 16668 2027 17154 2075
rect 15044 1999 15090 2022
rect 17222 1999 17498 2104
rect 17859 2068 17922 2260
tri 17922 2254 17928 2260 nw
tri 17991 2254 17997 2260 se
rect 17997 2254 18065 2260
tri 18065 2254 18071 2260 nw
tri 18163 2254 18169 2260 se
rect 18169 2254 19678 2260
tri 17973 2236 17991 2254 se
rect 17991 2236 18031 2254
tri 17957 2220 17973 2236 se
rect 17973 2220 18031 2236
tri 18031 2220 18065 2254 nw
tri 18160 2251 18163 2254 se
rect 18163 2251 18226 2254
tri 18226 2251 18229 2254 nw
rect 19672 2251 19678 2254
rect 19730 2251 19742 2303
rect 19794 2251 19800 2303
tri 18151 2242 18160 2251 se
rect 18160 2242 18217 2251
tri 18217 2242 18226 2251 nw
rect 23077 2242 23083 2294
rect 23135 2242 23155 2294
rect 23207 2242 23227 2294
rect 23279 2242 23299 2294
rect 23351 2242 23371 2294
rect 23423 2242 23442 2294
rect 23494 2242 23513 2294
rect 23565 2242 23584 2294
rect 23636 2242 23642 2294
tri 18143 2234 18151 2242 se
rect 18151 2234 18209 2242
tri 18209 2234 18217 2242 nw
tri 18129 2220 18143 2234 se
rect 18143 2220 18177 2234
rect 17773 2016 17779 2068
rect 17831 2016 17843 2068
rect 17895 2037 17922 2068
rect 17895 2016 17901 2037
tri 17901 2016 17922 2037 nw
tri 17954 2217 17957 2220 se
rect 17957 2217 18028 2220
tri 18028 2217 18031 2220 nw
tri 18126 2217 18129 2220 se
rect 18129 2217 18177 2220
rect 13836 1993 17498 1999
rect 13836 1984 15370 1993
rect 13836 1979 14114 1984
rect 13524 1953 14114 1979
rect 11959 1950 14114 1953
rect 14148 1950 14426 1984
rect 14460 1950 14738 1984
rect 14772 1950 15050 1984
rect 15084 1959 15370 1984
rect 15404 1959 15465 1993
rect 15499 1959 15559 1993
rect 15593 1987 17498 1993
rect 17954 1987 18006 2217
tri 18006 2195 18028 2217 nw
tri 18111 2202 18126 2217 se
rect 18126 2202 18177 2217
tri 18177 2202 18209 2234 nw
rect 18111 2195 18170 2202
tri 18170 2195 18177 2202 nw
rect 18111 2011 18157 2195
tri 18157 2182 18170 2195 nw
rect 20422 2105 20428 2157
rect 20480 2105 20492 2157
rect 20544 2154 20550 2157
rect 20544 2148 23599 2154
rect 20544 2114 20580 2148
rect 20614 2114 20653 2148
rect 20687 2114 20726 2148
rect 20760 2114 20799 2148
rect 20833 2114 20872 2148
rect 20906 2114 20945 2148
rect 20979 2114 21018 2148
rect 21052 2114 21091 2148
rect 21125 2114 21164 2148
rect 21198 2114 21237 2148
rect 21271 2114 21310 2148
rect 21344 2114 21383 2148
rect 21417 2114 21456 2148
rect 21490 2114 21529 2148
rect 21563 2114 21602 2148
rect 21636 2114 21675 2148
rect 21709 2114 21748 2148
rect 21782 2114 21821 2148
rect 21855 2114 21894 2148
rect 21928 2114 21967 2148
rect 22001 2114 22040 2148
rect 22074 2114 22113 2148
rect 22147 2114 22185 2148
rect 22219 2114 22257 2148
rect 22291 2114 22329 2148
rect 22363 2114 22401 2148
rect 22435 2114 22473 2148
rect 22507 2114 22545 2148
rect 22579 2114 22617 2148
rect 22651 2114 22689 2148
rect 22723 2114 22761 2148
rect 22795 2114 22833 2148
rect 22867 2114 22905 2148
rect 22939 2114 22977 2148
rect 23011 2114 23049 2148
rect 23083 2114 23121 2148
rect 23155 2114 23193 2148
rect 23227 2114 23265 2148
rect 23299 2114 23337 2148
rect 23371 2114 23409 2148
rect 23443 2114 23481 2148
rect 23515 2114 23553 2148
rect 23587 2114 23599 2148
rect 20544 2108 23599 2114
rect 20544 2105 20550 2108
tri 19472 2012 19483 2023 ne
rect 19483 2012 19566 2023
tri 18157 2011 18158 2012 sw
tri 19483 2011 19484 2012 ne
rect 19484 2011 19566 2012
rect 18111 1987 18158 2011
tri 18158 1987 18182 2011 sw
tri 19484 1987 19508 2011 ne
rect 19508 1987 19566 2011
tri 19566 1987 19602 2023 nw
rect 15593 1959 16411 1987
rect 15084 1953 16411 1959
rect 16445 1953 17498 1987
rect 15084 1950 17498 1953
rect 11959 1926 17498 1950
rect 17909 1935 17915 1987
rect 17967 1935 17979 1987
rect 18031 1935 18037 1987
rect 18111 1982 18182 1987
tri 18182 1982 18187 1987 sw
tri 18111 1981 18112 1982 ne
rect 18112 1981 18187 1982
tri 18187 1981 18188 1982 sw
tri 18112 1975 18118 1981 ne
rect 18118 1975 19356 1981
tri 18118 1941 18152 1975 ne
rect 18152 1941 18459 1975
rect 18493 1941 18537 1975
rect 18571 1941 18615 1975
rect 18649 1941 18693 1975
rect 18727 1941 18771 1975
rect 18805 1941 18848 1975
rect 18882 1941 18925 1975
rect 18959 1941 19002 1975
rect 19036 1941 19079 1975
rect 19113 1941 19156 1975
rect 19190 1941 19233 1975
rect 19267 1941 19310 1975
rect 19344 1941 19356 1975
tri 18152 1935 18158 1941 ne
rect 18158 1935 19356 1941
rect 11959 1917 13802 1926
rect 11959 1883 12495 1917
rect 12529 1913 13802 1917
rect 12529 1883 13178 1913
rect 11959 1879 13178 1883
rect 13212 1879 13490 1913
rect 13524 1892 13802 1913
rect 13836 1915 17498 1926
rect 13836 1912 16411 1915
rect 13836 1892 14114 1912
rect 13524 1879 14114 1892
rect 11959 1878 14114 1879
rect 14148 1878 14426 1912
rect 14460 1878 14738 1912
rect 14772 1878 15050 1912
rect 15084 1881 16411 1912
rect 16445 1881 17498 1915
tri 19476 1892 19511 1927 se
rect 19511 1892 19566 1927
tri 19566 1892 19601 1927 sw
rect 15084 1878 17498 1881
rect 11959 1873 17498 1878
rect 11959 1845 15370 1873
rect 11959 1811 12495 1845
rect 12529 1840 15370 1845
rect 12529 1811 13178 1840
rect 11959 1806 13178 1811
rect 13212 1806 13490 1840
rect 13524 1806 13802 1840
rect 13836 1806 14114 1840
rect 14148 1806 14426 1840
rect 14460 1806 14738 1840
rect 14772 1806 15050 1840
rect 15084 1839 15370 1840
rect 15404 1839 15465 1873
rect 15499 1839 15559 1873
rect 15593 1839 17498 1873
rect 15084 1806 17498 1839
rect 11959 1757 17498 1806
rect 11959 1723 12141 1757
rect 12175 1723 12214 1757
rect 12248 1723 12287 1757
rect 12321 1723 12360 1757
rect 12394 1723 12433 1757
rect 12467 1723 12506 1757
rect 12540 1723 12579 1757
rect 12613 1723 12652 1757
rect 12686 1723 12725 1757
rect 12759 1723 12798 1757
rect 12832 1723 12871 1757
rect 12905 1723 12944 1757
rect 12978 1723 13017 1757
rect 13051 1723 13090 1757
rect 13124 1723 13163 1757
rect 13197 1723 13236 1757
rect 13270 1723 13309 1757
rect 13343 1723 13382 1757
rect 13416 1723 13455 1757
rect 13489 1723 13528 1757
rect 13562 1723 13601 1757
rect 13635 1723 13674 1757
rect 13708 1723 13747 1757
rect 13781 1723 13820 1757
rect 13854 1723 13893 1757
rect 13927 1723 13966 1757
rect 14000 1723 14039 1757
rect 14073 1723 14112 1757
rect 14146 1723 14185 1757
rect 14219 1723 14258 1757
rect 14292 1723 14331 1757
rect 14365 1723 14404 1757
rect 14438 1723 14477 1757
rect 14511 1723 14550 1757
rect 14584 1723 14623 1757
rect 14657 1723 14696 1757
rect 14730 1723 14769 1757
rect 14803 1723 14842 1757
rect 14876 1723 14915 1757
rect 14949 1723 14988 1757
rect 15022 1723 15061 1757
rect 15095 1723 15134 1757
rect 15168 1723 15207 1757
rect 15241 1723 15280 1757
rect 15314 1723 15353 1757
rect 15387 1723 15426 1757
rect 15460 1723 15498 1757
rect 15532 1723 15570 1757
rect 15604 1723 15642 1757
rect 15676 1723 15714 1757
rect 15748 1723 15786 1757
rect 15820 1723 17498 1757
rect 11959 1716 17498 1723
rect 18113 1752 20495 1892
tri 20495 1810 20577 1892 sw
rect 18113 1716 20792 1752
tri 20792 1716 20828 1752 nw
rect 18113 1698 20774 1716
tri 20774 1698 20792 1716 nw
rect 18113 1692 20768 1698
tri 20768 1692 20774 1698 nw
rect 20947 1692 23607 1698
rect 18113 1691 20755 1692
rect 18113 1657 18160 1691
rect 18194 1657 18232 1691
rect 18266 1657 18304 1691
rect 18338 1657 18376 1691
rect 18410 1657 18448 1691
rect 18482 1657 18520 1691
rect 18554 1657 18592 1691
rect 18626 1657 18664 1691
rect 18698 1657 18736 1691
rect 18770 1657 18808 1691
rect 18842 1657 18880 1691
rect 18914 1657 18952 1691
rect 18986 1657 19024 1691
rect 19058 1657 19096 1691
rect 19130 1657 19168 1691
rect 19202 1657 19240 1691
rect 19274 1657 19312 1691
rect 19346 1657 19384 1691
rect 19418 1657 19456 1691
rect 19490 1657 19528 1691
rect 19562 1657 19600 1691
rect 19634 1657 19672 1691
rect 19706 1657 19744 1691
rect 19778 1657 19816 1691
rect 19850 1657 19888 1691
rect 19922 1657 19960 1691
rect 19994 1657 20032 1691
rect 20066 1657 20104 1691
rect 20138 1657 20176 1691
rect 20210 1657 20248 1691
rect 20282 1657 20320 1691
rect 20354 1657 20392 1691
rect 20426 1679 20464 1691
rect 20498 1679 20536 1691
rect 20570 1679 20608 1691
rect 20642 1679 20680 1691
rect 20714 1679 20755 1691
tri 20755 1679 20768 1692 nw
rect 20947 1679 20977 1692
rect 21011 1679 21051 1692
rect 20452 1657 20464 1679
rect 18113 1648 20400 1657
rect 20394 1627 20400 1648
rect 20452 1627 20467 1657
rect 20519 1627 20534 1679
rect 20586 1627 20600 1679
rect 20652 1627 20666 1679
rect 20718 1658 20734 1679
tri 20734 1658 20755 1679 nw
rect 20718 1651 20727 1658
tri 20727 1651 20734 1658 nw
rect 20718 1627 20724 1651
tri 20724 1648 20727 1651 nw
rect 20947 1627 20953 1679
rect 21011 1658 21017 1679
rect 21085 1658 21125 1692
rect 21159 1658 21199 1692
rect 21233 1658 21273 1692
rect 21307 1658 21347 1692
rect 21381 1658 21421 1692
rect 21455 1658 21495 1692
rect 21529 1658 21569 1692
rect 21603 1658 21643 1692
rect 21677 1658 21717 1692
rect 21751 1658 21791 1692
rect 21825 1658 21865 1692
rect 21899 1658 21939 1692
rect 21973 1658 22013 1692
rect 22047 1658 22087 1692
rect 22121 1658 22161 1692
rect 22195 1658 22235 1692
rect 22269 1658 22309 1692
rect 22343 1658 22383 1692
rect 22417 1658 22457 1692
rect 22491 1658 22531 1692
rect 22565 1658 22605 1692
rect 22639 1658 22679 1692
rect 22713 1658 22753 1692
rect 22787 1658 22827 1692
rect 22861 1658 22901 1692
rect 22935 1658 22975 1692
rect 23009 1658 23049 1692
rect 23083 1658 23123 1692
rect 23157 1658 23196 1692
rect 23230 1658 23269 1692
rect 23303 1658 23342 1692
rect 23376 1658 23415 1692
rect 23449 1658 23488 1692
rect 23522 1658 23561 1692
rect 23595 1658 23607 1692
rect 21005 1627 21017 1658
rect 21069 1652 23607 1658
rect 21069 1627 21075 1652
<< rmetal1 >>
rect 17387 2562 17389 2563
rect 17387 2512 17388 2562
rect 17387 2511 17389 2512
rect 17425 2562 17427 2563
rect 17426 2512 17427 2562
rect 17425 2511 17427 2512
rect 17787 2478 17789 2479
rect 17825 2478 17827 2479
rect 17787 2434 17788 2478
rect 17826 2434 17827 2478
rect 17787 2433 17789 2434
rect 17825 2433 17827 2434
rect 16628 2074 16630 2075
rect 16666 2074 16668 2075
rect 16628 2028 16629 2074
rect 16667 2028 16668 2074
rect 16628 2027 16630 2028
rect 16666 2027 16668 2028
<< via1 >>
rect 37702 16105 37754 16157
rect 37702 16041 37754 16093
rect 37702 15977 37754 16029
rect 35675 15117 35727 15126
rect 35742 15117 35794 15126
rect 35809 15117 35861 15126
rect 35877 15117 35929 15126
rect 35945 15117 35997 15126
rect 36013 15117 36065 15126
rect 36081 15117 36133 15126
rect 35675 15083 35681 15117
rect 35681 15083 35719 15117
rect 35719 15083 35727 15117
rect 35742 15083 35753 15117
rect 35753 15083 35791 15117
rect 35791 15083 35794 15117
rect 35809 15083 35825 15117
rect 35825 15083 35861 15117
rect 35877 15083 35897 15117
rect 35897 15083 35929 15117
rect 35945 15083 35969 15117
rect 35969 15083 35997 15117
rect 36013 15083 36041 15117
rect 36041 15083 36065 15117
rect 36081 15083 36113 15117
rect 36113 15083 36133 15117
rect 35675 15074 35727 15083
rect 35742 15074 35794 15083
rect 35809 15074 35861 15083
rect 35877 15074 35929 15083
rect 35945 15074 35997 15083
rect 36013 15074 36065 15083
rect 36081 15074 36133 15083
rect 36149 15117 36201 15126
rect 36149 15083 36151 15117
rect 36151 15083 36185 15117
rect 36185 15083 36201 15117
rect 36149 15074 36201 15083
rect 36217 15117 36269 15126
rect 36217 15083 36223 15117
rect 36223 15083 36257 15117
rect 36257 15083 36269 15117
rect 36217 15074 36269 15083
rect 36285 15117 36337 15126
rect 36285 15083 36295 15117
rect 36295 15083 36329 15117
rect 36329 15083 36337 15117
rect 36285 15074 36337 15083
rect 36353 15117 36405 15126
rect 36353 15083 36367 15117
rect 36367 15083 36401 15117
rect 36401 15083 36405 15117
rect 36353 15074 36405 15083
rect 36421 15117 36473 15126
rect 36421 15083 36439 15117
rect 36439 15083 36473 15117
rect 36421 15074 36473 15083
rect 36489 15117 36541 15126
rect 36489 15083 36511 15117
rect 36511 15083 36541 15117
rect 36489 15074 36541 15083
rect 37618 15060 37670 15066
rect 37618 15026 37627 15060
rect 37627 15026 37661 15060
rect 37661 15026 37670 15060
rect 37618 15014 37670 15026
rect 37618 14987 37670 15002
rect 36667 14961 36719 14970
rect 36732 14961 36784 14970
rect 36667 14927 36689 14961
rect 36689 14927 36719 14961
rect 36732 14927 36761 14961
rect 36761 14927 36784 14961
rect 36667 14918 36719 14927
rect 36732 14918 36784 14927
rect 36797 14961 36849 14970
rect 36797 14927 36799 14961
rect 36799 14927 36833 14961
rect 36833 14927 36849 14961
rect 36797 14918 36849 14927
rect 36862 14961 36914 14970
rect 36862 14927 36871 14961
rect 36871 14927 36905 14961
rect 36905 14927 36914 14961
rect 36862 14918 36914 14927
rect 36927 14961 36979 14970
rect 36927 14927 36943 14961
rect 36943 14927 36977 14961
rect 36977 14927 36979 14961
rect 36927 14918 36979 14927
rect 36992 14961 37044 14970
rect 37057 14961 37109 14970
rect 37122 14961 37174 14970
rect 37188 14961 37240 14970
rect 37254 14961 37306 14970
rect 37320 14961 37372 14970
rect 37386 14961 37438 14970
rect 37452 14961 37504 14970
rect 36992 14927 37015 14961
rect 37015 14927 37044 14961
rect 37057 14927 37087 14961
rect 37087 14927 37109 14961
rect 37122 14927 37159 14961
rect 37159 14927 37174 14961
rect 37188 14927 37193 14961
rect 37193 14927 37231 14961
rect 37231 14927 37240 14961
rect 37254 14927 37265 14961
rect 37265 14927 37303 14961
rect 37303 14927 37306 14961
rect 37320 14927 37337 14961
rect 37337 14927 37372 14961
rect 37386 14927 37409 14961
rect 37409 14927 37438 14961
rect 37452 14927 37481 14961
rect 37481 14927 37504 14961
rect 36992 14918 37044 14927
rect 37057 14918 37109 14927
rect 37122 14918 37174 14927
rect 37188 14918 37240 14927
rect 37254 14918 37306 14927
rect 37320 14918 37372 14927
rect 37386 14918 37438 14927
rect 37452 14918 37504 14927
rect 37618 14953 37627 14987
rect 37627 14953 37661 14987
rect 37661 14953 37670 14987
rect 37618 14950 37670 14953
rect 37618 14914 37670 14938
rect 37618 14886 37627 14914
rect 37627 14886 37661 14914
rect 37661 14886 37670 14914
rect 37618 14841 37670 14874
rect 37618 14822 37627 14841
rect 37627 14822 37661 14841
rect 37661 14822 37670 14841
rect 35675 14805 35727 14814
rect 35742 14805 35794 14814
rect 35809 14805 35861 14814
rect 35877 14805 35929 14814
rect 35945 14805 35997 14814
rect 36013 14805 36065 14814
rect 36081 14805 36133 14814
rect 35675 14771 35681 14805
rect 35681 14771 35719 14805
rect 35719 14771 35727 14805
rect 35742 14771 35753 14805
rect 35753 14771 35791 14805
rect 35791 14771 35794 14805
rect 35809 14771 35825 14805
rect 35825 14771 35861 14805
rect 35877 14771 35897 14805
rect 35897 14771 35929 14805
rect 35945 14771 35969 14805
rect 35969 14771 35997 14805
rect 36013 14771 36041 14805
rect 36041 14771 36065 14805
rect 36081 14771 36113 14805
rect 36113 14771 36133 14805
rect 35675 14762 35727 14771
rect 35742 14762 35794 14771
rect 35809 14762 35861 14771
rect 35877 14762 35929 14771
rect 35945 14762 35997 14771
rect 36013 14762 36065 14771
rect 36081 14762 36133 14771
rect 36149 14805 36201 14814
rect 36149 14771 36151 14805
rect 36151 14771 36185 14805
rect 36185 14771 36201 14805
rect 36149 14762 36201 14771
rect 36217 14805 36269 14814
rect 36217 14771 36223 14805
rect 36223 14771 36257 14805
rect 36257 14771 36269 14805
rect 36217 14762 36269 14771
rect 36285 14805 36337 14814
rect 36285 14771 36295 14805
rect 36295 14771 36329 14805
rect 36329 14771 36337 14805
rect 36285 14762 36337 14771
rect 36353 14805 36405 14814
rect 36353 14771 36367 14805
rect 36367 14771 36401 14805
rect 36401 14771 36405 14805
rect 36353 14762 36405 14771
rect 36421 14805 36473 14814
rect 36421 14771 36439 14805
rect 36439 14771 36473 14805
rect 36421 14762 36473 14771
rect 36489 14805 36541 14814
rect 36489 14771 36511 14805
rect 36511 14771 36541 14805
rect 36489 14762 36541 14771
rect 37618 14807 37627 14809
rect 37627 14807 37661 14809
rect 37661 14807 37670 14809
rect 37618 14768 37670 14807
rect 37618 14757 37627 14768
rect 37627 14757 37661 14768
rect 37661 14757 37670 14768
rect 37618 14734 37627 14744
rect 37627 14734 37661 14744
rect 37661 14734 37670 14744
rect 37618 14695 37670 14734
rect 37618 14692 37627 14695
rect 37627 14692 37661 14695
rect 37661 14692 37670 14695
rect 37618 14661 37627 14679
rect 37627 14661 37661 14679
rect 37661 14661 37670 14679
rect 36667 14649 36719 14658
rect 36732 14649 36784 14658
rect 36667 14615 36689 14649
rect 36689 14615 36719 14649
rect 36732 14615 36761 14649
rect 36761 14615 36784 14649
rect 36667 14606 36719 14615
rect 36732 14606 36784 14615
rect 36797 14649 36849 14658
rect 36797 14615 36799 14649
rect 36799 14615 36833 14649
rect 36833 14615 36849 14649
rect 36797 14606 36849 14615
rect 36862 14649 36914 14658
rect 36862 14615 36871 14649
rect 36871 14615 36905 14649
rect 36905 14615 36914 14649
rect 36862 14606 36914 14615
rect 36927 14649 36979 14658
rect 36927 14615 36943 14649
rect 36943 14615 36977 14649
rect 36977 14615 36979 14649
rect 36927 14606 36979 14615
rect 36992 14649 37044 14658
rect 37057 14649 37109 14658
rect 37122 14649 37174 14658
rect 37188 14649 37240 14658
rect 37254 14649 37306 14658
rect 37320 14649 37372 14658
rect 37386 14649 37438 14658
rect 37452 14649 37504 14658
rect 36992 14615 37015 14649
rect 37015 14615 37044 14649
rect 37057 14615 37087 14649
rect 37087 14615 37109 14649
rect 37122 14615 37159 14649
rect 37159 14615 37174 14649
rect 37188 14615 37193 14649
rect 37193 14615 37231 14649
rect 37231 14615 37240 14649
rect 37254 14615 37265 14649
rect 37265 14615 37303 14649
rect 37303 14615 37306 14649
rect 37320 14615 37337 14649
rect 37337 14615 37372 14649
rect 37386 14615 37409 14649
rect 37409 14615 37438 14649
rect 37452 14615 37481 14649
rect 37481 14615 37504 14649
rect 36992 14606 37044 14615
rect 37057 14606 37109 14615
rect 37122 14606 37174 14615
rect 37188 14606 37240 14615
rect 37254 14606 37306 14615
rect 37320 14606 37372 14615
rect 37386 14606 37438 14615
rect 37452 14606 37504 14615
rect 37618 14627 37670 14661
rect 37618 14588 37627 14614
rect 37627 14588 37661 14614
rect 37661 14588 37670 14614
rect 37618 14562 37670 14588
rect 37618 14515 37627 14549
rect 37627 14515 37661 14549
rect 37661 14515 37670 14549
rect 35675 14493 35727 14502
rect 35742 14493 35794 14502
rect 35809 14493 35861 14502
rect 35877 14493 35929 14502
rect 35945 14493 35997 14502
rect 36013 14493 36065 14502
rect 36081 14493 36133 14502
rect 35675 14459 35681 14493
rect 35681 14459 35719 14493
rect 35719 14459 35727 14493
rect 35742 14459 35753 14493
rect 35753 14459 35791 14493
rect 35791 14459 35794 14493
rect 35809 14459 35825 14493
rect 35825 14459 35861 14493
rect 35877 14459 35897 14493
rect 35897 14459 35929 14493
rect 35945 14459 35969 14493
rect 35969 14459 35997 14493
rect 36013 14459 36041 14493
rect 36041 14459 36065 14493
rect 36081 14459 36113 14493
rect 36113 14459 36133 14493
rect 35675 14450 35727 14459
rect 35742 14450 35794 14459
rect 35809 14450 35861 14459
rect 35877 14450 35929 14459
rect 35945 14450 35997 14459
rect 36013 14450 36065 14459
rect 36081 14450 36133 14459
rect 36149 14493 36201 14502
rect 36149 14459 36151 14493
rect 36151 14459 36185 14493
rect 36185 14459 36201 14493
rect 36149 14450 36201 14459
rect 36217 14493 36269 14502
rect 36217 14459 36223 14493
rect 36223 14459 36257 14493
rect 36257 14459 36269 14493
rect 36217 14450 36269 14459
rect 36285 14493 36337 14502
rect 36285 14459 36295 14493
rect 36295 14459 36329 14493
rect 36329 14459 36337 14493
rect 36285 14450 36337 14459
rect 36353 14493 36405 14502
rect 36353 14459 36367 14493
rect 36367 14459 36401 14493
rect 36401 14459 36405 14493
rect 36353 14450 36405 14459
rect 36421 14493 36473 14502
rect 36421 14459 36439 14493
rect 36439 14459 36473 14493
rect 36421 14450 36473 14459
rect 36489 14493 36541 14502
rect 36489 14459 36511 14493
rect 36511 14459 36541 14493
rect 36489 14450 36541 14459
rect 37618 14497 37670 14515
rect 37618 14476 37670 14484
rect 37618 14442 37627 14476
rect 37627 14442 37661 14476
rect 37661 14442 37670 14476
rect 37618 14432 37670 14442
rect 37618 14403 37670 14419
rect 37618 14369 37627 14403
rect 37627 14369 37661 14403
rect 37661 14369 37670 14403
rect 37618 14367 37670 14369
rect 36667 14337 36719 14346
rect 36732 14337 36784 14346
rect 36667 14303 36689 14337
rect 36689 14303 36719 14337
rect 36732 14303 36761 14337
rect 36761 14303 36784 14337
rect 36667 14294 36719 14303
rect 36732 14294 36784 14303
rect 36797 14337 36849 14346
rect 36797 14303 36799 14337
rect 36799 14303 36833 14337
rect 36833 14303 36849 14337
rect 36797 14294 36849 14303
rect 36862 14337 36914 14346
rect 36862 14303 36871 14337
rect 36871 14303 36905 14337
rect 36905 14303 36914 14337
rect 36862 14294 36914 14303
rect 36927 14337 36979 14346
rect 36927 14303 36943 14337
rect 36943 14303 36977 14337
rect 36977 14303 36979 14337
rect 36927 14294 36979 14303
rect 36992 14337 37044 14346
rect 37057 14337 37109 14346
rect 37122 14337 37174 14346
rect 37188 14337 37240 14346
rect 37254 14337 37306 14346
rect 37320 14337 37372 14346
rect 37386 14337 37438 14346
rect 37452 14337 37504 14346
rect 36992 14303 37015 14337
rect 37015 14303 37044 14337
rect 37057 14303 37087 14337
rect 37087 14303 37109 14337
rect 37122 14303 37159 14337
rect 37159 14303 37174 14337
rect 37188 14303 37193 14337
rect 37193 14303 37231 14337
rect 37231 14303 37240 14337
rect 37254 14303 37265 14337
rect 37265 14303 37303 14337
rect 37303 14303 37306 14337
rect 37320 14303 37337 14337
rect 37337 14303 37372 14337
rect 37386 14303 37409 14337
rect 37409 14303 37438 14337
rect 37452 14303 37481 14337
rect 37481 14303 37504 14337
rect 36992 14294 37044 14303
rect 37057 14294 37109 14303
rect 37122 14294 37174 14303
rect 37188 14294 37240 14303
rect 37254 14294 37306 14303
rect 37320 14294 37372 14303
rect 37386 14294 37438 14303
rect 37452 14294 37504 14303
rect 37618 14330 37670 14354
rect 37618 14302 37627 14330
rect 37627 14302 37661 14330
rect 37661 14302 37670 14330
rect 37618 14257 37670 14289
rect 37618 14237 37627 14257
rect 37627 14237 37661 14257
rect 37661 14237 37670 14257
rect 37618 14223 37627 14224
rect 37627 14223 37661 14224
rect 37661 14223 37670 14224
rect 35675 14181 35727 14190
rect 35742 14181 35794 14190
rect 35809 14181 35861 14190
rect 35877 14181 35929 14190
rect 35945 14181 35997 14190
rect 36013 14181 36065 14190
rect 36081 14181 36133 14190
rect 35675 14147 35681 14181
rect 35681 14147 35719 14181
rect 35719 14147 35727 14181
rect 35742 14147 35753 14181
rect 35753 14147 35791 14181
rect 35791 14147 35794 14181
rect 35809 14147 35825 14181
rect 35825 14147 35861 14181
rect 35877 14147 35897 14181
rect 35897 14147 35929 14181
rect 35945 14147 35969 14181
rect 35969 14147 35997 14181
rect 36013 14147 36041 14181
rect 36041 14147 36065 14181
rect 36081 14147 36113 14181
rect 36113 14147 36133 14181
rect 35675 14138 35727 14147
rect 35742 14138 35794 14147
rect 35809 14138 35861 14147
rect 35877 14138 35929 14147
rect 35945 14138 35997 14147
rect 36013 14138 36065 14147
rect 36081 14138 36133 14147
rect 36149 14181 36201 14190
rect 36149 14147 36151 14181
rect 36151 14147 36185 14181
rect 36185 14147 36201 14181
rect 36149 14138 36201 14147
rect 36217 14181 36269 14190
rect 36217 14147 36223 14181
rect 36223 14147 36257 14181
rect 36257 14147 36269 14181
rect 36217 14138 36269 14147
rect 36285 14181 36337 14190
rect 36285 14147 36295 14181
rect 36295 14147 36329 14181
rect 36329 14147 36337 14181
rect 36285 14138 36337 14147
rect 36353 14181 36405 14190
rect 36353 14147 36367 14181
rect 36367 14147 36401 14181
rect 36401 14147 36405 14181
rect 36353 14138 36405 14147
rect 36421 14181 36473 14190
rect 36421 14147 36439 14181
rect 36439 14147 36473 14181
rect 36421 14138 36473 14147
rect 36489 14181 36541 14190
rect 36489 14147 36511 14181
rect 36511 14147 36541 14181
rect 36489 14138 36541 14147
rect 37618 14184 37670 14223
rect 37618 14172 37627 14184
rect 37627 14172 37661 14184
rect 37661 14172 37670 14184
rect 37618 14150 37627 14159
rect 37627 14150 37661 14159
rect 37661 14150 37670 14159
rect 37618 14111 37670 14150
rect 37618 14107 37627 14111
rect 37627 14107 37661 14111
rect 37661 14107 37670 14111
rect 37618 14077 37627 14094
rect 37627 14077 37661 14094
rect 37661 14077 37670 14094
rect 37618 14042 37670 14077
rect 36667 14025 36719 14034
rect 36732 14025 36784 14034
rect 36667 13991 36689 14025
rect 36689 13991 36719 14025
rect 36732 13991 36761 14025
rect 36761 13991 36784 14025
rect 36667 13982 36719 13991
rect 36732 13982 36784 13991
rect 36797 14025 36849 14034
rect 36797 13991 36799 14025
rect 36799 13991 36833 14025
rect 36833 13991 36849 14025
rect 36797 13982 36849 13991
rect 36862 14025 36914 14034
rect 36862 13991 36871 14025
rect 36871 13991 36905 14025
rect 36905 13991 36914 14025
rect 36862 13982 36914 13991
rect 36927 14025 36979 14034
rect 36927 13991 36943 14025
rect 36943 13991 36977 14025
rect 36977 13991 36979 14025
rect 36927 13982 36979 13991
rect 36992 14025 37044 14034
rect 37057 14025 37109 14034
rect 37122 14025 37174 14034
rect 37188 14025 37240 14034
rect 37254 14025 37306 14034
rect 37320 14025 37372 14034
rect 37386 14025 37438 14034
rect 37452 14025 37504 14034
rect 36992 13991 37015 14025
rect 37015 13991 37044 14025
rect 37057 13991 37087 14025
rect 37087 13991 37109 14025
rect 37122 13991 37159 14025
rect 37159 13991 37174 14025
rect 37188 13991 37193 14025
rect 37193 13991 37231 14025
rect 37231 13991 37240 14025
rect 37254 13991 37265 14025
rect 37265 13991 37303 14025
rect 37303 13991 37306 14025
rect 37320 13991 37337 14025
rect 37337 13991 37372 14025
rect 37386 13991 37409 14025
rect 37409 13991 37438 14025
rect 37452 13991 37481 14025
rect 37481 13991 37504 14025
rect 36992 13982 37044 13991
rect 37057 13982 37109 13991
rect 37122 13982 37174 13991
rect 37188 13982 37240 13991
rect 37254 13982 37306 13991
rect 37320 13982 37372 13991
rect 37386 13982 37438 13991
rect 37452 13982 37504 13991
rect 37618 14004 37627 14029
rect 37627 14004 37661 14029
rect 37661 14004 37670 14029
rect 37618 13977 37670 14004
rect 37618 13931 37627 13964
rect 37627 13931 37661 13964
rect 37661 13931 37670 13964
rect 37618 13912 37670 13931
rect 37618 13892 37670 13899
rect 35675 13869 35727 13878
rect 35742 13869 35794 13878
rect 35809 13869 35861 13878
rect 35877 13869 35929 13878
rect 35945 13869 35997 13878
rect 36013 13869 36065 13878
rect 36081 13869 36133 13878
rect 35675 13835 35681 13869
rect 35681 13835 35719 13869
rect 35719 13835 35727 13869
rect 35742 13835 35753 13869
rect 35753 13835 35791 13869
rect 35791 13835 35794 13869
rect 35809 13835 35825 13869
rect 35825 13835 35861 13869
rect 35877 13835 35897 13869
rect 35897 13835 35929 13869
rect 35945 13835 35969 13869
rect 35969 13835 35997 13869
rect 36013 13835 36041 13869
rect 36041 13835 36065 13869
rect 36081 13835 36113 13869
rect 36113 13835 36133 13869
rect 35675 13826 35727 13835
rect 35742 13826 35794 13835
rect 35809 13826 35861 13835
rect 35877 13826 35929 13835
rect 35945 13826 35997 13835
rect 36013 13826 36065 13835
rect 36081 13826 36133 13835
rect 36149 13869 36201 13878
rect 36149 13835 36151 13869
rect 36151 13835 36185 13869
rect 36185 13835 36201 13869
rect 36149 13826 36201 13835
rect 36217 13869 36269 13878
rect 36217 13835 36223 13869
rect 36223 13835 36257 13869
rect 36257 13835 36269 13869
rect 36217 13826 36269 13835
rect 36285 13869 36337 13878
rect 36285 13835 36295 13869
rect 36295 13835 36329 13869
rect 36329 13835 36337 13869
rect 36285 13826 36337 13835
rect 36353 13869 36405 13878
rect 36353 13835 36367 13869
rect 36367 13835 36401 13869
rect 36401 13835 36405 13869
rect 36353 13826 36405 13835
rect 36421 13869 36473 13878
rect 36421 13835 36439 13869
rect 36439 13835 36473 13869
rect 36421 13826 36473 13835
rect 36489 13869 36541 13878
rect 36489 13835 36511 13869
rect 36511 13835 36541 13869
rect 36489 13826 36541 13835
rect 37618 13858 37627 13892
rect 37627 13858 37661 13892
rect 37661 13858 37670 13892
rect 37618 13847 37670 13858
rect 37618 13819 37670 13834
rect 37618 13785 37627 13819
rect 37627 13785 37661 13819
rect 37661 13785 37670 13819
rect 37618 13782 37670 13785
rect 37618 13746 37670 13769
rect 36667 13713 36719 13722
rect 36732 13713 36784 13722
rect 36667 13679 36689 13713
rect 36689 13679 36719 13713
rect 36732 13679 36761 13713
rect 36761 13679 36784 13713
rect 36667 13670 36719 13679
rect 36732 13670 36784 13679
rect 36797 13713 36849 13722
rect 36797 13679 36799 13713
rect 36799 13679 36833 13713
rect 36833 13679 36849 13713
rect 36797 13670 36849 13679
rect 36862 13713 36914 13722
rect 36862 13679 36871 13713
rect 36871 13679 36905 13713
rect 36905 13679 36914 13713
rect 36862 13670 36914 13679
rect 36927 13713 36979 13722
rect 36927 13679 36943 13713
rect 36943 13679 36977 13713
rect 36977 13679 36979 13713
rect 36927 13670 36979 13679
rect 36992 13713 37044 13722
rect 37057 13713 37109 13722
rect 37122 13713 37174 13722
rect 37188 13713 37240 13722
rect 37254 13713 37306 13722
rect 37320 13713 37372 13722
rect 37386 13713 37438 13722
rect 37452 13713 37504 13722
rect 36992 13679 37015 13713
rect 37015 13679 37044 13713
rect 37057 13679 37087 13713
rect 37087 13679 37109 13713
rect 37122 13679 37159 13713
rect 37159 13679 37174 13713
rect 37188 13679 37193 13713
rect 37193 13679 37231 13713
rect 37231 13679 37240 13713
rect 37254 13679 37265 13713
rect 37265 13679 37303 13713
rect 37303 13679 37306 13713
rect 37320 13679 37337 13713
rect 37337 13679 37372 13713
rect 37386 13679 37409 13713
rect 37409 13679 37438 13713
rect 37452 13679 37481 13713
rect 37481 13679 37504 13713
rect 36992 13670 37044 13679
rect 37057 13670 37109 13679
rect 37122 13670 37174 13679
rect 37188 13670 37240 13679
rect 37254 13670 37306 13679
rect 37320 13670 37372 13679
rect 37386 13670 37438 13679
rect 37452 13670 37504 13679
rect 37618 13717 37627 13746
rect 37627 13717 37661 13746
rect 37661 13717 37670 13746
rect 37618 13672 37670 13704
rect 37618 13652 37627 13672
rect 37627 13652 37661 13672
rect 37661 13652 37670 13672
rect 37618 13638 37627 13639
rect 37627 13638 37661 13639
rect 37661 13638 37670 13639
rect 37618 13598 37670 13638
rect 37618 13587 37627 13598
rect 37627 13587 37661 13598
rect 37661 13587 37670 13598
rect 35675 13557 35727 13566
rect 35742 13557 35794 13566
rect 35809 13557 35861 13566
rect 35877 13557 35929 13566
rect 35945 13557 35997 13566
rect 36013 13557 36065 13566
rect 36081 13557 36133 13566
rect 35675 13523 35681 13557
rect 35681 13523 35719 13557
rect 35719 13523 35727 13557
rect 35742 13523 35753 13557
rect 35753 13523 35791 13557
rect 35791 13523 35794 13557
rect 35809 13523 35825 13557
rect 35825 13523 35861 13557
rect 35877 13523 35897 13557
rect 35897 13523 35929 13557
rect 35945 13523 35969 13557
rect 35969 13523 35997 13557
rect 36013 13523 36041 13557
rect 36041 13523 36065 13557
rect 36081 13523 36113 13557
rect 36113 13523 36133 13557
rect 35675 13514 35727 13523
rect 35742 13514 35794 13523
rect 35809 13514 35861 13523
rect 35877 13514 35929 13523
rect 35945 13514 35997 13523
rect 36013 13514 36065 13523
rect 36081 13514 36133 13523
rect 36149 13557 36201 13566
rect 36149 13523 36151 13557
rect 36151 13523 36185 13557
rect 36185 13523 36201 13557
rect 36149 13514 36201 13523
rect 36217 13557 36269 13566
rect 36217 13523 36223 13557
rect 36223 13523 36257 13557
rect 36257 13523 36269 13557
rect 36217 13514 36269 13523
rect 36285 13557 36337 13566
rect 36285 13523 36295 13557
rect 36295 13523 36329 13557
rect 36329 13523 36337 13557
rect 36285 13514 36337 13523
rect 36353 13557 36405 13566
rect 36353 13523 36367 13557
rect 36367 13523 36401 13557
rect 36401 13523 36405 13557
rect 36353 13514 36405 13523
rect 36421 13557 36473 13566
rect 36421 13523 36439 13557
rect 36439 13523 36473 13557
rect 36421 13514 36473 13523
rect 36489 13557 36541 13566
rect 37618 13564 37627 13574
rect 37627 13564 37661 13574
rect 37661 13564 37670 13574
rect 36489 13523 36511 13557
rect 36511 13523 36541 13557
rect 36489 13514 36541 13523
rect 37618 13524 37670 13564
rect 37618 13522 37627 13524
rect 37627 13522 37661 13524
rect 37661 13522 37670 13524
rect 37618 13490 37627 13509
rect 37627 13490 37661 13509
rect 37661 13490 37670 13509
rect 37618 13457 37670 13490
rect 36667 13401 36719 13410
rect 36732 13401 36784 13410
rect 36667 13367 36689 13401
rect 36689 13367 36719 13401
rect 36732 13367 36761 13401
rect 36761 13367 36784 13401
rect 36667 13358 36719 13367
rect 36732 13358 36784 13367
rect 36797 13401 36849 13410
rect 36797 13367 36799 13401
rect 36799 13367 36833 13401
rect 36833 13367 36849 13401
rect 36797 13358 36849 13367
rect 36862 13401 36914 13410
rect 36862 13367 36871 13401
rect 36871 13367 36905 13401
rect 36905 13367 36914 13401
rect 36862 13358 36914 13367
rect 36927 13401 36979 13410
rect 36927 13367 36943 13401
rect 36943 13367 36977 13401
rect 36977 13367 36979 13401
rect 36927 13358 36979 13367
rect 36992 13401 37044 13410
rect 37057 13401 37109 13410
rect 37122 13401 37174 13410
rect 37188 13401 37240 13410
rect 37254 13401 37306 13410
rect 37320 13401 37372 13410
rect 37386 13401 37438 13410
rect 37452 13401 37504 13410
rect 36992 13367 37015 13401
rect 37015 13367 37044 13401
rect 37057 13367 37087 13401
rect 37087 13367 37109 13401
rect 37122 13367 37159 13401
rect 37159 13367 37174 13401
rect 37188 13367 37193 13401
rect 37193 13367 37231 13401
rect 37231 13367 37240 13401
rect 37254 13367 37265 13401
rect 37265 13367 37303 13401
rect 37303 13367 37306 13401
rect 37320 13367 37337 13401
rect 37337 13367 37372 13401
rect 37386 13367 37409 13401
rect 37409 13367 37438 13401
rect 37452 13367 37481 13401
rect 37481 13367 37504 13401
rect 36992 13358 37044 13367
rect 37057 13358 37109 13367
rect 37122 13358 37174 13367
rect 37188 13358 37240 13367
rect 37254 13358 37306 13367
rect 37320 13358 37372 13367
rect 37386 13358 37438 13367
rect 37452 13358 37504 13367
rect 37618 13416 37627 13444
rect 37627 13416 37661 13444
rect 37661 13416 37670 13444
rect 37618 13392 37670 13416
rect 37618 13376 37670 13379
rect 37618 13342 37627 13376
rect 37627 13342 37661 13376
rect 37661 13342 37670 13376
rect 37618 13327 37670 13342
rect 37618 13302 37670 13314
rect 37618 13268 37627 13302
rect 37627 13268 37661 13302
rect 37661 13268 37670 13302
rect 37618 13262 37670 13268
rect 35675 13245 35727 13254
rect 35742 13245 35794 13254
rect 35809 13245 35861 13254
rect 35877 13245 35929 13254
rect 35945 13245 35997 13254
rect 36013 13245 36065 13254
rect 36081 13245 36133 13254
rect 35675 13211 35681 13245
rect 35681 13211 35719 13245
rect 35719 13211 35727 13245
rect 35742 13211 35753 13245
rect 35753 13211 35791 13245
rect 35791 13211 35794 13245
rect 35809 13211 35825 13245
rect 35825 13211 35861 13245
rect 35877 13211 35897 13245
rect 35897 13211 35929 13245
rect 35945 13211 35969 13245
rect 35969 13211 35997 13245
rect 36013 13211 36041 13245
rect 36041 13211 36065 13245
rect 36081 13211 36113 13245
rect 36113 13211 36133 13245
rect 35675 13202 35727 13211
rect 35742 13202 35794 13211
rect 35809 13202 35861 13211
rect 35877 13202 35929 13211
rect 35945 13202 35997 13211
rect 36013 13202 36065 13211
rect 36081 13202 36133 13211
rect 36149 13245 36201 13254
rect 36149 13211 36151 13245
rect 36151 13211 36185 13245
rect 36185 13211 36201 13245
rect 36149 13202 36201 13211
rect 36217 13245 36269 13254
rect 36217 13211 36223 13245
rect 36223 13211 36257 13245
rect 36257 13211 36269 13245
rect 36217 13202 36269 13211
rect 36285 13245 36337 13254
rect 36285 13211 36295 13245
rect 36295 13211 36329 13245
rect 36329 13211 36337 13245
rect 36285 13202 36337 13211
rect 36353 13245 36405 13254
rect 36353 13211 36367 13245
rect 36367 13211 36401 13245
rect 36401 13211 36405 13245
rect 36353 13202 36405 13211
rect 36421 13245 36473 13254
rect 36421 13211 36439 13245
rect 36439 13211 36473 13245
rect 36421 13202 36473 13211
rect 36489 13245 36541 13254
rect 36489 13211 36511 13245
rect 36511 13211 36541 13245
rect 36489 13202 36541 13211
rect 17637 3351 17689 3403
rect 17701 3351 17753 3403
rect 17917 3351 17969 3403
rect 17981 3351 18033 3403
rect 17658 3271 17710 3323
rect 17722 3271 17774 3323
rect 18157 3265 18209 3317
rect 18157 3201 18209 3253
rect 19678 2294 19730 2303
rect 19678 2260 19682 2294
rect 19682 2260 19716 2294
rect 19716 2260 19730 2294
rect 19678 2251 19730 2260
rect 19742 2294 19794 2303
rect 19742 2260 19754 2294
rect 19754 2260 19788 2294
rect 19788 2260 19794 2294
rect 19742 2251 19794 2260
rect 23083 2242 23135 2294
rect 23155 2242 23207 2294
rect 23227 2242 23279 2294
rect 23299 2242 23351 2294
rect 23371 2242 23423 2294
rect 23442 2242 23494 2294
rect 23513 2242 23565 2294
rect 23584 2242 23636 2294
rect 17779 2016 17831 2068
rect 17843 2016 17895 2068
rect 20428 2148 20480 2157
rect 20428 2114 20434 2148
rect 20434 2114 20468 2148
rect 20468 2114 20480 2148
rect 20428 2105 20480 2114
rect 20492 2148 20544 2157
rect 20492 2114 20507 2148
rect 20507 2114 20541 2148
rect 20541 2114 20544 2148
rect 20492 2105 20544 2114
rect 17915 1935 17967 1987
rect 17979 1935 18031 1987
rect 20400 1657 20426 1679
rect 20426 1657 20452 1679
rect 20467 1657 20498 1679
rect 20498 1657 20519 1679
rect 20400 1627 20452 1657
rect 20467 1627 20519 1657
rect 20534 1657 20536 1679
rect 20536 1657 20570 1679
rect 20570 1657 20586 1679
rect 20534 1627 20586 1657
rect 20600 1657 20608 1679
rect 20608 1657 20642 1679
rect 20642 1657 20652 1679
rect 20600 1627 20652 1657
rect 20666 1657 20680 1679
rect 20680 1657 20714 1679
rect 20714 1657 20718 1679
rect 20666 1627 20718 1657
rect 20953 1658 20977 1679
rect 20977 1658 21005 1679
rect 21017 1658 21051 1679
rect 21051 1658 21069 1679
rect 20953 1627 21005 1658
rect 21017 1627 21069 1658
<< metal2 >>
rect 37686 16157 37770 16163
rect 37686 16105 37702 16157
rect 37754 16105 37770 16157
rect 37686 16093 37770 16105
rect 37686 16041 37702 16093
rect 37754 16041 37770 16093
rect 37686 16029 37770 16041
rect 37686 15977 37702 16029
rect 37754 15977 37770 16029
rect 37686 15971 37770 15977
tri 37700 15962 37709 15971 ne
tri 37692 15412 37709 15429 se
rect 37709 15412 37754 15971
tri 37621 15341 37692 15412 se
rect 37692 15403 37754 15412
tri 37692 15341 37754 15403 nw
rect 35669 15126 36547 15153
rect 35669 15074 35675 15126
rect 35727 15074 35742 15126
rect 35794 15074 35809 15126
rect 35861 15074 35877 15126
rect 35929 15074 35945 15126
rect 35997 15074 36013 15126
rect 36065 15074 36081 15126
rect 36133 15074 36149 15126
rect 36201 15074 36217 15126
rect 36269 15074 36285 15126
rect 36337 15074 36353 15126
rect 36405 15074 36421 15126
rect 36473 15074 36489 15126
rect 36541 15074 36547 15126
rect 35669 14814 36547 15074
rect 37621 15072 37673 15341
tri 37673 15322 37692 15341 nw
rect 37618 15066 37670 15072
rect 37618 15002 37670 15014
rect 35669 14762 35675 14814
rect 35727 14762 35742 14814
rect 35794 14762 35809 14814
rect 35861 14762 35877 14814
rect 35929 14762 35945 14814
rect 35997 14762 36013 14814
rect 36065 14762 36081 14814
rect 36133 14762 36149 14814
rect 36201 14762 36217 14814
rect 36269 14762 36285 14814
rect 36337 14762 36353 14814
rect 36405 14762 36421 14814
rect 36473 14762 36489 14814
rect 36541 14762 36547 14814
rect 35669 14502 36547 14762
rect 35669 14450 35675 14502
rect 35727 14450 35742 14502
rect 35794 14450 35809 14502
rect 35861 14450 35877 14502
rect 35929 14450 35945 14502
rect 35997 14450 36013 14502
rect 36065 14450 36081 14502
rect 36133 14450 36149 14502
rect 36201 14450 36217 14502
rect 36269 14450 36285 14502
rect 36337 14450 36353 14502
rect 36405 14450 36421 14502
rect 36473 14450 36489 14502
rect 36541 14450 36547 14502
rect 35669 14190 36547 14450
rect 35669 14138 35675 14190
rect 35727 14138 35742 14190
rect 35794 14138 35809 14190
rect 35861 14138 35877 14190
rect 35929 14138 35945 14190
rect 35997 14138 36013 14190
rect 36065 14138 36081 14190
rect 36133 14138 36149 14190
rect 36201 14138 36217 14190
rect 36269 14138 36285 14190
rect 36337 14138 36353 14190
rect 36405 14138 36421 14190
rect 36473 14138 36489 14190
rect 36541 14138 36547 14190
tri 35628 13982 35669 14023 se
rect 35669 13982 36547 14138
tri 35623 13977 35628 13982 se
rect 35628 13977 36547 13982
tri 35610 13964 35623 13977 se
rect 35623 13964 36547 13977
tri 35558 13912 35610 13964 se
rect 35610 13912 36547 13964
tri 35545 13899 35558 13912 se
rect 35558 13899 36547 13912
tri 35524 13878 35545 13899 se
rect 35545 13878 36547 13899
tri 35472 13826 35524 13878 se
rect 35524 13826 35675 13878
rect 35727 13826 35742 13878
rect 35794 13826 35809 13878
rect 35861 13826 35877 13878
rect 35929 13826 35945 13878
rect 35997 13826 36013 13878
rect 36065 13826 36081 13878
rect 36133 13826 36149 13878
rect 36201 13826 36217 13878
rect 36269 13826 36285 13878
rect 36337 13826 36353 13878
rect 36405 13826 36421 13878
rect 36473 13826 36489 13878
rect 36541 13826 36547 13878
tri 35428 13782 35472 13826 se
rect 35472 13782 36547 13826
tri 35415 13769 35428 13782 se
rect 35428 13769 36547 13782
tri 35368 13722 35415 13769 se
rect 35415 13722 36547 13769
tri 35344 13698 35368 13722 se
rect 35368 13698 36547 13722
rect 31824 13694 36547 13698
rect 31820 13638 31829 13694
rect 31885 13638 31911 13694
rect 31967 13638 31993 13694
rect 32049 13638 32075 13694
rect 32131 13638 32157 13694
rect 32213 13638 32239 13694
rect 32295 13638 32321 13694
rect 32377 13638 32403 13694
rect 32459 13638 32486 13694
rect 32542 13638 32569 13694
rect 32625 13638 32652 13694
rect 32708 13638 36547 13694
rect 31820 13566 36547 13638
rect 31820 13560 35675 13566
rect 31820 13504 31829 13560
rect 31885 13504 31911 13560
rect 31967 13504 31993 13560
rect 32049 13504 32075 13560
rect 32131 13504 32157 13560
rect 32213 13504 32239 13560
rect 32295 13504 32321 13560
rect 32377 13504 32403 13560
rect 32459 13504 32486 13560
rect 32542 13504 32569 13560
rect 32625 13504 32652 13560
rect 32708 13514 35675 13560
rect 35727 13514 35742 13566
rect 35794 13514 35809 13566
rect 35861 13514 35877 13566
rect 35929 13514 35945 13566
rect 35997 13514 36013 13566
rect 36065 13514 36081 13566
rect 36133 13514 36149 13566
rect 36201 13514 36217 13566
rect 36269 13514 36285 13566
rect 36337 13514 36353 13566
rect 36405 13514 36421 13566
rect 36473 13514 36489 13566
rect 36541 13514 36547 13566
rect 32708 13504 36547 13514
rect 31824 13500 36547 13504
tri 35356 13457 35399 13500 ne
rect 35399 13457 36547 13500
tri 35399 13444 35412 13457 ne
rect 35412 13444 36547 13457
tri 35412 13410 35446 13444 ne
rect 35446 13410 36547 13444
tri 35446 13358 35498 13410 ne
rect 35498 13358 36547 13410
tri 35498 13327 35529 13358 ne
rect 35529 13327 36547 13358
rect 36661 14918 36667 14970
rect 36719 14918 36732 14970
rect 36784 14918 36797 14970
rect 36849 14918 36862 14970
rect 36914 14918 36927 14970
rect 36979 14918 36992 14970
rect 37044 14918 37057 14970
rect 37109 14918 37122 14970
rect 37174 14918 37188 14970
rect 37240 14918 37254 14970
rect 37306 14918 37320 14970
rect 37372 14918 37386 14970
rect 37438 14918 37452 14970
rect 37504 14918 37510 14970
rect 36661 14658 37510 14918
rect 36661 14606 36667 14658
rect 36719 14606 36732 14658
rect 36784 14606 36797 14658
rect 36849 14606 36862 14658
rect 36914 14606 36927 14658
rect 36979 14606 36992 14658
rect 37044 14606 37057 14658
rect 37109 14606 37122 14658
rect 37174 14606 37188 14658
rect 37240 14606 37254 14658
rect 37306 14606 37320 14658
rect 37372 14606 37386 14658
rect 37438 14606 37452 14658
rect 37504 14606 37510 14658
rect 36661 14346 37510 14606
rect 36661 14294 36667 14346
rect 36719 14294 36732 14346
rect 36784 14294 36797 14346
rect 36849 14294 36862 14346
rect 36914 14294 36927 14346
rect 36979 14294 36992 14346
rect 37044 14294 37057 14346
rect 37109 14294 37122 14346
rect 37174 14294 37188 14346
rect 37240 14294 37254 14346
rect 37306 14294 37320 14346
rect 37372 14294 37386 14346
rect 37438 14294 37452 14346
rect 37504 14294 37510 14346
rect 36661 14034 37510 14294
rect 36661 13982 36667 14034
rect 36719 13982 36732 14034
rect 36784 13982 36797 14034
rect 36849 13982 36862 14034
rect 36914 13982 36927 14034
rect 36979 13982 36992 14034
rect 37044 13982 37057 14034
rect 37109 13982 37122 14034
rect 37174 13982 37188 14034
rect 37240 13982 37254 14034
rect 37306 13982 37320 14034
rect 37372 13982 37386 14034
rect 37438 13982 37452 14034
rect 37504 13982 37510 14034
rect 36661 13722 37510 13982
rect 36661 13670 36667 13722
rect 36719 13670 36732 13722
rect 36784 13670 36797 13722
rect 36849 13670 36862 13722
rect 36914 13670 36927 13722
rect 36979 13670 36992 13722
rect 37044 13670 37057 13722
rect 37109 13670 37122 13722
rect 37174 13670 37188 13722
rect 37240 13670 37254 13722
rect 37306 13670 37320 13722
rect 37372 13670 37386 13722
rect 37438 13670 37452 13722
rect 37504 13670 37510 13722
rect 36661 13410 37510 13670
rect 36661 13358 36667 13410
rect 36719 13358 36732 13410
rect 36784 13358 36797 13410
rect 36849 13358 36862 13410
rect 36914 13358 36927 13410
rect 36979 13358 36992 13410
rect 37044 13358 37057 13410
rect 37109 13358 37122 13410
rect 37174 13358 37188 13410
rect 37240 13358 37254 13410
rect 37306 13358 37320 13410
rect 37372 13358 37386 13410
rect 37438 13358 37452 13410
rect 37504 13358 37510 13410
rect 36661 13342 37510 13358
rect 37618 14938 37670 14950
rect 37618 14874 37670 14886
rect 37618 14809 37670 14822
rect 37618 14744 37670 14757
rect 37618 14679 37670 14692
rect 37618 14614 37670 14627
rect 37618 14549 37670 14562
rect 37618 14484 37670 14497
rect 37618 14419 37670 14432
rect 37618 14354 37670 14367
rect 37618 14289 37670 14302
rect 37618 14224 37670 14237
rect 37618 14159 37670 14172
rect 37618 14094 37670 14107
rect 37618 14029 37670 14042
rect 37618 13964 37670 13977
rect 37618 13899 37670 13912
rect 37618 13834 37670 13847
rect 37618 13769 37670 13782
rect 37618 13704 37670 13717
rect 37618 13639 37670 13652
rect 37618 13574 37670 13587
rect 37618 13509 37670 13522
rect 37618 13444 37670 13457
rect 37618 13379 37670 13392
tri 35529 13314 35542 13327 ne
rect 35542 13314 36547 13327
tri 35542 13262 35594 13314 ne
rect 35594 13262 36547 13314
tri 35594 13254 35602 13262 ne
rect 35602 13254 36547 13262
rect 37618 13314 37670 13327
rect 37618 13256 37670 13262
tri 35602 13202 35654 13254 ne
rect 35654 13202 35675 13254
rect 35727 13202 35742 13254
rect 35794 13202 35809 13254
rect 35861 13202 35877 13254
rect 35929 13202 35945 13254
rect 35997 13202 36013 13254
rect 36065 13202 36081 13254
rect 36133 13202 36149 13254
rect 36201 13202 36217 13254
rect 36269 13202 36285 13254
rect 36337 13202 36353 13254
rect 36405 13202 36421 13254
rect 36473 13202 36489 13254
rect 36541 13202 36547 13254
tri 35654 13133 35723 13202 ne
rect 17631 3351 17637 3403
rect 17689 3351 17701 3403
rect 17753 3351 17917 3403
rect 17969 3351 17981 3403
rect 18033 3351 18039 3403
rect 17652 3271 17658 3323
rect 17710 3271 17722 3323
rect 17774 3317 18209 3323
rect 17774 3271 18157 3317
rect 18157 3253 18209 3265
rect 18157 3195 18209 3201
rect 19672 2251 19678 2303
rect 19730 2251 19742 2303
rect 19794 2294 20003 2303
tri 20003 2294 20012 2303 sw
rect 19794 2251 20012 2294
tri 20012 2251 20055 2294 sw
tri 21440 2251 21483 2294 se
rect 21483 2251 23083 2294
tri 19989 2242 19998 2251 ne
rect 19998 2242 20055 2251
tri 20055 2242 20064 2251 sw
tri 21431 2242 21440 2251 se
rect 21440 2242 23083 2251
rect 23135 2242 23155 2294
rect 23207 2242 23227 2294
rect 23279 2242 23299 2294
rect 23351 2242 23371 2294
rect 23423 2242 23442 2294
rect 23494 2242 23513 2294
rect 23565 2242 23584 2294
rect 23636 2242 23647 2294
tri 19998 2185 20055 2242 ne
rect 20055 2185 20064 2242
tri 20064 2185 20121 2242 sw
tri 21409 2220 21431 2242 se
rect 21431 2220 21483 2242
tri 21483 2220 21505 2242 nw
tri 21374 2185 21409 2220 se
tri 20055 2157 20083 2185 ne
rect 20083 2157 20121 2185
tri 20121 2157 20149 2185 sw
tri 21346 2157 21374 2185 se
rect 21374 2157 21409 2185
tri 20083 2119 20121 2157 ne
rect 20121 2119 20428 2157
tri 20121 2105 20135 2119 ne
rect 20135 2105 20428 2119
rect 20480 2105 20492 2157
rect 20544 2105 20550 2157
tri 21335 2146 21346 2157 se
rect 21346 2146 21409 2157
tri 21409 2146 21483 2220 nw
tri 21294 2105 21335 2146 se
tri 21261 2072 21294 2105 se
rect 21294 2072 21335 2105
tri 21335 2072 21409 2146 nw
tri 21257 2068 21261 2072 se
rect 17773 2016 17779 2068
rect 17831 2016 17843 2068
rect 17895 2016 17901 2068
tri 21205 2016 21257 2068 se
rect 21257 2016 21261 2068
tri 21187 1998 21205 2016 se
rect 21205 1998 21261 2016
tri 21261 1998 21335 2072 nw
tri 21176 1987 21187 1998 se
rect 21187 1987 21250 1998
tri 21250 1987 21261 1998 nw
rect 17909 1935 17915 1987
rect 17967 1935 17979 1987
rect 18031 1937 21200 1987
tri 21200 1937 21250 1987 nw
rect 18031 1935 18037 1937
rect 20394 1627 20400 1679
rect 20452 1627 20467 1679
rect 20519 1627 20534 1679
rect 20586 1627 20600 1679
rect 20652 1627 20666 1679
rect 20718 1627 20953 1679
rect 21005 1627 21017 1679
rect 21069 1627 21147 1679
<< via2 >>
rect 31829 13638 31885 13694
rect 31911 13638 31967 13694
rect 31993 13638 32049 13694
rect 32075 13638 32131 13694
rect 32157 13638 32213 13694
rect 32239 13638 32295 13694
rect 32321 13638 32377 13694
rect 32403 13638 32459 13694
rect 32486 13638 32542 13694
rect 32569 13638 32625 13694
rect 32652 13638 32708 13694
rect 31829 13504 31885 13560
rect 31911 13504 31967 13560
rect 31993 13504 32049 13560
rect 32075 13504 32131 13560
rect 32157 13504 32213 13560
rect 32239 13504 32295 13560
rect 32321 13504 32377 13560
rect 32403 13504 32459 13560
rect 32486 13504 32542 13560
rect 32569 13504 32625 13560
rect 32652 13504 32708 13560
<< metal3 >>
rect 31824 13694 32713 13699
rect 31824 13638 31829 13694
rect 31885 13638 31911 13694
rect 31967 13638 31993 13694
rect 32049 13638 32075 13694
rect 32131 13638 32157 13694
rect 32213 13638 32239 13694
rect 32295 13638 32321 13694
rect 32377 13638 32403 13694
rect 32459 13638 32486 13694
rect 32542 13638 32569 13694
rect 32625 13638 32652 13694
rect 32708 13638 32713 13694
rect 31824 13560 32713 13638
rect 31824 13504 31829 13560
rect 31885 13504 31911 13560
rect 31967 13504 31993 13560
rect 32049 13504 32075 13560
rect 32131 13504 32157 13560
rect 32213 13504 32239 13560
rect 32295 13504 32321 13560
rect 32377 13504 32403 13560
rect 32459 13504 32486 13560
rect 32542 13504 32569 13560
rect 32625 13504 32652 13560
rect 32708 13504 32713 13560
rect 31824 13499 32713 13504
use sky130_fd_pr__pfet_01v8__example_55959141808126  sky130_fd_pr__pfet_01v8__example_55959141808126_0
timestamp 1619729480
transform -1 0 13479 0 1 1831
box -28 0 284 267
use sky130_fd_pr__pfet_01v8__example_55959141808126  sky130_fd_pr__pfet_01v8__example_55959141808126_1
timestamp 1619729480
transform -1 0 13791 0 1 1831
box -28 0 284 267
use sky130_fd_pr__pfet_01v8__example_55959141808125  sky130_fd_pr__pfet_01v8__example_55959141808125_0
timestamp 1619729480
transform -1 0 14415 0 1 1831
box -28 0 596 267
use sky130_fd_pr__pfet_01v8__example_55959141808124  sky130_fd_pr__pfet_01v8__example_55959141808124_0
timestamp 1619729480
transform 1 0 12724 0 1 2137
box -28 0 228 29
use sky130_fd_pr__pfet_01v8__example_55959141808124  sky130_fd_pr__pfet_01v8__example_55959141808124_1
timestamp 1619729480
transform -1 0 12668 0 1 2137
box -28 0 228 29
use sky130_fd_pr__pfet_01v8__example_55959141808121  sky130_fd_pr__pfet_01v8__example_55959141808121_0
timestamp 1619729480
transform 1 0 12542 0 -1 1940
box -28 0 428 29
use sky130_fd_pr__pfet_01v8__example_55959141808121  sky130_fd_pr__pfet_01v8__example_55959141808121_1
timestamp 1619729480
transform -1 0 12486 0 -1 1940
box -28 0 428 29
use sky130_fd_pr__pfet_01v8__example_55959141808120  sky130_fd_pr__pfet_01v8__example_55959141808120_0
timestamp 1619729480
transform -1 0 15039 0 1 1831
box -28 0 596 267
use sky130_fd_pr__pfet_01v8__example_55959141808119  sky130_fd_pr__pfet_01v8__example_55959141808119_0
timestamp 1619729480
transform 0 1 35579 1 0 13256
box -28 0 1844 985
use sky130_fd_pr__nfet_01v8__example_55959141808118  sky130_fd_pr__nfet_01v8__example_55959141808118_0
timestamp 1619729480
transform 1 0 13042 0 -1 3566
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_5595914180888  sky130_fd_pr__nfet_01v8__example_5595914180888_0
timestamp 1619729480
transform 1 0 13198 0 -1 3566
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_5595914180888  sky130_fd_pr__nfet_01v8__example_5595914180888_1
timestamp 1619729480
transform 1 0 13510 0 -1 3566
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_5595914180888  sky130_fd_pr__nfet_01v8__example_5595914180888_2
timestamp 1619729480
transform 1 0 14419 0 -1 3566
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_5595914180888  sky130_fd_pr__nfet_01v8__example_5595914180888_3
timestamp 1619729480
transform 1 0 14263 0 -1 3566
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_5595914180888  sky130_fd_pr__nfet_01v8__example_5595914180888_4
timestamp 1619729480
transform 1 0 13354 0 -1 3566
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_55959141808117  sky130_fd_pr__nfet_01v8__example_55959141808117_0
timestamp 1619729480
transform 1 0 12724 0 -1 2492
box -28 0 228 29
use sky130_fd_pr__nfet_01v8__example_55959141808117  sky130_fd_pr__nfet_01v8__example_55959141808117_1
timestamp 1619729480
transform -1 0 12668 0 -1 2492
box -28 0 228 29
use sky130_fd_pr__nfet_01v8__example_55959141808116  sky130_fd_pr__nfet_01v8__example_55959141808116_0
timestamp 1619729480
transform 1 0 14087 0 -1 3566
box -28 0 148 267
use sky130_fd_pr__nfet_01v8__example_55959141808116  sky130_fd_pr__nfet_01v8__example_55959141808116_1
timestamp 1619729480
transform -1 0 13907 0 -1 3566
box -28 0 148 267
use sky130_fd_pr__nfet_01v8__example_55959141808114  sky130_fd_pr__nfet_01v8__example_55959141808114_0
timestamp 1619729480
transform 1 0 12418 0 -1 3566
box -28 0 284 267
use sky130_fd_pr__nfet_01v8__example_55959141808114  sky130_fd_pr__nfet_01v8__example_55959141808114_1
timestamp 1619729480
transform 1 0 11794 0 -1 3566
box -28 0 284 267
use sky130_fd_pr__nfet_01v8__example_55959141808114  sky130_fd_pr__nfet_01v8__example_55959141808114_2
timestamp 1619729480
transform 1 0 12730 0 -1 3566
box -28 0 284 267
use sky130_fd_pr__nfet_01v8__example_55959141808114  sky130_fd_pr__nfet_01v8__example_55959141808114_3
timestamp 1619729480
transform 1 0 12106 0 -1 3566
box -28 0 284 267
use sky130_fd_io__sio_hotswap_hys  sky130_fd_io__sio_hotswap_hys_0
timestamp 1619729480
transform -1 0 16518 0 -1 2448
box 0 -76 1215 674
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_0
timestamp 1619729480
transform 0 1 16629 1 0 2280
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_1
timestamp 1619729480
transform 0 1 16629 -1 0 2280
box -107 21 267 1369
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_0
timestamp 1619729480
transform 1 0 17335 0 -1 2563
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_0
timestamp 1619729480
transform 1 0 17735 0 1 2433
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180896  sky130_fd_io__tk_em1s_cdns_5595914180896_0
timestamp 1619729480
transform 1 0 16576 0 1 2027
box 0 24 144 28
use sky130_fd_io__sio_hotswap_wpd_ovtv2  sky130_fd_io__sio_hotswap_wpd_ovtv2_0
timestamp 1619729480
transform 1 0 18201 0 1 1641
box 32 52 1830 1178
use sky130_fd_io__sio_hotswap_wpd_ovtv2_1  sky130_fd_io__sio_hotswap_wpd_ovtv2_1_0
timestamp 1619729480
transform 1 0 20285 0 -1 2186
box -150 -571 3405 495
use sky130_fd_io__gpio_ovtv2_hotswap_pghspd  sky130_fd_io__gpio_ovtv2_hotswap_pghspd_0
timestamp 1619729480
transform 1 0 14575 0 -1 3623
box 65 -57 3367 835
<< labels >>
flabel metal2 s 35954 14244 36173 14437 3 FreeSans 520 0 0 0 VCC_IO
flabel metal1 s 14753 2474 14811 2516 0 FreeSans 400 0 0 0 PAD_ESD
flabel metal1 s 19011 2257 19069 2299 0 FreeSans 440 0 0 0 VPWR_KA
flabel metal1 s 14291 2844 14349 2886 0 FreeSans 440 0 0 0 ENHS_H
flabel metal1 s 12079 2880 12137 2922 0 FreeSans 440 0 0 0 EXITHS_H
flabel metal1 s 13283 2880 13341 2922 0 FreeSans 440 0 0 0 ENHS_H_N
flabel metal1 s 12690 2880 12748 2922 0 FreeSans 440 0 0 0 DISHS_H
flabel metal1 s 14111 2474 14169 2516 0 FreeSans 440 180 0 0 DISHS_H_N
flabel metal1 s 12460 2480 12693 2595 3 FreeSans 520 0 0 0 VGND
flabel metal1 s 17102 2590 17180 2642 3 FreeSans 520 0 0 0 ENHS_LATHYS_H_N
flabel metal1 s 18012 2517 18062 2563 3 FreeSans 520 0 0 0 ENHS_LAT_H_N
flabel metal1 s 14672 3518 14905 3649 3 FreeSans 520 0 0 0 VGND
flabel metal1 s 14199 1792 14418 1985 3 FreeSans 520 0 0 0 VCC_IO
flabel metal1 s 12623 3171 12733 3217 3 FreeSans 520 0 0 0 PGHS_H
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 40195864
string GDS_START 40098232
<< end >>
