magic
tech sky130A
magscale 1 2
timestamp 1619729579
<< nwell >>
rect -66 377 3042 897
<< pwell >>
rect 0 -17 2976 17
<< locali >>
rect 121 441 551 504
rect 720 443 839 553
rect 121 371 610 405
rect 121 289 359 371
rect 544 219 610 371
rect 869 235 935 337
rect 2732 439 2804 747
rect 2770 356 2804 439
rect 2770 301 2951 356
rect 2732 123 2804 301
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 2976 831
rect 182 735 372 741
rect 182 701 188 735
rect 222 701 260 735
rect 294 701 332 735
rect 366 701 372 735
rect 25 253 76 685
rect 182 585 372 701
rect 727 735 917 747
rect 727 701 733 735
rect 767 701 805 735
rect 839 701 877 735
rect 911 701 917 735
rect 480 619 546 685
rect 480 585 680 619
rect 727 589 917 701
rect 646 407 680 585
rect 953 553 1019 747
rect 1063 735 1181 747
rect 1063 701 1069 735
rect 1103 701 1141 735
rect 1175 701 1181 735
rect 1063 589 1181 701
rect 1219 701 1285 747
rect 1806 741 1996 751
rect 1806 707 1812 741
rect 1846 707 1884 741
rect 1918 707 1956 741
rect 1990 707 1996 741
rect 1806 701 1996 707
rect 2396 735 2586 747
rect 2396 701 2402 735
rect 2436 701 2474 735
rect 2508 701 2546 735
rect 2580 701 2586 735
rect 1219 667 1465 701
rect 1219 589 1285 667
rect 953 519 1121 553
rect 1055 443 1121 519
rect 1322 539 1395 631
rect 1322 407 1356 539
rect 1431 503 1465 667
rect 2064 665 2290 699
rect 1392 445 1465 503
rect 1501 535 1551 635
rect 1608 631 2098 665
rect 395 253 461 335
rect 25 219 461 253
rect 646 373 1356 407
rect 25 103 91 219
rect 646 183 680 373
rect 1108 265 1174 337
rect 971 231 1174 265
rect 181 113 371 183
rect 181 79 187 113
rect 221 79 259 113
rect 293 79 331 113
rect 365 79 371 113
rect 479 149 680 183
rect 479 99 545 149
rect 716 113 897 199
rect 971 195 1005 231
rect 1313 199 1356 373
rect 181 73 371 79
rect 716 79 718 113
rect 752 79 790 113
rect 824 79 862 113
rect 896 79 897 113
rect 933 103 1005 195
rect 1043 113 1161 195
rect 716 73 897 79
rect 1043 79 1049 113
rect 1083 79 1121 113
rect 1155 79 1161 113
rect 1043 73 1161 79
rect 1199 87 1265 195
rect 1313 123 1379 199
rect 1415 87 1449 445
rect 1501 355 1535 535
rect 1608 499 1642 631
rect 1962 535 2028 595
rect 1576 391 1642 499
rect 1724 425 1790 511
rect 1962 425 1996 535
rect 2064 499 2098 631
rect 2134 535 2215 629
rect 2032 461 2098 499
rect 1724 391 2129 425
rect 1501 321 1937 355
rect 1501 199 1551 321
rect 2009 285 2059 355
rect 1485 123 1551 199
rect 1587 251 2059 285
rect 1587 87 1642 251
rect 2095 215 2129 391
rect 1199 53 1642 87
rect 1736 113 1926 215
rect 1736 79 1742 113
rect 1776 79 1814 113
rect 1848 79 1886 113
rect 1920 79 1926 113
rect 1962 181 2129 215
rect 1962 99 2028 181
rect 2165 133 2215 535
rect 2251 217 2290 665
rect 2396 539 2586 701
rect 2326 469 2586 503
rect 2326 133 2360 469
rect 2396 331 2462 431
rect 2520 369 2586 469
rect 2622 403 2688 747
rect 2840 735 2958 747
rect 2840 701 2846 735
rect 2880 701 2918 735
rect 2952 701 2958 735
rect 2840 439 2958 701
rect 2622 337 2734 403
rect 2622 331 2688 337
rect 2396 297 2688 331
rect 2165 99 2360 133
rect 2396 113 2586 261
rect 1736 73 1926 79
rect 2396 79 2402 113
rect 2436 79 2474 113
rect 2508 79 2546 113
rect 2580 79 2586 113
rect 2622 103 2688 297
rect 2840 113 2958 265
rect 2396 73 2586 79
rect 2840 79 2846 113
rect 2880 79 2918 113
rect 2952 79 2958 113
rect 2840 73 2958 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 188 701 222 735
rect 260 701 294 735
rect 332 701 366 735
rect 733 701 767 735
rect 805 701 839 735
rect 877 701 911 735
rect 1069 701 1103 735
rect 1141 701 1175 735
rect 1812 707 1846 741
rect 1884 707 1918 741
rect 1956 707 1990 741
rect 2402 701 2436 735
rect 2474 701 2508 735
rect 2546 701 2580 735
rect 187 79 221 113
rect 259 79 293 113
rect 331 79 365 113
rect 718 79 752 113
rect 790 79 824 113
rect 862 79 896 113
rect 1049 79 1083 113
rect 1121 79 1155 113
rect 1742 79 1776 113
rect 1814 79 1848 113
rect 1886 79 1920 113
rect 2846 701 2880 735
rect 2918 701 2952 735
rect 2402 79 2436 113
rect 2474 79 2508 113
rect 2546 79 2580 113
rect 2846 79 2880 113
rect 2918 79 2952 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
<< metal1 >>
rect 0 831 2976 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 2976 831
rect 0 791 2976 797
rect 0 741 2976 763
rect 0 735 1812 741
rect 0 701 188 735
rect 222 701 260 735
rect 294 701 332 735
rect 366 701 733 735
rect 767 701 805 735
rect 839 701 877 735
rect 911 701 1069 735
rect 1103 701 1141 735
rect 1175 707 1812 735
rect 1846 707 1884 741
rect 1918 707 1956 741
rect 1990 735 2976 741
rect 1990 707 2402 735
rect 1175 701 2402 707
rect 2436 701 2474 735
rect 2508 701 2546 735
rect 2580 701 2846 735
rect 2880 701 2918 735
rect 2952 701 2976 735
rect 0 689 2976 701
rect 0 113 2976 125
rect 0 79 187 113
rect 221 79 259 113
rect 293 79 331 113
rect 365 79 718 113
rect 752 79 790 113
rect 824 79 862 113
rect 896 79 1049 113
rect 1083 79 1121 113
rect 1155 79 1742 113
rect 1776 79 1814 113
rect 1848 79 1886 113
rect 1920 79 2402 113
rect 2436 79 2474 113
rect 2508 79 2546 113
rect 2580 79 2846 113
rect 2880 79 2918 113
rect 2952 79 2976 113
rect 0 51 2976 79
rect 0 17 2976 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
rect 0 -23 2976 -17
<< labels >>
rlabel locali s 121 441 551 504 6 D
port 2 nsew signal input
rlabel locali s 2770 356 2804 439 6 Q
port 9 nsew signal output
rlabel locali s 2770 301 2951 356 6 Q
port 9 nsew signal output
rlabel locali s 2732 439 2804 747 6 Q
port 9 nsew signal output
rlabel locali s 2732 123 2804 301 6 Q
port 9 nsew signal output
rlabel locali s 720 443 839 553 6 SCD
port 3 nsew signal input
rlabel locali s 544 219 610 371 6 SCE
port 4 nsew signal input
rlabel locali s 121 371 610 405 6 SCE
port 4 nsew signal input
rlabel locali s 121 289 359 371 6 SCE
port 4 nsew signal input
rlabel locali s 869 235 935 337 6 CLK
port 1 nsew clock input
rlabel metal1 s 0 51 2976 125 6 VGND
port 5 nsew ground bidirectional
rlabel pwell s 0 -17 2976 17 8 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 -23 2976 23 8 VNB
port 6 nsew ground bidirectional
rlabel nwell s -66 377 3042 897 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 791 2976 837 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 689 2976 763 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 2976 814
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_END 794358
string GDS_START 765370
<< end >>
