magic
tech sky130A
magscale 1 2
timestamp 1640697980
<< nwell >>
rect -38 261 130 827
rect 384 261 596 827
rect 850 261 1481 827
<< pwell >>
rect 3 893 89 1050
rect 511 885 1111 1067
rect 1383 893 1469 1050
rect 3 38 89 195
rect 601 192 1425 203
rect 398 56 1425 192
rect 601 21 1425 56
<< locali >>
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1472 1105
rect 17 926 75 1071
rect 529 903 581 1071
rect 715 903 753 1071
rect 889 903 991 1071
rect 1397 926 1455 1071
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 378 561
rect 412 532 562 750
rect 412 467 478 532
rect 276 457 478 467
rect 276 423 284 457
rect 318 423 356 457
rect 390 423 428 457
rect 462 423 478 457
rect 276 413 478 423
rect 412 327 478 413
rect 17 17 75 162
rect 404 17 470 179
rect 594 214 658 308
rect 978 561 1024 748
rect 978 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 978 325 1024 527
rect 1072 282 1127 474
rect 1181 322 1215 527
rect 1256 282 1311 474
rect 1351 322 1387 527
rect 1072 217 1311 282
rect 1072 196 1127 217
rect 623 17 689 180
rect 795 17 861 112
rect 967 17 1033 180
rect 1067 51 1127 196
rect 1165 17 1231 169
rect 1267 51 1311 217
rect 1351 17 1401 185
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 1071 63 1105
rect 121 1071 155 1105
rect 213 1071 247 1105
rect 305 1071 339 1105
rect 397 1071 431 1105
rect 489 1071 523 1105
rect 581 1071 615 1105
rect 673 1071 707 1105
rect 765 1071 799 1105
rect 857 1071 891 1105
rect 949 1071 983 1105
rect 1041 1071 1075 1105
rect 1133 1071 1167 1105
rect 1225 1071 1259 1105
rect 1317 1071 1351 1105
rect 1409 1071 1443 1105
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 284 423 318 457
rect 356 423 390 457
rect 428 423 462 457
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< obsli1 >>
rect 615 865 681 1037
rect 787 865 853 1037
rect 1027 964 1097 1032
rect 1027 892 1139 964
rect 1027 881 1153 892
rect 615 853 853 865
rect 1072 871 1153 881
rect 629 831 839 853
rect 17 731 75 794
rect 17 697 28 731
rect 62 697 75 731
rect 17 597 75 697
rect 612 474 678 793
rect 804 762 838 831
rect 1072 825 1217 871
rect 882 728 944 748
rect 736 694 944 728
rect 736 515 770 694
rect 804 583 838 660
rect 878 617 944 694
rect 804 549 928 583
rect 736 481 838 515
rect 512 426 678 474
rect 512 75 560 426
rect 804 196 838 481
rect 894 325 928 549
rect 1072 614 1110 825
rect 1397 731 1455 791
rect 1397 697 1398 731
rect 1432 697 1455 731
rect 1397 597 1455 697
rect 723 146 933 196
rect 723 51 761 146
rect 895 51 933 146
<< obsli1c >>
rect 28 697 62 731
rect 1398 697 1432 731
<< metal1 >>
rect 0 1105 1472 1136
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1317 1105
rect 1351 1071 1409 1105
rect 1443 1071 1472 1105
rect 0 1040 1472 1071
rect 16 731 74 737
rect 16 728 28 731
rect 14 700 28 728
rect 16 697 28 700
rect 62 728 74 731
rect 1386 731 1444 737
rect 1386 728 1398 731
rect 62 700 1398 728
rect 62 697 74 700
rect 16 691 74 697
rect 1386 697 1398 700
rect 1432 728 1444 731
rect 1432 700 1458 728
rect 1432 697 1444 700
rect 1386 691 1444 697
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 272 457 474 463
rect 272 456 284 457
rect 14 428 284 456
rect 272 423 284 428
rect 318 423 356 457
rect 390 423 428 457
rect 462 456 474 457
rect 462 428 1458 456
rect 462 423 474 428
rect 272 417 474 423
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
rlabel locali s 594 214 658 308 6 A
port 1 nsew signal input
rlabel metal1 s 272 417 474 428 6 LOWLVPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 14 428 1458 456 6 LOWLVPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 272 456 474 463 6 LOWLVPWR
port 2 nsew power bidirectional abutment
rlabel nwell s 384 261 596 827 6 LOWLVPWR
port 2 nsew power bidirectional abutment
rlabel viali s 428 423 462 457 6 LOWLVPWR
port 2 nsew power bidirectional abutment
rlabel viali s 356 423 390 457 6 LOWLVPWR
port 2 nsew power bidirectional abutment
rlabel viali s 284 423 318 457 6 LOWLVPWR
port 2 nsew power bidirectional abutment
rlabel locali s 412 327 478 413 6 LOWLVPWR
port 2 nsew power bidirectional abutment
rlabel locali s 276 413 478 467 6 LOWLVPWR
port 2 nsew power bidirectional abutment
rlabel locali s 412 467 478 532 6 LOWLVPWR
port 2 nsew power bidirectional abutment
rlabel locali s 412 532 562 750 6 LOWLVPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 1040 1472 1136 6 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 1383 893 1469 1050 6 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 3 893 89 1050 6 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1472 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 3 38 89 195 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1409 1071 1443 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1317 1071 1351 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1225 1071 1259 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1133 1071 1167 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1041 1071 1075 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 949 1071 983 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 857 1071 891 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 765 1071 799 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 673 1071 707 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 581 1071 615 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 489 1071 523 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 397 1071 431 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 305 1071 339 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 213 1071 247 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 121 1071 155 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 29 1071 63 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1397 926 1455 1071 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 889 903 991 1071 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 715 903 753 1071 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 529 903 581 1071 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 17 926 75 1071 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 1071 1472 1105 6 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1409 -17 1443 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1317 -17 1351 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1225 -17 1259 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1133 -17 1167 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1041 -17 1075 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 949 -17 983 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 857 -17 891 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 765 -17 799 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 673 -17 707 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 581 -17 615 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 489 -17 523 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 397 -17 431 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 305 -17 339 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 213 -17 247 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 121 -17 155 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 29 -17 63 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 1472 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1351 17 1401 185 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1165 17 1231 169 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 967 17 1033 180 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 795 17 861 112 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 623 17 689 180 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 404 17 470 179 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 17 17 75 162 6 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 1386 691 1444 700 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 16 691 74 700 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 14 700 1458 728 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 1386 728 1444 737 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 16 728 74 737 6 VPB
port 4 nsew power bidirectional
rlabel nwell s 850 261 1481 827 6 VPB
port 4 nsew power bidirectional
rlabel nwell s -38 261 130 827 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 1472 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1409 527 1443 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1317 527 1351 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1225 527 1259 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1133 527 1167 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 1041 527 1075 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1351 322 1387 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1181 322 1215 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 978 325 1024 527 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 978 527 1472 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 978 561 1024 748 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 305 527 339 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 213 527 247 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 121 527 155 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel viali s 29 527 63 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 0 527 378 561 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1267 51 1311 217 6 X
port 6 nsew signal output
rlabel locali s 1067 51 1127 196 6 X
port 6 nsew signal output
rlabel locali s 1072 196 1127 217 6 X
port 6 nsew signal output
rlabel locali s 1072 217 1311 282 6 X
port 6 nsew signal output
rlabel locali s 1256 282 1311 474 6 X
port 6 nsew signal output
rlabel locali s 1072 282 1127 474 6 X
port 6 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE WELLTAP
string FIXED_BBOX 0 0 1472 1088
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1635856
string GDS_START 1621350
<< end >>
