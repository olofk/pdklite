magic
tech sky130A
magscale 1 2
timestamp 1640697850
<< nwell >>
rect 2166 493 2524 1225
<< pwell >>
rect 867 -1510 1119 -1232
<< mvnmos >>
rect 893 -1431 1093 -1311
<< mvpmos >>
rect 2285 559 2405 1159
<< mvndiff >>
rect 893 -1266 1093 -1258
rect 893 -1300 905 -1266
rect 939 -1300 973 -1266
rect 1007 -1300 1041 -1266
rect 1075 -1300 1093 -1266
rect 893 -1311 1093 -1300
rect 893 -1442 1093 -1431
rect 893 -1476 905 -1442
rect 939 -1476 973 -1442
rect 1007 -1476 1041 -1442
rect 1075 -1476 1093 -1442
rect 893 -1484 1093 -1476
<< mvpdiff >>
rect 2232 1147 2285 1159
rect 2232 1113 2240 1147
rect 2274 1113 2285 1147
rect 2232 1079 2285 1113
rect 2232 1045 2240 1079
rect 2274 1045 2285 1079
rect 2232 1011 2285 1045
rect 2232 977 2240 1011
rect 2274 977 2285 1011
rect 2232 943 2285 977
rect 2232 909 2240 943
rect 2274 909 2285 943
rect 2232 875 2285 909
rect 2232 841 2240 875
rect 2274 841 2285 875
rect 2232 807 2285 841
rect 2232 773 2240 807
rect 2274 773 2285 807
rect 2232 739 2285 773
rect 2232 705 2240 739
rect 2274 705 2285 739
rect 2232 671 2285 705
rect 2232 637 2240 671
rect 2274 637 2285 671
rect 2232 559 2285 637
rect 2405 1147 2458 1159
rect 2405 1113 2416 1147
rect 2450 1113 2458 1147
rect 2405 1079 2458 1113
rect 2405 1045 2416 1079
rect 2450 1045 2458 1079
rect 2405 1011 2458 1045
rect 2405 977 2416 1011
rect 2450 977 2458 1011
rect 2405 943 2458 977
rect 2405 909 2416 943
rect 2450 909 2458 943
rect 2405 875 2458 909
rect 2405 841 2416 875
rect 2450 841 2458 875
rect 2405 807 2458 841
rect 2405 773 2416 807
rect 2450 773 2458 807
rect 2405 739 2458 773
rect 2405 705 2416 739
rect 2450 705 2458 739
rect 2405 671 2458 705
rect 2405 637 2416 671
rect 2450 637 2458 671
rect 2405 559 2458 637
<< mvndiffc >>
rect 905 -1300 939 -1266
rect 973 -1300 1007 -1266
rect 1041 -1300 1075 -1266
rect 905 -1476 939 -1442
rect 973 -1476 1007 -1442
rect 1041 -1476 1075 -1442
<< mvpdiffc >>
rect 2240 1113 2274 1147
rect 2240 1045 2274 1079
rect 2240 977 2274 1011
rect 2240 909 2274 943
rect 2240 841 2274 875
rect 2240 773 2274 807
rect 2240 705 2274 739
rect 2240 637 2274 671
rect 2416 1113 2450 1147
rect 2416 1045 2450 1079
rect 2416 977 2450 1011
rect 2416 909 2450 943
rect 2416 841 2450 875
rect 2416 773 2450 807
rect 2416 705 2450 739
rect 2416 637 2450 671
<< poly >>
rect 2285 1159 2405 1185
rect 2285 503 2405 559
rect 2285 469 2334 503
rect 2368 469 2405 503
rect 2285 435 2405 469
rect 2285 401 2334 435
rect 2368 401 2405 435
rect 2285 391 2405 401
rect 2318 385 2384 391
rect 867 -1431 893 -1311
rect 1093 -1362 1263 -1311
rect 1093 -1396 1141 -1362
rect 1175 -1396 1209 -1362
rect 1243 -1396 1263 -1362
rect 1093 -1431 1263 -1396
<< polycont >>
rect 2334 469 2368 503
rect 2334 401 2368 435
rect 1141 -1396 1175 -1362
rect 1209 -1396 1243 -1362
<< locali >>
rect 2241 1163 2275 1183
rect 2240 1147 2275 1163
rect 2274 1145 2275 1147
rect 2240 1111 2241 1113
rect 2240 1079 2275 1111
rect 2274 1073 2275 1079
rect 2240 1039 2241 1045
rect 2401 1147 2453 1174
rect 2401 1113 2416 1147
rect 2450 1113 2453 1147
rect 2401 1079 2453 1113
rect 2401 1045 2416 1079
rect 2450 1045 2453 1079
rect 2240 1011 2274 1039
rect 2240 943 2274 977
rect 2240 875 2274 909
rect 2240 807 2274 841
rect 2240 739 2274 773
rect 2240 671 2274 705
rect 2240 621 2274 637
rect 2401 1011 2453 1045
rect 2401 977 2416 1011
rect 2450 977 2453 1011
rect 2401 953 2453 977
rect 2401 919 2411 953
rect 2445 943 2453 953
rect 2401 909 2416 919
rect 2450 909 2453 943
rect 2401 877 2453 909
rect 2401 843 2411 877
rect 2445 875 2453 877
rect 2401 841 2416 843
rect 2450 841 2453 875
rect 2401 807 2453 841
rect 2401 801 2416 807
rect 2401 767 2411 801
rect 2450 773 2453 807
rect 2445 767 2453 773
rect 2401 739 2453 767
rect 2401 725 2416 739
rect 2401 691 2411 725
rect 2450 705 2453 739
rect 2445 691 2453 705
rect 2401 671 2453 691
rect 2401 650 2416 671
rect 2401 616 2411 650
rect 2450 637 2453 671
rect 2445 616 2453 637
rect 2401 604 2453 616
rect 2201 434 2235 472
rect 2334 503 2368 519
rect 2334 435 2368 469
rect 2334 385 2368 401
rect 1007 -1110 1045 -1076
rect 889 -1300 905 -1266
rect 939 -1300 973 -1266
rect 1007 -1300 1041 -1266
rect 1079 -1300 1091 -1266
rect 1125 -1396 1141 -1362
rect 1178 -1396 1209 -1362
rect 1250 -1396 1259 -1362
rect 889 -1476 905 -1442
rect 939 -1476 973 -1442
rect 1007 -1476 1041 -1442
rect 1079 -1476 1091 -1442
<< viali >>
rect 2241 1183 2275 1217
rect 2241 1113 2274 1145
rect 2274 1113 2275 1145
rect 2241 1111 2275 1113
rect 2241 1045 2274 1073
rect 2274 1045 2275 1073
rect 2241 1039 2275 1045
rect 2411 943 2445 953
rect 2411 919 2416 943
rect 2416 919 2445 943
rect 2411 875 2445 877
rect 2411 843 2416 875
rect 2416 843 2445 875
rect 2411 773 2416 801
rect 2416 773 2445 801
rect 2411 767 2445 773
rect 2411 705 2416 725
rect 2416 705 2445 725
rect 2411 691 2445 705
rect 2411 637 2416 650
rect 2416 637 2445 650
rect 2411 616 2445 637
rect 2201 472 2235 506
rect 2201 400 2235 434
rect 973 -1110 1007 -1076
rect 1045 -1110 1079 -1076
rect 973 -1300 1007 -1266
rect 1045 -1300 1075 -1266
rect 1075 -1300 1079 -1266
rect 1144 -1396 1175 -1362
rect 1175 -1396 1178 -1362
rect 1216 -1396 1243 -1362
rect 1243 -1396 1250 -1362
rect 973 -1476 1007 -1442
rect 1045 -1476 1075 -1442
rect 1075 -1476 1079 -1442
<< metal1 >>
rect 2197 1217 2624 1229
rect 2197 1183 2241 1217
rect 2275 1183 2624 1217
rect 2197 1145 2624 1183
rect 2197 1111 2241 1145
rect 2275 1111 2624 1145
rect 2197 1073 2624 1111
rect 2197 1039 2241 1073
rect 2275 1039 2624 1073
rect 2197 1026 2624 1039
rect 2405 953 2451 965
rect 2405 919 2411 953
rect 2445 919 2451 953
rect 2405 877 2451 919
rect 2405 843 2411 877
rect 2445 843 2451 877
rect 2405 801 2451 843
rect 2405 767 2411 801
rect 2445 767 2451 801
rect 2405 725 2451 767
rect 2405 691 2411 725
rect 2445 691 2451 725
rect 2405 650 2451 691
rect 2405 616 2411 650
rect 2445 616 2451 650
rect 2192 506 2244 519
rect 2192 472 2201 506
rect 2235 472 2244 506
rect 2192 434 2244 472
rect 2192 400 2201 434
rect 2235 400 2244 434
tri 2110 177 2192 259 se
rect 2192 187 2244 400
rect 2192 177 2234 187
tri 2234 177 2244 187 nw
rect 976 125 982 177
rect 1034 125 1046 177
rect 1098 125 2182 177
tri 2182 125 2234 177 nw
rect 2405 79 2451 616
rect 878 27 884 79
rect 936 27 948 79
rect 1000 27 2451 79
rect 961 -1076 975 -1067
rect 961 -1110 973 -1076
rect 961 -1119 975 -1110
rect 1027 -1119 1039 -1067
rect 1091 -1119 1097 -1067
tri 825 -1257 860 -1222 sw
rect 825 -1266 1097 -1257
rect 825 -1300 973 -1266
rect 1007 -1300 1045 -1266
rect 1079 -1300 1097 -1266
rect 825 -1309 1097 -1300
tri 825 -1344 860 -1309 nw
rect 1132 -1405 1138 -1353
rect 1190 -1405 1202 -1353
rect 1254 -1356 1260 -1353
rect 1254 -1402 1262 -1356
rect 1254 -1405 1260 -1402
rect 878 -1458 884 -1406
rect 936 -1458 948 -1406
rect 1000 -1433 1006 -1406
tri 1006 -1433 1033 -1406 sw
rect 1000 -1442 1097 -1433
rect 878 -1476 973 -1458
rect 1007 -1476 1045 -1442
rect 1079 -1476 1097 -1442
rect 878 -1485 1097 -1476
<< via1 >>
rect 982 125 1034 177
rect 1046 125 1098 177
rect 884 27 936 79
rect 948 27 1000 79
rect 975 -1076 1027 -1067
rect 975 -1110 1007 -1076
rect 1007 -1110 1027 -1076
rect 975 -1119 1027 -1110
rect 1039 -1076 1091 -1067
rect 1039 -1110 1045 -1076
rect 1045 -1110 1079 -1076
rect 1079 -1110 1091 -1076
rect 1039 -1119 1091 -1110
rect 1138 -1362 1190 -1353
rect 1138 -1396 1144 -1362
rect 1144 -1396 1178 -1362
rect 1178 -1396 1190 -1362
rect 1138 -1405 1190 -1396
rect 1202 -1362 1254 -1353
rect 1202 -1396 1216 -1362
rect 1216 -1396 1250 -1362
rect 1250 -1396 1254 -1362
rect 1202 -1405 1254 -1396
rect 884 -1458 936 -1406
rect 948 -1442 1000 -1406
rect 948 -1458 973 -1442
rect 973 -1458 1000 -1442
<< metal2 >>
rect 976 125 982 177
rect 1034 125 1046 177
rect 1098 125 1104 177
rect 878 27 884 79
rect 936 27 948 79
rect 1000 27 1006 79
rect 878 -1405 930 27
tri 930 -14 971 27 nw
tri 1018 -1067 1052 -1033 se
rect 1052 -1067 1104 125
rect 969 -1119 975 -1067
rect 1027 -1119 1039 -1067
rect 1091 -1119 1104 -1067
tri 1018 -1153 1052 -1119 ne
rect 1052 -1353 1104 -1119
tri 1104 -1353 1141 -1316 sw
tri 930 -1405 975 -1360 sw
rect 1052 -1405 1138 -1353
rect 1190 -1405 1202 -1353
rect 1254 -1405 1260 -1353
rect 878 -1406 975 -1405
tri 975 -1406 976 -1405 sw
rect 878 -1458 884 -1406
rect 936 -1458 948 -1406
rect 1000 -1458 1006 -1406
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1640697850
transform 0 -1 2275 -1 0 1217
box 0 0 1 1
use sky130_fd_pr__model__nfet_highvoltage__example_5595914180899  sky130_fd_pr__model__nfet_highvoltage__example_5595914180899_0
timestamp 1640697850
transform 0 1 893 1 0 -1431
box -28 0 148 97
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808101  sky130_fd_pr__model__pfet_highvoltage__example_55959141808101_0
timestamp 1640697850
transform 1 0 2285 0 -1 1159
box -28 0 148 267
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 37331040
string GDS_START 37326146
<< end >>
