magic
tech sky130A
magscale 1 2
timestamp 1640697864
<< metal3 >>
rect 10078 2988 14858 3676
<< obsm3 >>
rect 99 2988 4879 3676
<< metal4 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 19000
rect 14746 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 11647 254 12537
rect 14746 11647 15000 12537
rect 0 11281 15000 11347
rect 0 10625 15000 11221
rect 0 10329 254 10565
rect 14746 10329 15000 10565
rect 0 9673 15000 10269
rect 0 9547 15000 9613
rect 0 8317 254 9247
rect 14746 8317 15000 9247
rect 0 7347 254 8037
rect 14746 7347 15000 8037
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 5167 254 6097
rect 14746 5167 15000 6097
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 2987 4874 3677
rect 10083 2987 15000 3677
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< obsm4 >>
rect 334 35077 14666 40000
rect 254 19080 14746 35077
rect 334 13927 14666 19080
rect 254 13787 14746 13927
rect 334 12737 14666 13787
rect 254 12617 14746 12737
rect 334 11567 14666 12617
rect 254 11427 14746 11567
rect 334 10349 14666 10545
rect 254 9327 14746 9467
rect 334 8237 14666 9327
rect 254 8117 14746 8237
rect 334 7267 14666 8117
rect 254 7147 14746 7267
rect 334 6297 14666 7147
rect 254 6177 14746 6297
rect 334 5087 14666 6177
rect 254 4967 14746 5087
rect 334 3877 14666 4967
rect 254 3757 14746 3877
rect 4954 2907 10003 3757
rect 254 2787 14746 2907
rect 334 1697 14666 2787
rect 254 1577 14746 1697
rect 334 407 14666 1577
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 18997
rect 0 12837 254 13687
rect 0 11667 254 12517
rect 0 9547 254 11347
rect 0 8337 254 9227
rect 0 7368 254 8017
rect 14746 14007 15000 18997
rect 14746 12837 15000 13687
rect 14746 11667 15000 12517
rect 14746 9547 15000 11347
rect 14746 8337 15000 9227
rect 14746 7368 15000 8017
rect 0 6397 254 7047
rect 0 5187 254 6077
rect 0 3977 254 4867
rect 14746 6397 15000 7047
rect 14746 5187 15000 6077
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 0 427 254 1477
rect 14746 1797 15000 2687
rect 14746 427 15000 1477
<< obsm5 >>
rect 574 34837 14426 40000
rect 0 19317 15000 34837
rect 574 7368 14426 19317
rect 0 7367 15000 7368
rect 574 3657 14426 7367
rect 513 3007 14487 3657
rect 574 427 14426 3007
<< labels >>
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 1 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 1 nsew power bidirectional
rlabel metal4 s 14746 1777 15000 2707 6 VCCD
port 1 nsew power bidirectional
rlabel metal4 s 0 1777 254 2707 6 VCCD
port 1 nsew power bidirectional
rlabel metal4 s 14746 1777 15000 2707 6 VCCD
port 1 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 1 nsew power bidirectional
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 1 nsew power bidirectional
rlabel metal4 s 14746 1777 15000 2707 6 VCCD
port 1 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 1 nsew power bidirectional
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 1 nsew power bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 2 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 2 nsew power bidirectional
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 2 nsew power bidirectional
rlabel metal4 s 0 6377 254 7067 6 VSWITCH
port 2 nsew power bidirectional
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 2 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 2 nsew power bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 2 nsew power bidirectional
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 2 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 2 nsew power bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 2 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal4 s 0 407 254 1497 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 9547 15000 9613 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 11281 15000 11347 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 7347 254 8037 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14746 7347 15000 8037 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14746 9547 15000 9613 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14746 11281 15000 11347 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 9547 254 9613 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 11281 254 11347 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14746 7347 15000 8037 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14746 9547 15000 9613 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14746 11281 15000 11347 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 9547 254 9613 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 11281 254 11347 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14746 7347 15000 8037 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14746 9547 15000 9613 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14746 11281 15000 11347 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 5 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 5 nsew power bidirectional
rlabel metal4 s 0 2987 193 3677 6 VDDA
port 5 nsew power bidirectional
rlabel metal4 s 14807 2987 15000 3677 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10078 2988 14858 3676 6 VDDA
port 5 nsew power bidirectional
rlabel metal4 s 0 2987 4874 3677 6 VDDA
port 5 nsew power bidirectional
rlabel metal4 s 10083 2987 15000 3677 6 VDDA
port 5 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 5 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3620 14840 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3532 14840 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3444 14840 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3356 14840 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3268 14840 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3180 14840 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3092 14840 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3004 14840 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3620 14759 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3532 14759 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3444 14759 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3356 14759 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3268 14759 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3180 14759 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3092 14759 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3004 14759 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3620 14678 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3532 14678 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3444 14678 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3356 14678 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3268 14678 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3180 14678 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3092 14678 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3004 14678 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3620 14597 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3532 14597 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3444 14597 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3356 14597 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3268 14597 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3180 14597 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3092 14597 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3004 14597 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3620 14516 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3532 14516 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3444 14516 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3356 14516 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3268 14516 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3180 14516 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3092 14516 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3004 14516 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3620 14435 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3532 14435 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3444 14435 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3356 14435 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3268 14435 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3180 14435 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3092 14435 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3004 14435 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3620 14354 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3532 14354 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3444 14354 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3356 14354 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3268 14354 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3180 14354 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3092 14354 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3004 14354 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3620 14273 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3532 14273 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3444 14273 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3356 14273 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3268 14273 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3180 14273 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3092 14273 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3004 14273 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3620 14192 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3532 14192 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3444 14192 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3356 14192 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3268 14192 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3180 14192 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3092 14192 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3004 14192 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3620 14111 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3532 14111 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3444 14111 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3356 14111 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3268 14111 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3180 14111 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3092 14111 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3004 14111 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3620 14030 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3532 14030 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3444 14030 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3356 14030 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3268 14030 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3180 14030 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3092 14030 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3004 14030 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3620 13949 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3532 13949 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3444 13949 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3356 13949 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3268 13949 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3180 13949 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3092 13949 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3004 13949 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3620 13868 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3532 13868 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3444 13868 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3356 13868 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3268 13868 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3180 13868 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3092 13868 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3004 13868 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3620 13787 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3532 13787 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3444 13787 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3356 13787 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3268 13787 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3180 13787 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3092 13787 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3004 13787 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3620 13706 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3532 13706 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3444 13706 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3356 13706 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3268 13706 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3180 13706 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3092 13706 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3004 13706 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3620 13625 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3532 13625 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3444 13625 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3356 13625 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3268 13625 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3180 13625 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3092 13625 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3004 13625 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3620 13544 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3532 13544 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3444 13544 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3356 13544 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3268 13544 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3180 13544 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3092 13544 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3004 13544 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3620 13463 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3532 13463 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3444 13463 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3356 13463 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3268 13463 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3180 13463 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3092 13463 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3004 13463 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3620 13382 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3532 13382 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3444 13382 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3356 13382 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3268 13382 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3180 13382 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3092 13382 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3004 13382 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3620 13301 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3532 13301 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3444 13301 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3356 13301 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3268 13301 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3180 13301 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3092 13301 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3004 13301 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3620 13220 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3532 13220 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3444 13220 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3356 13220 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3268 13220 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3180 13220 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3092 13220 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3004 13220 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3620 13139 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3532 13139 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3444 13139 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3356 13139 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3268 13139 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3180 13139 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3092 13139 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3004 13139 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3620 13058 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3532 13058 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3444 13058 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3356 13058 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3268 13058 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3180 13058 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3092 13058 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3004 13058 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3620 12977 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3532 12977 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3444 12977 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3356 12977 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3268 12977 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3180 12977 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3092 12977 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3004 12977 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3620 12896 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3532 12896 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3444 12896 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3356 12896 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3268 12896 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3180 12896 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3092 12896 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3004 12896 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3620 12815 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3532 12815 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3444 12815 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3356 12815 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3268 12815 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3180 12815 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3092 12815 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3004 12815 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3620 12734 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3532 12734 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3444 12734 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3356 12734 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3268 12734 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3180 12734 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3092 12734 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3004 12734 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3620 12653 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3532 12653 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3444 12653 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3356 12653 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3268 12653 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3180 12653 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3092 12653 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3004 12653 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3620 12572 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3532 12572 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3444 12572 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3356 12572 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3268 12572 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3180 12572 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3092 12572 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3004 12572 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3620 12491 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3532 12491 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3444 12491 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3356 12491 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3268 12491 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3180 12491 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3092 12491 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3004 12491 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3620 12410 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3532 12410 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3444 12410 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3356 12410 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3268 12410 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3180 12410 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3092 12410 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3004 12410 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3620 12329 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3532 12329 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3444 12329 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3356 12329 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3268 12329 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3180 12329 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3092 12329 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3004 12329 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3620 12248 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3532 12248 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3444 12248 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3356 12248 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3268 12248 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3180 12248 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3092 12248 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3004 12248 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3620 12167 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3532 12167 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3444 12167 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3356 12167 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3268 12167 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3180 12167 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3092 12167 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3004 12167 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3620 12086 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3532 12086 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3444 12086 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3356 12086 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3268 12086 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3180 12086 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3092 12086 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3004 12086 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3620 12005 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3532 12005 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3444 12005 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3356 12005 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3268 12005 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3180 12005 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3092 12005 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3004 12005 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3620 11924 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3532 11924 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3444 11924 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3356 11924 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3268 11924 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3180 11924 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3092 11924 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3004 11924 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3620 11843 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3532 11843 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3444 11843 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3356 11843 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3268 11843 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3180 11843 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3092 11843 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3004 11843 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3620 11762 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3532 11762 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3444 11762 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3356 11762 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3268 11762 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3180 11762 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3092 11762 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3004 11762 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3620 11681 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3532 11681 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3444 11681 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3356 11681 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3268 11681 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3180 11681 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3092 11681 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3004 11681 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3620 11600 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3532 11600 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3444 11600 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3356 11600 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3268 11600 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3180 11600 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3092 11600 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3004 11600 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3620 11519 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3532 11519 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3444 11519 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3356 11519 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3268 11519 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3180 11519 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3092 11519 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3004 11519 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3620 11438 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3532 11438 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3444 11438 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3356 11438 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3268 11438 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3180 11438 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3092 11438 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3004 11438 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3620 11357 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3532 11357 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3444 11357 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3356 11357 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3268 11357 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3180 11357 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3092 11357 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3004 11357 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3620 11276 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3532 11276 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3444 11276 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3356 11276 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3268 11276 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3180 11276 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3092 11276 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3004 11276 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3620 11195 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3532 11195 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3444 11195 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3356 11195 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3268 11195 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3180 11195 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3092 11195 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3004 11195 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3620 11114 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3532 11114 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3444 11114 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3356 11114 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3268 11114 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3180 11114 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3092 11114 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3004 11114 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3620 11033 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3532 11033 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3444 11033 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3356 11033 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3268 11033 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3180 11033 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3092 11033 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3004 11033 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3620 10952 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3532 10952 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3444 10952 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3356 10952 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3268 10952 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3180 10952 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3092 10952 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3004 10952 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3620 10871 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3532 10871 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3444 10871 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3356 10871 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3268 10871 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3180 10871 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3092 10871 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3004 10871 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3620 10790 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3532 10790 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3444 10790 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3356 10790 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3268 10790 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3180 10790 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3092 10790 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3004 10790 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3620 10709 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3532 10709 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3444 10709 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3356 10709 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3268 10709 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3180 10709 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3092 10709 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3004 10709 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3620 10628 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3532 10628 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3444 10628 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3356 10628 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3268 10628 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3180 10628 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3092 10628 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3004 10628 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3620 10546 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3532 10546 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3444 10546 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3356 10546 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3268 10546 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3180 10546 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3092 10546 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3004 10546 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3620 10464 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3532 10464 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3444 10464 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3356 10464 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3268 10464 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3180 10464 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3092 10464 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3004 10464 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3620 10382 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3532 10382 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3444 10382 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3356 10382 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3268 10382 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3180 10382 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3092 10382 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3004 10382 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3620 10300 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3532 10300 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3444 10300 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3356 10300 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3268 10300 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3180 10300 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3092 10300 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3004 10300 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3620 10218 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3532 10218 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3444 10218 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3356 10218 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3268 10218 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3180 10218 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3092 10218 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3004 10218 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3620 10136 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3532 10136 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3444 10136 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3356 10136 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3268 10136 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3180 10136 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3092 10136 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3004 10136 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4809 3608 4873 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4809 3520 4873 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4809 3432 4873 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4809 3344 4873 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4809 3256 4873 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4809 3168 4873 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4809 3080 4873 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4809 2992 4873 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4728 3608 4792 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4728 3520 4792 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4728 3432 4792 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4728 3344 4792 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4728 3256 4792 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4728 3168 4792 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4728 3080 4792 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4728 2992 4792 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4647 3608 4711 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4647 3520 4711 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4647 3432 4711 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4647 3344 4711 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4647 3256 4711 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4647 3168 4711 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4647 3080 4711 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4647 2992 4711 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4566 3608 4630 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4566 3520 4630 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4566 3432 4630 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4566 3344 4630 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4566 3256 4630 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4566 3168 4630 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4566 3080 4630 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4566 2992 4630 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4485 3608 4549 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4485 3520 4549 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4485 3432 4549 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4485 3344 4549 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4485 3256 4549 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4485 3168 4549 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4485 3080 4549 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4485 2992 4549 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4404 3608 4468 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4404 3520 4468 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4404 3432 4468 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4404 3344 4468 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4404 3256 4468 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4404 3168 4468 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4404 3080 4468 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4404 2992 4468 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4323 3608 4387 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4323 3520 4387 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4323 3432 4387 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4323 3344 4387 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4323 3256 4387 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4323 3168 4387 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4323 3080 4387 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4323 2992 4387 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4242 3608 4306 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4242 3520 4306 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4242 3432 4306 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4242 3344 4306 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4242 3256 4306 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4242 3168 4306 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4242 3080 4306 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4242 2992 4306 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4161 3608 4225 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4161 3520 4225 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4161 3432 4225 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4161 3344 4225 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4161 3256 4225 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4161 3168 4225 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4161 3080 4225 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4161 2992 4225 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4080 3608 4144 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4080 3520 4144 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4080 3432 4144 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4080 3344 4144 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4080 3256 4144 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4080 3168 4144 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4080 3080 4144 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4080 2992 4144 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3999 3608 4063 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3999 3520 4063 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3999 3432 4063 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3999 3344 4063 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3999 3256 4063 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3999 3168 4063 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3999 3080 4063 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3999 2992 4063 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3918 3608 3982 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3918 3520 3982 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3918 3432 3982 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3918 3344 3982 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3918 3256 3982 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3918 3168 3982 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3918 3080 3982 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3918 2992 3982 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3837 3608 3901 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3837 3520 3901 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3837 3432 3901 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3837 3344 3901 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3837 3256 3901 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3837 3168 3901 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3837 3080 3901 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3837 2992 3901 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3756 3608 3820 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3756 3520 3820 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3756 3432 3820 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3756 3344 3820 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3756 3256 3820 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3756 3168 3820 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3756 3080 3820 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3756 2992 3820 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3675 3608 3739 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3675 3520 3739 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3675 3432 3739 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3675 3344 3739 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3675 3256 3739 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3675 3168 3739 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3675 3080 3739 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3675 2992 3739 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3594 3608 3658 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3594 3520 3658 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3594 3432 3658 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3594 3344 3658 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3594 3256 3658 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3594 3168 3658 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3594 3080 3658 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3594 2992 3658 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3513 3608 3577 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3513 3520 3577 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3513 3432 3577 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3513 3344 3577 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3513 3256 3577 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3513 3168 3577 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3513 3080 3577 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3513 2992 3577 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3432 3608 3496 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3432 3520 3496 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3432 3432 3496 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3432 3344 3496 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3432 3256 3496 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3432 3168 3496 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3432 3080 3496 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3432 2992 3496 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3351 3608 3415 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3351 3520 3415 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3351 3432 3415 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3351 3344 3415 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3351 3256 3415 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3351 3168 3415 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3351 3080 3415 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3351 2992 3415 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3270 3608 3334 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3270 3520 3334 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3270 3432 3334 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3270 3344 3334 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3270 3256 3334 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3270 3168 3334 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3270 3080 3334 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3270 2992 3334 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3189 3608 3253 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3189 3520 3253 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3189 3432 3253 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3189 3344 3253 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3189 3256 3253 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3189 3168 3253 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3189 3080 3253 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3189 2992 3253 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3108 3608 3172 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3108 3520 3172 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3108 3432 3172 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3108 3344 3172 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3108 3256 3172 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3108 3168 3172 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3108 3080 3172 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3108 2992 3172 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3027 3608 3091 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3027 3520 3091 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3027 3432 3091 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3027 3344 3091 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3027 3256 3091 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3027 3168 3091 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3027 3080 3091 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3027 2992 3091 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2946 3608 3010 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2946 3520 3010 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2946 3432 3010 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2946 3344 3010 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2946 3256 3010 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2946 3168 3010 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2946 3080 3010 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2946 2992 3010 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2865 3608 2929 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2865 3520 2929 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2865 3432 2929 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2865 3344 2929 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2865 3256 2929 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2865 3168 2929 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2865 3080 2929 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2865 2992 2929 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2784 3608 2848 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2784 3520 2848 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2784 3432 2848 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2784 3344 2848 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2784 3256 2848 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2784 3168 2848 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2784 3080 2848 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2784 2992 2848 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2703 3608 2767 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2703 3520 2767 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2703 3432 2767 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2703 3344 2767 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2703 3256 2767 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2703 3168 2767 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2703 3080 2767 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2703 2992 2767 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2622 3608 2686 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2622 3520 2686 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2622 3432 2686 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2622 3344 2686 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2622 3256 2686 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2622 3168 2686 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2622 3080 2686 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2622 2992 2686 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2541 3608 2605 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2541 3520 2605 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2541 3432 2605 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2541 3344 2605 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2541 3256 2605 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2541 3168 2605 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2541 3080 2605 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2541 2992 2605 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2460 3608 2524 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2460 3520 2524 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2460 3432 2524 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2460 3344 2524 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2460 3256 2524 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2460 3168 2524 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2460 3080 2524 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2460 2992 2524 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2379 3608 2443 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2379 3520 2443 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2379 3432 2443 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2379 3344 2443 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2379 3256 2443 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2379 3168 2443 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2379 3080 2443 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2379 2992 2443 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2298 3608 2362 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2298 3520 2362 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2298 3432 2362 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2298 3344 2362 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2298 3256 2362 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2298 3168 2362 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2298 3080 2362 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2298 2992 2362 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2217 3608 2281 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2217 3520 2281 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2217 3432 2281 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2217 3344 2281 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2217 3256 2281 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2217 3168 2281 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2217 3080 2281 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2217 2992 2281 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2136 3608 2200 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2136 3520 2200 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2136 3432 2200 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2136 3344 2200 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2136 3256 2200 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2136 3168 2200 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2136 3080 2200 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2136 2992 2200 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2055 3608 2119 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2055 3520 2119 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2055 3432 2119 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2055 3344 2119 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2055 3256 2119 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2055 3168 2119 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2055 3080 2119 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2055 2992 2119 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1974 3608 2038 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1974 3520 2038 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1974 3432 2038 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1974 3344 2038 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1974 3256 2038 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1974 3168 2038 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1974 3080 2038 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1974 2992 2038 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1893 3608 1957 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1893 3520 1957 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1893 3432 1957 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1893 3344 1957 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1893 3256 1957 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1893 3168 1957 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1893 3080 1957 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1893 2992 1957 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1812 3608 1876 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1812 3520 1876 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1812 3432 1876 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1812 3344 1876 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1812 3256 1876 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1812 3168 1876 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1812 3080 1876 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1812 2992 1876 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1731 3608 1795 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1731 3520 1795 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1731 3432 1795 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1731 3344 1795 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1731 3256 1795 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1731 3168 1795 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1731 3080 1795 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1731 2992 1795 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1650 3608 1714 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1650 3520 1714 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1650 3432 1714 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1650 3344 1714 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1650 3256 1714 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1650 3168 1714 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1650 3080 1714 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1650 2992 1714 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1569 3608 1633 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1569 3520 1633 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1569 3432 1633 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1569 3344 1633 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1569 3256 1633 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1569 3168 1633 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1569 3080 1633 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1569 2992 1633 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1488 3608 1552 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1488 3520 1552 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1488 3432 1552 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1488 3344 1552 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1488 3256 1552 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1488 3168 1552 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1488 3080 1552 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1488 2992 1552 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1407 3608 1471 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1407 3520 1471 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1407 3432 1471 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1407 3344 1471 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1407 3256 1471 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1407 3168 1471 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1407 3080 1471 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1407 2992 1471 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1326 3608 1390 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1326 3520 1390 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1326 3432 1390 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1326 3344 1390 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1326 3256 1390 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1326 3168 1390 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1326 3080 1390 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1326 2992 1390 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1245 3608 1309 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1245 3520 1309 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1245 3432 1309 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1245 3344 1309 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1245 3256 1309 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1245 3168 1309 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1245 3080 1309 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1245 2992 1309 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1164 3608 1228 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1164 3520 1228 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1164 3432 1228 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1164 3344 1228 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1164 3256 1228 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1164 3168 1228 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1164 3080 1228 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1164 2992 1228 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1083 3608 1147 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1083 3520 1147 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1083 3432 1147 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1083 3344 1147 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1083 3256 1147 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1083 3168 1147 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1083 3080 1147 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1083 2992 1147 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1002 3608 1066 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1002 3520 1066 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1002 3432 1066 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1002 3344 1066 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1002 3256 1066 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1002 3168 1066 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1002 3080 1066 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1002 2992 1066 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 921 3608 985 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 921 3520 985 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 921 3432 985 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 921 3344 985 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 921 3256 985 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 921 3168 985 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 921 3080 985 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 921 2992 985 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 840 3608 904 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 840 3520 904 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 840 3432 904 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 840 3344 904 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 840 3256 904 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 840 3168 904 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 840 3080 904 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 840 2992 904 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 759 3608 823 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 759 3520 823 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 759 3432 823 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 759 3344 823 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 759 3256 823 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 759 3168 823 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 759 3080 823 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 759 2992 823 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 678 3608 742 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 678 3520 742 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 678 3432 742 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 678 3344 742 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 678 3256 742 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 678 3168 742 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 678 3080 742 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 678 2992 742 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 597 3608 661 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 597 3520 661 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 597 3432 661 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 597 3344 661 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 597 3256 661 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 597 3168 661 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 597 3080 661 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 597 2992 661 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 515 3608 579 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 515 3520 579 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 515 3432 579 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 515 3344 579 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 515 3256 579 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 515 3168 579 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 515 3080 579 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 515 2992 579 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 433 3608 497 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 433 3520 497 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 433 3432 497 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 433 3344 497 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 433 3256 497 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 433 3168 497 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 433 3080 497 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 433 2992 497 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 351 3608 415 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 351 3520 415 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 351 3432 415 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 351 3344 415 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 351 3256 415 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 351 3168 415 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 351 3080 415 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 351 2992 415 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 269 3608 333 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 269 3520 333 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 269 3432 333 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 269 3344 333 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 269 3256 333 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 269 3168 333 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 269 3080 333 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 269 2992 333 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 187 3608 251 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 187 3520 251 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 187 3432 251 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 187 3344 251 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 187 3256 251 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 187 3168 251 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 187 3080 251 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 187 2992 251 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 105 3608 169 3672 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 105 3520 169 3584 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 105 3432 169 3496 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 105 3344 169 3408 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 105 3256 169 3320 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 105 3168 169 3232 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 105 3080 169 3144 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 105 2992 169 3056 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10078 2988 14858 3676 6 VDDA
port 5 nsew power bidirectional
rlabel metal4 s 0 2987 4874 3677 6 VDDA
port 5 nsew power bidirectional
rlabel metal4 s 10083 2987 15000 3677 6 VDDA
port 5 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 5 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3620 14840 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3532 14840 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3444 14840 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3356 14840 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3268 14840 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3180 14840 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3092 14840 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14800 3004 14840 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3620 14759 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3532 14759 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3444 14759 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3356 14759 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3268 14759 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3180 14759 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3092 14759 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14719 3004 14759 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3620 14678 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3532 14678 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3444 14678 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3356 14678 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3268 14678 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3180 14678 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3092 14678 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14638 3004 14678 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3620 14597 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3532 14597 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3444 14597 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3356 14597 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3268 14597 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3180 14597 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3092 14597 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14557 3004 14597 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3620 14516 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3532 14516 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3444 14516 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3356 14516 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3268 14516 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3180 14516 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3092 14516 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14476 3004 14516 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3620 14435 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3532 14435 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3444 14435 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3356 14435 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3268 14435 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3180 14435 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3092 14435 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14395 3004 14435 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3620 14354 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3532 14354 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3444 14354 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3356 14354 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3268 14354 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3180 14354 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3092 14354 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14314 3004 14354 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3620 14273 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3532 14273 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3444 14273 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3356 14273 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3268 14273 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3180 14273 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3092 14273 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14233 3004 14273 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3620 14192 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3532 14192 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3444 14192 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3356 14192 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3268 14192 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3180 14192 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3092 14192 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14152 3004 14192 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3620 14111 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3532 14111 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3444 14111 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3356 14111 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3268 14111 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3180 14111 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3092 14111 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 14071 3004 14111 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3620 14030 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3532 14030 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3444 14030 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3356 14030 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3268 14030 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3180 14030 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3092 14030 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13990 3004 14030 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3620 13949 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3532 13949 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3444 13949 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3356 13949 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3268 13949 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3180 13949 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3092 13949 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13909 3004 13949 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3620 13868 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3532 13868 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3444 13868 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3356 13868 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3268 13868 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3180 13868 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3092 13868 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13828 3004 13868 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3620 13787 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3532 13787 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3444 13787 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3356 13787 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3268 13787 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3180 13787 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3092 13787 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13747 3004 13787 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3620 13706 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3532 13706 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3444 13706 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3356 13706 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3268 13706 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3180 13706 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3092 13706 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13666 3004 13706 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3620 13625 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3532 13625 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3444 13625 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3356 13625 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3268 13625 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3180 13625 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3092 13625 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13585 3004 13625 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3620 13544 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3532 13544 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3444 13544 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3356 13544 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3268 13544 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3180 13544 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3092 13544 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13504 3004 13544 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3620 13463 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3532 13463 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3444 13463 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3356 13463 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3268 13463 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3180 13463 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3092 13463 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13423 3004 13463 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3620 13382 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3532 13382 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3444 13382 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3356 13382 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3268 13382 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3180 13382 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3092 13382 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13342 3004 13382 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3620 13301 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3532 13301 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3444 13301 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3356 13301 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3268 13301 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3180 13301 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3092 13301 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13261 3004 13301 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3620 13220 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3532 13220 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3444 13220 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3356 13220 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3268 13220 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3180 13220 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3092 13220 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13180 3004 13220 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3620 13139 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3532 13139 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3444 13139 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3356 13139 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3268 13139 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3180 13139 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3092 13139 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13099 3004 13139 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3620 13058 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3532 13058 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3444 13058 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3356 13058 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3268 13058 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3180 13058 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3092 13058 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 13018 3004 13058 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3620 12977 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3532 12977 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3444 12977 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3356 12977 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3268 12977 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3180 12977 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3092 12977 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12937 3004 12977 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3620 12896 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3532 12896 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3444 12896 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3356 12896 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3268 12896 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3180 12896 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3092 12896 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12856 3004 12896 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3620 12815 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3532 12815 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3444 12815 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3356 12815 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3268 12815 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3180 12815 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3092 12815 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12775 3004 12815 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3620 12734 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3532 12734 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3444 12734 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3356 12734 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3268 12734 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3180 12734 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3092 12734 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12694 3004 12734 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3620 12653 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3532 12653 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3444 12653 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3356 12653 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3268 12653 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3180 12653 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3092 12653 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12613 3004 12653 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3620 12572 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3532 12572 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3444 12572 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3356 12572 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3268 12572 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3180 12572 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3092 12572 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12532 3004 12572 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3620 12491 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3532 12491 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3444 12491 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3356 12491 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3268 12491 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3180 12491 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3092 12491 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12451 3004 12491 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3620 12410 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3532 12410 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3444 12410 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3356 12410 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3268 12410 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3180 12410 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3092 12410 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12370 3004 12410 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3620 12329 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3532 12329 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3444 12329 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3356 12329 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3268 12329 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3180 12329 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3092 12329 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12289 3004 12329 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3620 12248 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3532 12248 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3444 12248 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3356 12248 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3268 12248 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3180 12248 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3092 12248 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12208 3004 12248 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3620 12167 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3532 12167 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3444 12167 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3356 12167 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3268 12167 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3180 12167 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3092 12167 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12127 3004 12167 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3620 12086 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3532 12086 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3444 12086 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3356 12086 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3268 12086 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3180 12086 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3092 12086 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 12046 3004 12086 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3620 12005 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3532 12005 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3444 12005 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3356 12005 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3268 12005 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3180 12005 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3092 12005 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11965 3004 12005 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3620 11924 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3532 11924 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3444 11924 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3356 11924 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3268 11924 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3180 11924 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3092 11924 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11884 3004 11924 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3620 11843 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3532 11843 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3444 11843 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3356 11843 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3268 11843 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3180 11843 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3092 11843 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11803 3004 11843 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3620 11762 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3532 11762 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3444 11762 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3356 11762 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3268 11762 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3180 11762 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3092 11762 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11722 3004 11762 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3620 11681 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3532 11681 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3444 11681 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3356 11681 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3268 11681 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3180 11681 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3092 11681 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11641 3004 11681 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3620 11600 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3532 11600 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3444 11600 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3356 11600 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3268 11600 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3180 11600 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3092 11600 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11560 3004 11600 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3620 11519 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3532 11519 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3444 11519 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3356 11519 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3268 11519 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3180 11519 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3092 11519 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11479 3004 11519 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3620 11438 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3532 11438 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3444 11438 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3356 11438 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3268 11438 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3180 11438 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3092 11438 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11398 3004 11438 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3620 11357 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3532 11357 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3444 11357 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3356 11357 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3268 11357 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3180 11357 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3092 11357 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11317 3004 11357 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3620 11276 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3532 11276 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3444 11276 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3356 11276 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3268 11276 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3180 11276 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3092 11276 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11236 3004 11276 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3620 11195 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3532 11195 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3444 11195 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3356 11195 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3268 11195 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3180 11195 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3092 11195 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11155 3004 11195 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3620 11114 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3532 11114 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3444 11114 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3356 11114 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3268 11114 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3180 11114 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3092 11114 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 11074 3004 11114 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3620 11033 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3532 11033 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3444 11033 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3356 11033 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3268 11033 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3180 11033 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3092 11033 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10993 3004 11033 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3620 10952 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3532 10952 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3444 10952 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3356 10952 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3268 10952 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3180 10952 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3092 10952 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10912 3004 10952 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3620 10871 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3532 10871 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3444 10871 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3356 10871 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3268 10871 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3180 10871 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3092 10871 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10831 3004 10871 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3620 10790 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3532 10790 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3444 10790 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3356 10790 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3268 10790 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3180 10790 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3092 10790 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10750 3004 10790 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3620 10709 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3532 10709 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3444 10709 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3356 10709 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3268 10709 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3180 10709 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3092 10709 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10669 3004 10709 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3620 10628 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3532 10628 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3444 10628 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3356 10628 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3268 10628 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3180 10628 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3092 10628 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10588 3004 10628 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3620 10546 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3532 10546 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3444 10546 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3356 10546 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3268 10546 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3180 10546 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3092 10546 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10506 3004 10546 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3620 10464 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3532 10464 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3444 10464 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3356 10464 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3268 10464 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3180 10464 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3092 10464 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10424 3004 10464 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3620 10382 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3532 10382 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3444 10382 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3356 10382 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3268 10382 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3180 10382 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3092 10382 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10342 3004 10382 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3620 10300 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3532 10300 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3444 10300 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3356 10300 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3268 10300 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3180 10300 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3092 10300 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10260 3004 10300 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3620 10218 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3532 10218 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3444 10218 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3356 10218 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3268 10218 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3180 10218 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3092 10218 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10178 3004 10218 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3620 10136 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3532 10136 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3444 10136 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3356 10136 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3268 10136 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3180 10136 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3092 10136 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 10096 3004 10136 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4821 3620 4861 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4821 3532 4861 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4821 3444 4861 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4821 3356 4861 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4821 3268 4861 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4821 3180 4861 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4821 3092 4861 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4821 3004 4861 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4740 3620 4780 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4740 3532 4780 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4740 3444 4780 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4740 3356 4780 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4740 3268 4780 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4740 3180 4780 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4740 3092 4780 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4740 3004 4780 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4659 3620 4699 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4659 3532 4699 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4659 3444 4699 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4659 3356 4699 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4659 3268 4699 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4659 3180 4699 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4659 3092 4699 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4659 3004 4699 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4578 3620 4618 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4578 3532 4618 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4578 3444 4618 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4578 3356 4618 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4578 3268 4618 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4578 3180 4618 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4578 3092 4618 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4578 3004 4618 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4497 3620 4537 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4497 3532 4537 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4497 3444 4537 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4497 3356 4537 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4497 3268 4537 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4497 3180 4537 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4497 3092 4537 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4497 3004 4537 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4416 3620 4456 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4416 3532 4456 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4416 3444 4456 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4416 3356 4456 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4416 3268 4456 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4416 3180 4456 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4416 3092 4456 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4416 3004 4456 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4335 3620 4375 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4335 3532 4375 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4335 3444 4375 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4335 3356 4375 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4335 3268 4375 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4335 3180 4375 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4335 3092 4375 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4335 3004 4375 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4254 3620 4294 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4254 3532 4294 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4254 3444 4294 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4254 3356 4294 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4254 3268 4294 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4254 3180 4294 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4254 3092 4294 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4254 3004 4294 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4173 3620 4213 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4173 3532 4213 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4173 3444 4213 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4173 3356 4213 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4173 3268 4213 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4173 3180 4213 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4173 3092 4213 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4173 3004 4213 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4092 3620 4132 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4092 3532 4132 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4092 3444 4132 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4092 3356 4132 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4092 3268 4132 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4092 3180 4132 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4092 3092 4132 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4092 3004 4132 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4011 3620 4051 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4011 3532 4051 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4011 3444 4051 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4011 3356 4051 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4011 3268 4051 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4011 3180 4051 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4011 3092 4051 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 4011 3004 4051 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3930 3620 3970 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3930 3532 3970 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3930 3444 3970 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3930 3356 3970 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3930 3268 3970 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3930 3180 3970 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3930 3092 3970 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3930 3004 3970 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3849 3620 3889 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3849 3532 3889 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3849 3444 3889 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3849 3356 3889 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3849 3268 3889 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3849 3180 3889 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3849 3092 3889 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3849 3004 3889 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3768 3620 3808 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3768 3532 3808 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3768 3444 3808 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3768 3356 3808 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3768 3268 3808 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3768 3180 3808 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3768 3092 3808 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3768 3004 3808 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3687 3620 3727 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3687 3532 3727 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3687 3444 3727 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3687 3356 3727 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3687 3268 3727 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3687 3180 3727 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3687 3092 3727 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3687 3004 3727 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3606 3620 3646 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3606 3532 3646 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3606 3444 3646 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3606 3356 3646 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3606 3268 3646 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3606 3180 3646 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3606 3092 3646 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3606 3004 3646 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3525 3620 3565 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3525 3532 3565 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3525 3444 3565 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3525 3356 3565 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3525 3268 3565 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3525 3180 3565 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3525 3092 3565 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3525 3004 3565 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3444 3620 3484 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3444 3532 3484 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3444 3444 3484 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3444 3356 3484 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3444 3268 3484 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3444 3180 3484 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3444 3092 3484 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3444 3004 3484 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3363 3620 3403 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3363 3532 3403 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3363 3444 3403 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3363 3356 3403 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3363 3268 3403 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3363 3180 3403 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3363 3092 3403 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3363 3004 3403 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3282 3620 3322 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3282 3532 3322 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3282 3444 3322 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3282 3356 3322 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3282 3268 3322 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3282 3180 3322 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3282 3092 3322 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3282 3004 3322 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3201 3620 3241 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3201 3532 3241 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3201 3444 3241 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3201 3356 3241 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3201 3268 3241 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3201 3180 3241 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3201 3092 3241 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3201 3004 3241 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3120 3620 3160 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3120 3532 3160 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3120 3444 3160 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3120 3356 3160 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3120 3268 3160 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3120 3180 3160 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3120 3092 3160 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3120 3004 3160 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3039 3620 3079 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3039 3532 3079 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3039 3444 3079 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3039 3356 3079 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3039 3268 3079 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3039 3180 3079 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3039 3092 3079 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 3039 3004 3079 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2958 3620 2998 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2958 3532 2998 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2958 3444 2998 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2958 3356 2998 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2958 3268 2998 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2958 3180 2998 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2958 3092 2998 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2958 3004 2998 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2877 3620 2917 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2877 3532 2917 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2877 3444 2917 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2877 3356 2917 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2877 3268 2917 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2877 3180 2917 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2877 3092 2917 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2877 3004 2917 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2796 3620 2836 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2796 3532 2836 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2796 3444 2836 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2796 3356 2836 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2796 3268 2836 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2796 3180 2836 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2796 3092 2836 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2796 3004 2836 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2715 3620 2755 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2715 3532 2755 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2715 3444 2755 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2715 3356 2755 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2715 3268 2755 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2715 3180 2755 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2715 3092 2755 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2715 3004 2755 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2634 3620 2674 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2634 3532 2674 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2634 3444 2674 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2634 3356 2674 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2634 3268 2674 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2634 3180 2674 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2634 3092 2674 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2634 3004 2674 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2553 3620 2593 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2553 3532 2593 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2553 3444 2593 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2553 3356 2593 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2553 3268 2593 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2553 3180 2593 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2553 3092 2593 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2553 3004 2593 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2472 3620 2512 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2472 3532 2512 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2472 3444 2512 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2472 3356 2512 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2472 3268 2512 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2472 3180 2512 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2472 3092 2512 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2472 3004 2512 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2391 3620 2431 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2391 3532 2431 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2391 3444 2431 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2391 3356 2431 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2391 3268 2431 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2391 3180 2431 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2391 3092 2431 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2391 3004 2431 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2310 3620 2350 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2310 3532 2350 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2310 3444 2350 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2310 3356 2350 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2310 3268 2350 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2310 3180 2350 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2310 3092 2350 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2310 3004 2350 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2229 3620 2269 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2229 3532 2269 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2229 3444 2269 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2229 3356 2269 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2229 3268 2269 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2229 3180 2269 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2229 3092 2269 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2229 3004 2269 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2148 3620 2188 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2148 3532 2188 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2148 3444 2188 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2148 3356 2188 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2148 3268 2188 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2148 3180 2188 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2148 3092 2188 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2148 3004 2188 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2067 3620 2107 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2067 3532 2107 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2067 3444 2107 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2067 3356 2107 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2067 3268 2107 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2067 3180 2107 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2067 3092 2107 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 2067 3004 2107 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1986 3620 2026 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1986 3532 2026 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1986 3444 2026 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1986 3356 2026 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1986 3268 2026 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1986 3180 2026 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1986 3092 2026 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1986 3004 2026 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1905 3620 1945 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1905 3532 1945 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1905 3444 1945 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1905 3356 1945 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1905 3268 1945 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1905 3180 1945 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1905 3092 1945 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1905 3004 1945 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1824 3620 1864 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1824 3532 1864 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1824 3444 1864 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1824 3356 1864 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1824 3268 1864 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1824 3180 1864 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1824 3092 1864 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1824 3004 1864 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1743 3620 1783 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1743 3532 1783 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1743 3444 1783 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1743 3356 1783 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1743 3268 1783 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1743 3180 1783 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1743 3092 1783 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1743 3004 1783 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1662 3620 1702 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1662 3532 1702 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1662 3444 1702 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1662 3356 1702 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1662 3268 1702 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1662 3180 1702 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1662 3092 1702 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1662 3004 1702 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1581 3620 1621 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1581 3532 1621 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1581 3444 1621 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1581 3356 1621 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1581 3268 1621 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1581 3180 1621 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1581 3092 1621 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1581 3004 1621 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1500 3620 1540 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1500 3532 1540 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1500 3444 1540 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1500 3356 1540 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1500 3268 1540 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1500 3180 1540 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1500 3092 1540 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1500 3004 1540 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1419 3620 1459 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1419 3532 1459 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1419 3444 1459 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1419 3356 1459 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1419 3268 1459 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1419 3180 1459 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1419 3092 1459 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1419 3004 1459 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1338 3620 1378 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1338 3532 1378 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1338 3444 1378 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1338 3356 1378 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1338 3268 1378 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1338 3180 1378 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1338 3092 1378 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1338 3004 1378 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1257 3620 1297 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1257 3532 1297 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1257 3444 1297 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1257 3356 1297 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1257 3268 1297 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1257 3180 1297 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1257 3092 1297 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1257 3004 1297 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1176 3620 1216 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1176 3532 1216 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1176 3444 1216 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1176 3356 1216 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1176 3268 1216 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1176 3180 1216 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1176 3092 1216 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1176 3004 1216 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1095 3620 1135 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1095 3532 1135 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1095 3444 1135 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1095 3356 1135 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1095 3268 1135 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1095 3180 1135 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1095 3092 1135 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1095 3004 1135 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1014 3620 1054 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1014 3532 1054 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1014 3444 1054 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1014 3356 1054 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1014 3268 1054 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1014 3180 1054 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1014 3092 1054 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 1014 3004 1054 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 933 3620 973 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 933 3532 973 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 933 3444 973 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 933 3356 973 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 933 3268 973 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 933 3180 973 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 933 3092 973 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 933 3004 973 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 852 3620 892 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 852 3532 892 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 852 3444 892 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 852 3356 892 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 852 3268 892 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 852 3180 892 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 852 3092 892 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 852 3004 892 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 771 3620 811 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 771 3532 811 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 771 3444 811 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 771 3356 811 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 771 3268 811 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 771 3180 811 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 771 3092 811 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 771 3004 811 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 690 3620 730 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 690 3532 730 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 690 3444 730 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 690 3356 730 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 690 3268 730 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 690 3180 730 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 690 3092 730 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 690 3004 730 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 609 3620 649 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 609 3532 649 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 609 3444 649 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 609 3356 649 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 609 3268 649 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 609 3180 649 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 609 3092 649 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 609 3004 649 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 527 3620 567 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 527 3532 567 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 527 3444 567 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 527 3356 567 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 527 3268 567 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 527 3180 567 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 527 3092 567 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 527 3004 567 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 445 3620 485 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 445 3532 485 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 445 3444 485 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 445 3356 485 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 445 3268 485 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 445 3180 485 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 445 3092 485 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 445 3004 485 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 363 3620 403 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 363 3532 403 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 363 3444 403 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 363 3356 403 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 363 3268 403 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 363 3180 403 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 363 3092 403 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 363 3004 403 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 281 3620 321 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 281 3532 321 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 281 3444 321 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 281 3356 321 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 281 3268 321 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 281 3180 321 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 281 3092 321 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 281 3004 321 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 199 3620 239 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 199 3532 239 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 199 3444 239 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 199 3356 239 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 199 3268 239 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 199 3180 239 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 199 3092 239 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 199 3004 239 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 117 3620 157 3660 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 117 3532 157 3572 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 117 3444 157 3484 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 117 3356 157 3396 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 117 3268 157 3308 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 117 3180 157 3220 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 117 3092 157 3132 6 VDDA
port 5 nsew power bidirectional
rlabel metal3 s 117 3004 157 3044 6 VDDA
port 5 nsew power bidirectional
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 6 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 6 nsew ground bidirectional
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 6 nsew ground bidirectional
rlabel metal4 s 0 8317 254 9247 6 VSSD
port 6 nsew ground bidirectional
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 6 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 6 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 6 nsew ground bidirectional
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 6 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 6 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 6 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal4 s 14746 5167 15000 6097 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal4 s 0 35157 254 40000 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 40000 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 40000 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal4 s 14746 5167 15000 6097 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 40000 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal4 s 14746 5167 15000 6097 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 7 nsew ground bidirectional
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 3957 254 4887 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal4 s 14746 11647 15000 12537 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal4 s 0 11647 254 12537 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal4 s 14746 11647 15000 12537 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal4 s 14746 11647 15000 12537 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal4 s 0 12817 254 13707 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal4 s 0 10625 15000 11221 6 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 14746 10625 15000 11221 6 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 14746 10625 15000 11221 6 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 14746 10625 15000 11221 6 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 0 9673 15000 10269 6 AMUXBUS_B
port 12 nsew signal bidirectional
rlabel metal4 s 0 9673 254 10269 6 AMUXBUS_B
port 12 nsew signal bidirectional
rlabel metal4 s 14746 9673 15000 10269 6 AMUXBUS_B
port 12 nsew signal bidirectional
rlabel metal4 s 14746 9673 15000 10269 6 AMUXBUS_B
port 12 nsew signal bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 15000 40000
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 607034
string GDS_START 538154
<< end >>
