magic
tech sky130A
magscale 1 2
timestamp 1640697850
use sky130_fd_pr__hvdftpl1s2__example_55959141808506  sky130_fd_pr__hvdftpl1s2__example_55959141808506_0
timestamp 1640697850
transform 1 0 320 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808316  sky130_fd_pr__hvdfl1sd2__example_55959141808316_0
timestamp 1640697850
transform 1 0 132 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808137  sky130_fd_pr__hvdfl1sd__example_55959141808137_0
timestamp 1640697850
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 450 97 450 97 0 FreeSans 300 0 0 0 S
flabel comment s 160 97 160 97 0 FreeSans 300 0 0 0 D
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 48478706
string GDS_START 48477004
<< end >>
