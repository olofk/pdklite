magic
tech sky130A
magscale 1 2
timestamp 1640697850
<< nwell >>
rect -520 1854 3426 1950
rect -520 1552 374 1854
rect 658 1768 3338 1854
rect 3396 1768 3426 1854
rect 658 1552 4208 1768
rect -520 1076 1616 1552
rect -520 774 1743 1076
rect -520 526 616 774
<< pwell >>
rect -506 262 -420 465
rect 606 262 692 466
rect -506 -390 692 262
rect -506 -420 -420 -390
rect 606 -419 692 -390
<< mvnmos >>
rect -319 -364 -199 236
rect -143 -364 -23 236
rect 33 -364 153 236
rect 209 -364 329 236
rect 385 -364 505 236
<< mvpmos >>
rect -313 1218 -213 1818
rect -157 1218 -57 1818
rect -1 1218 99 1818
rect 155 1218 255 1818
rect 777 1618 877 1818
rect 933 1618 1133 1818
rect 1189 1618 1389 1818
rect 1563 1618 2363 1818
rect 2419 1618 3219 1818
rect 3289 1618 4089 1702
rect 777 1089 877 1289
rect 933 1089 1133 1289
rect 1189 1089 1389 1289
<< mvndiff >>
rect -372 158 -319 236
rect -372 124 -364 158
rect -330 124 -319 158
rect -372 90 -319 124
rect -372 56 -364 90
rect -330 56 -319 90
rect -372 22 -319 56
rect -372 -12 -364 22
rect -330 -12 -319 22
rect -372 -46 -319 -12
rect -372 -80 -364 -46
rect -330 -80 -319 -46
rect -372 -114 -319 -80
rect -372 -148 -364 -114
rect -330 -148 -319 -114
rect -372 -182 -319 -148
rect -372 -216 -364 -182
rect -330 -216 -319 -182
rect -372 -250 -319 -216
rect -372 -284 -364 -250
rect -330 -284 -319 -250
rect -372 -318 -319 -284
rect -372 -352 -364 -318
rect -330 -352 -319 -318
rect -372 -364 -319 -352
rect -199 158 -143 236
rect -199 124 -188 158
rect -154 124 -143 158
rect -199 90 -143 124
rect -199 56 -188 90
rect -154 56 -143 90
rect -199 22 -143 56
rect -199 -12 -188 22
rect -154 -12 -143 22
rect -199 -46 -143 -12
rect -199 -80 -188 -46
rect -154 -80 -143 -46
rect -199 -114 -143 -80
rect -199 -148 -188 -114
rect -154 -148 -143 -114
rect -199 -182 -143 -148
rect -199 -216 -188 -182
rect -154 -216 -143 -182
rect -199 -250 -143 -216
rect -199 -284 -188 -250
rect -154 -284 -143 -250
rect -199 -318 -143 -284
rect -199 -352 -188 -318
rect -154 -352 -143 -318
rect -199 -364 -143 -352
rect -23 158 33 236
rect -23 124 -12 158
rect 22 124 33 158
rect -23 90 33 124
rect -23 56 -12 90
rect 22 56 33 90
rect -23 22 33 56
rect -23 -12 -12 22
rect 22 -12 33 22
rect -23 -46 33 -12
rect -23 -80 -12 -46
rect 22 -80 33 -46
rect -23 -114 33 -80
rect -23 -148 -12 -114
rect 22 -148 33 -114
rect -23 -182 33 -148
rect -23 -216 -12 -182
rect 22 -216 33 -182
rect -23 -250 33 -216
rect -23 -284 -12 -250
rect 22 -284 33 -250
rect -23 -318 33 -284
rect -23 -352 -12 -318
rect 22 -352 33 -318
rect -23 -364 33 -352
rect 153 158 209 236
rect 153 124 164 158
rect 198 124 209 158
rect 153 90 209 124
rect 153 56 164 90
rect 198 56 209 90
rect 153 22 209 56
rect 153 -12 164 22
rect 198 -12 209 22
rect 153 -46 209 -12
rect 153 -80 164 -46
rect 198 -80 209 -46
rect 153 -114 209 -80
rect 153 -148 164 -114
rect 198 -148 209 -114
rect 153 -182 209 -148
rect 153 -216 164 -182
rect 198 -216 209 -182
rect 153 -250 209 -216
rect 153 -284 164 -250
rect 198 -284 209 -250
rect 153 -318 209 -284
rect 153 -352 164 -318
rect 198 -352 209 -318
rect 153 -364 209 -352
rect 329 158 385 236
rect 329 124 340 158
rect 374 124 385 158
rect 329 90 385 124
rect 329 56 340 90
rect 374 56 385 90
rect 329 22 385 56
rect 329 -12 340 22
rect 374 -12 385 22
rect 329 -46 385 -12
rect 329 -80 340 -46
rect 374 -80 385 -46
rect 329 -114 385 -80
rect 329 -148 340 -114
rect 374 -148 385 -114
rect 329 -182 385 -148
rect 329 -216 340 -182
rect 374 -216 385 -182
rect 329 -250 385 -216
rect 329 -284 340 -250
rect 374 -284 385 -250
rect 329 -318 385 -284
rect 329 -352 340 -318
rect 374 -352 385 -318
rect 329 -364 385 -352
rect 505 158 558 236
rect 505 124 516 158
rect 550 124 558 158
rect 505 90 558 124
rect 505 56 516 90
rect 550 56 558 90
rect 505 22 558 56
rect 505 -12 516 22
rect 550 -12 558 22
rect 505 -46 558 -12
rect 505 -80 516 -46
rect 550 -80 558 -46
rect 505 -114 558 -80
rect 505 -148 516 -114
rect 550 -148 558 -114
rect 505 -182 558 -148
rect 505 -216 516 -182
rect 550 -216 558 -182
rect 505 -250 558 -216
rect 505 -284 516 -250
rect 550 -284 558 -250
rect 505 -318 558 -284
rect 505 -352 516 -318
rect 550 -352 558 -318
rect 505 -364 558 -352
<< mvpdiff >>
rect -366 1806 -313 1818
rect -366 1772 -358 1806
rect -324 1772 -313 1806
rect -366 1738 -313 1772
rect -366 1704 -358 1738
rect -324 1704 -313 1738
rect -366 1670 -313 1704
rect -366 1636 -358 1670
rect -324 1636 -313 1670
rect -366 1602 -313 1636
rect -366 1568 -358 1602
rect -324 1568 -313 1602
rect -366 1534 -313 1568
rect -366 1500 -358 1534
rect -324 1500 -313 1534
rect -366 1466 -313 1500
rect -366 1432 -358 1466
rect -324 1432 -313 1466
rect -366 1398 -313 1432
rect -366 1364 -358 1398
rect -324 1364 -313 1398
rect -366 1330 -313 1364
rect -366 1296 -358 1330
rect -324 1296 -313 1330
rect -366 1218 -313 1296
rect -213 1806 -157 1818
rect -213 1772 -202 1806
rect -168 1772 -157 1806
rect -213 1738 -157 1772
rect -213 1704 -202 1738
rect -168 1704 -157 1738
rect -213 1670 -157 1704
rect -213 1636 -202 1670
rect -168 1636 -157 1670
rect -213 1602 -157 1636
rect -213 1568 -202 1602
rect -168 1568 -157 1602
rect -213 1534 -157 1568
rect -213 1500 -202 1534
rect -168 1500 -157 1534
rect -213 1466 -157 1500
rect -213 1432 -202 1466
rect -168 1432 -157 1466
rect -213 1398 -157 1432
rect -213 1364 -202 1398
rect -168 1364 -157 1398
rect -213 1330 -157 1364
rect -213 1296 -202 1330
rect -168 1296 -157 1330
rect -213 1218 -157 1296
rect -57 1806 -1 1818
rect -57 1772 -46 1806
rect -12 1772 -1 1806
rect -57 1738 -1 1772
rect -57 1704 -46 1738
rect -12 1704 -1 1738
rect -57 1670 -1 1704
rect -57 1636 -46 1670
rect -12 1636 -1 1670
rect -57 1602 -1 1636
rect -57 1568 -46 1602
rect -12 1568 -1 1602
rect -57 1534 -1 1568
rect -57 1500 -46 1534
rect -12 1500 -1 1534
rect -57 1466 -1 1500
rect -57 1432 -46 1466
rect -12 1432 -1 1466
rect -57 1398 -1 1432
rect -57 1364 -46 1398
rect -12 1364 -1 1398
rect -57 1330 -1 1364
rect -57 1296 -46 1330
rect -12 1296 -1 1330
rect -57 1218 -1 1296
rect 99 1806 155 1818
rect 99 1772 110 1806
rect 144 1772 155 1806
rect 99 1738 155 1772
rect 99 1704 110 1738
rect 144 1704 155 1738
rect 99 1670 155 1704
rect 99 1636 110 1670
rect 144 1636 155 1670
rect 99 1602 155 1636
rect 99 1568 110 1602
rect 144 1568 155 1602
rect 99 1534 155 1568
rect 99 1500 110 1534
rect 144 1500 155 1534
rect 99 1466 155 1500
rect 99 1432 110 1466
rect 144 1432 155 1466
rect 99 1398 155 1432
rect 99 1364 110 1398
rect 144 1364 155 1398
rect 99 1330 155 1364
rect 99 1296 110 1330
rect 144 1296 155 1330
rect 99 1218 155 1296
rect 255 1806 308 1818
rect 255 1772 266 1806
rect 300 1772 308 1806
rect 255 1738 308 1772
rect 255 1704 266 1738
rect 300 1704 308 1738
rect 255 1670 308 1704
rect 255 1636 266 1670
rect 300 1636 308 1670
rect 255 1602 308 1636
rect 724 1806 777 1818
rect 724 1772 732 1806
rect 766 1772 777 1806
rect 724 1738 777 1772
rect 724 1704 732 1738
rect 766 1704 777 1738
rect 724 1670 777 1704
rect 724 1636 732 1670
rect 766 1636 777 1670
rect 724 1618 777 1636
rect 877 1806 933 1818
rect 877 1772 888 1806
rect 922 1772 933 1806
rect 877 1738 933 1772
rect 877 1704 888 1738
rect 922 1704 933 1738
rect 877 1670 933 1704
rect 877 1636 888 1670
rect 922 1636 933 1670
rect 877 1618 933 1636
rect 1133 1806 1189 1818
rect 1133 1772 1144 1806
rect 1178 1772 1189 1806
rect 1133 1738 1189 1772
rect 1133 1704 1144 1738
rect 1178 1704 1189 1738
rect 1133 1670 1189 1704
rect 1133 1636 1144 1670
rect 1178 1636 1189 1670
rect 1133 1618 1189 1636
rect 1389 1806 1442 1818
rect 1389 1772 1400 1806
rect 1434 1772 1442 1806
rect 1389 1738 1442 1772
rect 1389 1704 1400 1738
rect 1434 1704 1442 1738
rect 1389 1670 1442 1704
rect 1389 1636 1400 1670
rect 1434 1636 1442 1670
rect 1389 1618 1442 1636
rect 1510 1800 1563 1818
rect 1510 1766 1518 1800
rect 1552 1766 1563 1800
rect 1510 1732 1563 1766
rect 1510 1698 1518 1732
rect 1552 1698 1563 1732
rect 1510 1664 1563 1698
rect 1510 1630 1518 1664
rect 1552 1630 1563 1664
rect 1510 1618 1563 1630
rect 2363 1800 2419 1818
rect 2363 1766 2374 1800
rect 2408 1766 2419 1800
rect 2363 1732 2419 1766
rect 2363 1698 2374 1732
rect 2408 1698 2419 1732
rect 2363 1664 2419 1698
rect 2363 1630 2374 1664
rect 2408 1630 2419 1664
rect 2363 1618 2419 1630
rect 3219 1800 3272 1818
rect 3219 1766 3230 1800
rect 3264 1766 3272 1800
rect 3219 1732 3272 1766
rect 3219 1698 3230 1732
rect 3264 1702 3272 1732
rect 3264 1698 3289 1702
rect 3219 1664 3289 1698
rect 3219 1630 3230 1664
rect 3264 1630 3289 1664
rect 3219 1618 3289 1630
rect 4089 1664 4142 1702
rect 4089 1630 4100 1664
rect 4134 1630 4142 1664
rect 4089 1618 4142 1630
rect 255 1568 266 1602
rect 300 1568 308 1602
rect 255 1534 308 1568
rect 255 1500 266 1534
rect 300 1500 308 1534
rect 255 1466 308 1500
rect 255 1432 266 1466
rect 300 1432 308 1466
rect 255 1398 308 1432
rect 255 1364 266 1398
rect 300 1364 308 1398
rect 255 1330 308 1364
rect 255 1296 266 1330
rect 300 1296 308 1330
rect 255 1218 308 1296
rect 724 1277 777 1289
rect 724 1243 732 1277
rect 766 1243 777 1277
rect 724 1209 777 1243
rect 724 1175 732 1209
rect 766 1175 777 1209
rect 724 1141 777 1175
rect 724 1107 732 1141
rect 766 1107 777 1141
rect 724 1089 777 1107
rect 877 1277 933 1289
rect 877 1243 888 1277
rect 922 1243 933 1277
rect 877 1209 933 1243
rect 877 1175 888 1209
rect 922 1175 933 1209
rect 877 1141 933 1175
rect 877 1107 888 1141
rect 922 1107 933 1141
rect 877 1089 933 1107
rect 1133 1277 1189 1289
rect 1133 1243 1144 1277
rect 1178 1243 1189 1277
rect 1133 1209 1189 1243
rect 1133 1175 1144 1209
rect 1178 1175 1189 1209
rect 1133 1141 1189 1175
rect 1133 1107 1144 1141
rect 1178 1107 1189 1141
rect 1133 1089 1189 1107
rect 1389 1277 1442 1289
rect 1389 1243 1400 1277
rect 1434 1243 1442 1277
rect 1389 1209 1442 1243
rect 1389 1175 1400 1209
rect 1434 1175 1442 1209
rect 1389 1141 1442 1175
rect 1389 1107 1400 1141
rect 1434 1107 1442 1141
rect 1389 1089 1442 1107
<< mvndiffc >>
rect -364 124 -330 158
rect -364 56 -330 90
rect -364 -12 -330 22
rect -364 -80 -330 -46
rect -364 -148 -330 -114
rect -364 -216 -330 -182
rect -364 -284 -330 -250
rect -364 -352 -330 -318
rect -188 124 -154 158
rect -188 56 -154 90
rect -188 -12 -154 22
rect -188 -80 -154 -46
rect -188 -148 -154 -114
rect -188 -216 -154 -182
rect -188 -284 -154 -250
rect -188 -352 -154 -318
rect -12 124 22 158
rect -12 56 22 90
rect -12 -12 22 22
rect -12 -80 22 -46
rect -12 -148 22 -114
rect -12 -216 22 -182
rect -12 -284 22 -250
rect -12 -352 22 -318
rect 164 124 198 158
rect 164 56 198 90
rect 164 -12 198 22
rect 164 -80 198 -46
rect 164 -148 198 -114
rect 164 -216 198 -182
rect 164 -284 198 -250
rect 164 -352 198 -318
rect 340 124 374 158
rect 340 56 374 90
rect 340 -12 374 22
rect 340 -80 374 -46
rect 340 -148 374 -114
rect 340 -216 374 -182
rect 340 -284 374 -250
rect 340 -352 374 -318
rect 516 124 550 158
rect 516 56 550 90
rect 516 -12 550 22
rect 516 -80 550 -46
rect 516 -148 550 -114
rect 516 -216 550 -182
rect 516 -284 550 -250
rect 516 -352 550 -318
<< mvpdiffc >>
rect -358 1772 -324 1806
rect -358 1704 -324 1738
rect -358 1636 -324 1670
rect -358 1568 -324 1602
rect -358 1500 -324 1534
rect -358 1432 -324 1466
rect -358 1364 -324 1398
rect -358 1296 -324 1330
rect -202 1772 -168 1806
rect -202 1704 -168 1738
rect -202 1636 -168 1670
rect -202 1568 -168 1602
rect -202 1500 -168 1534
rect -202 1432 -168 1466
rect -202 1364 -168 1398
rect -202 1296 -168 1330
rect -46 1772 -12 1806
rect -46 1704 -12 1738
rect -46 1636 -12 1670
rect -46 1568 -12 1602
rect -46 1500 -12 1534
rect -46 1432 -12 1466
rect -46 1364 -12 1398
rect -46 1296 -12 1330
rect 110 1772 144 1806
rect 110 1704 144 1738
rect 110 1636 144 1670
rect 110 1568 144 1602
rect 110 1500 144 1534
rect 110 1432 144 1466
rect 110 1364 144 1398
rect 110 1296 144 1330
rect 266 1772 300 1806
rect 266 1704 300 1738
rect 266 1636 300 1670
rect 732 1772 766 1806
rect 732 1704 766 1738
rect 732 1636 766 1670
rect 888 1772 922 1806
rect 888 1704 922 1738
rect 888 1636 922 1670
rect 1144 1772 1178 1806
rect 1144 1704 1178 1738
rect 1144 1636 1178 1670
rect 1400 1772 1434 1806
rect 1400 1704 1434 1738
rect 1400 1636 1434 1670
rect 1518 1766 1552 1800
rect 1518 1698 1552 1732
rect 1518 1630 1552 1664
rect 2374 1766 2408 1800
rect 2374 1698 2408 1732
rect 2374 1630 2408 1664
rect 3230 1766 3264 1800
rect 3230 1698 3264 1732
rect 3230 1630 3264 1664
rect 4100 1630 4134 1664
rect 266 1568 300 1602
rect 266 1500 300 1534
rect 266 1432 300 1466
rect 266 1364 300 1398
rect 266 1296 300 1330
rect 732 1243 766 1277
rect 732 1175 766 1209
rect 732 1107 766 1141
rect 888 1243 922 1277
rect 888 1175 922 1209
rect 888 1107 922 1141
rect 1144 1243 1178 1277
rect 1144 1175 1178 1209
rect 1144 1107 1178 1141
rect 1400 1243 1434 1277
rect 1400 1175 1434 1209
rect 1400 1107 1434 1141
<< mvpsubdiff >>
rect -480 405 -446 439
rect 632 406 666 440
rect -480 337 -446 371
rect -480 269 -446 303
rect 632 338 666 372
rect 632 270 666 304
rect -480 201 -446 235
rect -480 133 -446 167
rect -480 65 -446 99
rect -480 -3 -446 31
rect -480 -71 -446 -37
rect -480 -139 -446 -105
rect -480 -207 -446 -173
rect -480 -275 -446 -241
rect -480 -394 -446 -309
rect 632 202 666 236
rect 632 134 666 168
rect 632 66 666 100
rect 632 -2 666 32
rect 632 -70 666 -36
rect 632 -138 666 -104
rect 632 -206 666 -172
rect 632 -274 666 -240
rect 632 -393 666 -308
<< mvnsubdiff >>
rect -454 1794 -420 1818
rect -454 1722 -420 1760
rect -454 1650 -420 1688
rect -454 1578 -420 1616
rect -454 1506 -420 1544
rect -454 1434 -420 1472
rect -454 1362 -420 1400
rect -454 1290 -420 1328
rect -454 1218 -420 1256
rect 512 1228 546 1252
rect -454 1147 -420 1184
rect -454 1090 -420 1113
rect 512 1157 546 1194
rect -454 1076 -334 1090
rect -420 1066 -334 1076
rect -420 1042 -368 1066
rect -454 1032 -368 1042
rect -454 1005 -334 1032
rect -420 971 -334 1005
rect -454 952 -334 971
rect -454 934 -368 952
rect -420 918 -368 934
rect -420 900 -334 918
rect -454 894 -334 900
rect -192 1060 -158 1084
rect -192 980 -158 1026
rect -192 900 -158 946
rect -454 863 -420 894
rect -454 792 -420 829
rect -454 721 -420 758
rect -454 650 -420 687
rect -454 592 -420 616
rect -16 1060 18 1084
rect -16 952 18 1026
rect -16 894 18 918
rect 160 1060 194 1084
rect 160 980 194 1026
rect 160 900 194 946
rect -192 820 -158 866
rect -192 741 -158 786
rect -192 662 -158 707
rect -192 604 -158 628
rect 336 1066 370 1090
rect 336 952 370 1032
rect 336 894 370 918
rect 512 1086 546 1123
rect 512 1015 546 1052
rect 546 981 580 1010
rect 512 944 580 981
rect 546 910 580 944
rect 160 820 194 866
rect 160 741 194 786
rect 160 662 194 707
rect 160 604 194 628
rect 512 873 580 910
rect 546 840 580 873
rect 1022 976 1057 1010
rect 1091 976 1126 1010
rect 1160 976 1195 1010
rect 1229 976 1264 1010
rect 1298 976 1333 1010
rect 1367 976 1402 1010
rect 1436 976 1471 1010
rect 1505 976 1540 1010
rect 1574 976 1609 1010
rect 1643 976 1682 1010
rect 1022 942 1682 976
rect 1022 908 1057 942
rect 1091 908 1126 942
rect 1160 908 1195 942
rect 1229 908 1264 942
rect 1298 908 1333 942
rect 1367 908 1402 942
rect 1436 908 1471 942
rect 1505 908 1540 942
rect 1574 908 1609 942
rect 1643 908 1682 942
rect 1022 874 1682 908
rect 1022 840 1057 874
rect 1091 840 1126 874
rect 1160 840 1195 874
rect 1229 840 1264 874
rect 1298 840 1333 874
rect 1367 840 1402 874
rect 1436 840 1471 874
rect 1505 840 1540 874
rect 1574 840 1609 874
rect 1643 848 1682 874
rect 1643 840 1677 848
rect 512 802 546 839
rect 512 732 546 768
rect 512 662 546 698
rect 512 604 546 628
<< mvpsubdiffcont >>
rect -480 371 -446 405
rect -480 303 -446 337
rect -480 235 -446 269
rect 632 372 666 406
rect 632 304 666 338
rect 632 236 666 270
rect -480 167 -446 201
rect -480 99 -446 133
rect -480 31 -446 65
rect -480 -37 -446 -3
rect -480 -105 -446 -71
rect -480 -173 -446 -139
rect -480 -241 -446 -207
rect -480 -309 -446 -275
rect 632 168 666 202
rect 632 100 666 134
rect 632 32 666 66
rect 632 -36 666 -2
rect 632 -104 666 -70
rect 632 -172 666 -138
rect 632 -240 666 -206
rect 632 -308 666 -274
<< mvnsubdiffcont >>
rect -454 1760 -420 1794
rect -454 1688 -420 1722
rect -454 1616 -420 1650
rect -454 1544 -420 1578
rect -454 1472 -420 1506
rect -454 1400 -420 1434
rect -454 1328 -420 1362
rect -454 1256 -420 1290
rect -454 1184 -420 1218
rect -454 1113 -420 1147
rect 512 1194 546 1228
rect 512 1123 546 1157
rect -454 1042 -420 1076
rect -368 1032 -334 1066
rect -454 971 -420 1005
rect -454 900 -420 934
rect -368 918 -334 952
rect -192 1026 -158 1060
rect -192 946 -158 980
rect -454 829 -420 863
rect -454 758 -420 792
rect -454 687 -420 721
rect -454 616 -420 650
rect -192 866 -158 900
rect -16 1026 18 1060
rect -16 918 18 952
rect 160 1026 194 1060
rect 160 946 194 980
rect -192 786 -158 820
rect -192 707 -158 741
rect -192 628 -158 662
rect 160 866 194 900
rect 336 1032 370 1066
rect 336 918 370 952
rect 512 1052 546 1086
rect 512 981 546 1015
rect 512 910 546 944
rect 160 786 194 820
rect 160 707 194 741
rect 160 628 194 662
rect 512 839 546 873
rect 580 840 1022 1010
rect 1057 976 1091 1010
rect 1126 976 1160 1010
rect 1195 976 1229 1010
rect 1264 976 1298 1010
rect 1333 976 1367 1010
rect 1402 976 1436 1010
rect 1471 976 1505 1010
rect 1540 976 1574 1010
rect 1609 976 1643 1010
rect 1057 908 1091 942
rect 1126 908 1160 942
rect 1195 908 1229 942
rect 1264 908 1298 942
rect 1333 908 1367 942
rect 1402 908 1436 942
rect 1471 908 1505 942
rect 1540 908 1574 942
rect 1609 908 1643 942
rect 1057 840 1091 874
rect 1126 840 1160 874
rect 1195 840 1229 874
rect 1264 840 1298 874
rect 1333 840 1367 874
rect 1402 840 1436 874
rect 1471 840 1505 874
rect 1540 840 1574 874
rect 1609 840 1643 874
rect 512 768 546 802
rect 512 698 546 732
rect 512 628 546 662
<< poly >>
rect -313 1900 255 1916
rect -313 1866 -282 1900
rect -248 1866 -214 1900
rect -180 1866 -146 1900
rect -112 1866 -78 1900
rect -44 1866 -10 1900
rect 24 1866 58 1900
rect 92 1866 126 1900
rect 160 1866 194 1900
rect 228 1866 255 1900
rect -313 1844 255 1866
rect 681 1900 877 1916
rect 681 1866 697 1900
rect 731 1866 827 1900
rect 861 1866 877 1900
rect 681 1850 877 1866
rect -313 1818 -213 1844
rect -157 1818 -57 1844
rect -1 1818 99 1844
rect 155 1818 255 1844
rect 777 1818 877 1850
rect 933 1900 1389 1916
rect 933 1866 949 1900
rect 983 1866 1027 1900
rect 1061 1866 1105 1900
rect 1139 1866 1183 1900
rect 1217 1866 1261 1900
rect 1295 1866 1339 1900
rect 1373 1866 1389 1900
rect 933 1844 1389 1866
rect 933 1818 1133 1844
rect 1189 1818 1389 1844
rect 1563 1900 2363 1916
rect 1563 1866 1611 1900
rect 1645 1866 1679 1900
rect 1713 1866 1747 1900
rect 1781 1866 1815 1900
rect 1849 1866 1883 1900
rect 1917 1866 1951 1900
rect 1985 1866 2019 1900
rect 2053 1866 2087 1900
rect 2121 1866 2155 1900
rect 2189 1866 2223 1900
rect 2257 1866 2291 1900
rect 2325 1866 2363 1900
rect 1563 1818 2363 1866
rect 2419 1900 3219 1916
rect 2419 1866 2450 1900
rect 2484 1866 2518 1900
rect 2552 1866 2586 1900
rect 2620 1866 2654 1900
rect 2688 1866 2722 1900
rect 2756 1866 2790 1900
rect 2824 1866 2858 1900
rect 2892 1866 2926 1900
rect 2960 1866 2994 1900
rect 3028 1866 3062 1900
rect 3096 1866 3130 1900
rect 3164 1866 3219 1900
rect 2419 1818 3219 1866
rect 3289 1784 4089 1800
rect 3289 1750 3321 1784
rect 3355 1750 3395 1784
rect 3429 1750 3469 1784
rect 3503 1750 3544 1784
rect 3578 1750 3619 1784
rect 3653 1750 3694 1784
rect 3728 1750 3769 1784
rect 3803 1750 3844 1784
rect 3878 1750 3919 1784
rect 3953 1750 3994 1784
rect 4028 1750 4089 1784
rect 3289 1702 4089 1750
rect 777 1592 877 1618
rect 933 1592 1133 1618
rect 1189 1592 1389 1618
rect 1563 1592 2363 1618
rect 2419 1592 3219 1618
rect 3289 1592 4089 1618
rect 677 1421 877 1437
rect 677 1387 693 1421
rect 727 1387 827 1421
rect 861 1387 877 1421
rect 677 1371 877 1387
rect 777 1289 877 1371
rect 933 1421 1389 1437
rect 933 1387 949 1421
rect 983 1387 1027 1421
rect 1061 1387 1105 1421
rect 1139 1387 1183 1421
rect 1217 1387 1261 1421
rect 1295 1387 1339 1421
rect 1373 1387 1389 1421
rect 933 1315 1389 1387
rect 933 1289 1133 1315
rect 1189 1289 1389 1315
rect -313 1202 -213 1218
rect -157 1202 -57 1218
rect -1 1202 99 1218
rect 155 1202 255 1218
rect -313 1158 255 1202
rect -313 1124 -271 1158
rect -237 1124 -203 1158
rect -169 1124 -135 1158
rect -101 1124 -67 1158
rect -33 1124 1 1158
rect 35 1124 69 1158
rect 103 1124 137 1158
rect 171 1124 205 1158
rect 239 1124 255 1158
rect -313 1108 255 1124
rect 777 1063 877 1089
rect 933 1063 1133 1089
rect 1189 1063 1389 1089
rect -319 386 -199 402
rect -319 352 -276 386
rect -242 352 -199 386
rect -319 318 -199 352
rect -319 284 -276 318
rect -242 284 -199 318
rect -319 236 -199 284
rect -143 386 -23 402
rect -143 352 -100 386
rect -66 352 -23 386
rect -143 318 -23 352
rect -143 284 -100 318
rect -66 284 -23 318
rect -143 236 -23 284
rect 33 386 153 402
rect 33 352 76 386
rect 110 352 153 386
rect 33 318 153 352
rect 33 284 76 318
rect 110 284 153 318
rect 33 236 153 284
rect 209 386 329 402
rect 209 352 252 386
rect 286 352 329 386
rect 209 318 329 352
rect 209 284 252 318
rect 286 284 329 318
rect 209 236 329 284
rect 385 386 505 402
rect 385 352 428 386
rect 462 352 505 386
rect 385 318 505 352
rect 385 284 428 318
rect 462 284 505 318
rect 385 236 505 284
rect -319 -390 -199 -364
rect -143 -390 -23 -364
rect 33 -390 153 -364
rect 209 -390 329 -364
rect 385 -390 505 -364
<< polycont >>
rect -282 1866 -248 1900
rect -214 1866 -180 1900
rect -146 1866 -112 1900
rect -78 1866 -44 1900
rect -10 1866 24 1900
rect 58 1866 92 1900
rect 126 1866 160 1900
rect 194 1866 228 1900
rect 697 1866 731 1900
rect 827 1866 861 1900
rect 949 1866 983 1900
rect 1027 1866 1061 1900
rect 1105 1866 1139 1900
rect 1183 1866 1217 1900
rect 1261 1866 1295 1900
rect 1339 1866 1373 1900
rect 1611 1866 1645 1900
rect 1679 1866 1713 1900
rect 1747 1866 1781 1900
rect 1815 1866 1849 1900
rect 1883 1866 1917 1900
rect 1951 1866 1985 1900
rect 2019 1866 2053 1900
rect 2087 1866 2121 1900
rect 2155 1866 2189 1900
rect 2223 1866 2257 1900
rect 2291 1866 2325 1900
rect 2450 1866 2484 1900
rect 2518 1866 2552 1900
rect 2586 1866 2620 1900
rect 2654 1866 2688 1900
rect 2722 1866 2756 1900
rect 2790 1866 2824 1900
rect 2858 1866 2892 1900
rect 2926 1866 2960 1900
rect 2994 1866 3028 1900
rect 3062 1866 3096 1900
rect 3130 1866 3164 1900
rect 3321 1750 3355 1784
rect 3395 1750 3429 1784
rect 3469 1750 3503 1784
rect 3544 1750 3578 1784
rect 3619 1750 3653 1784
rect 3694 1750 3728 1784
rect 3769 1750 3803 1784
rect 3844 1750 3878 1784
rect 3919 1750 3953 1784
rect 3994 1750 4028 1784
rect 693 1387 727 1421
rect 827 1387 861 1421
rect 949 1387 983 1421
rect 1027 1387 1061 1421
rect 1105 1387 1139 1421
rect 1183 1387 1217 1421
rect 1261 1387 1295 1421
rect 1339 1387 1373 1421
rect -271 1124 -237 1158
rect -203 1124 -169 1158
rect -135 1124 -101 1158
rect -67 1124 -33 1158
rect 1 1124 35 1158
rect 69 1124 103 1158
rect 137 1124 171 1158
rect 205 1124 239 1158
rect -276 352 -242 386
rect -276 284 -242 318
rect -100 352 -66 386
rect -100 284 -66 318
rect 76 352 110 386
rect 76 284 110 318
rect 252 352 286 386
rect 252 284 286 318
rect 428 352 462 386
rect 428 284 462 318
<< locali >>
rect -265 1900 -227 1901
rect -193 1900 -155 1901
rect -121 1900 -83 1901
rect -49 1900 -11 1901
rect 23 1900 61 1901
rect 95 1900 133 1901
rect 167 1900 205 1901
rect 1621 1900 1659 1901
rect 1693 1900 1731 1901
rect 1765 1900 1803 1901
rect 1837 1900 1875 1901
rect 1909 1900 1947 1901
rect 1981 1900 2019 1901
rect 2053 1900 2091 1901
rect 2125 1900 2163 1901
rect 2197 1900 2235 1901
rect 2269 1900 2307 1901
rect -248 1867 -227 1900
rect -180 1867 -155 1900
rect -112 1867 -83 1900
rect -44 1867 -11 1900
rect -298 1866 -282 1867
rect -248 1866 -214 1867
rect -180 1866 -146 1867
rect -112 1866 -78 1867
rect -44 1866 -10 1867
rect 24 1866 58 1900
rect 95 1867 126 1900
rect 167 1867 194 1900
rect 239 1867 244 1900
rect 92 1866 126 1867
rect 160 1866 194 1867
rect 228 1866 244 1867
rect 681 1866 697 1900
rect 731 1866 827 1900
rect 861 1866 877 1900
rect 933 1866 949 1900
rect 983 1866 1027 1900
rect 1061 1866 1105 1900
rect 1139 1866 1183 1900
rect 1217 1866 1261 1900
rect 1295 1866 1339 1900
rect 1373 1866 1389 1900
rect 1645 1867 1659 1900
rect 1713 1867 1731 1900
rect 1781 1867 1803 1900
rect 1849 1867 1875 1900
rect 1917 1867 1947 1900
rect 1595 1866 1611 1867
rect 1645 1866 1679 1867
rect 1713 1866 1747 1867
rect 1781 1866 1815 1867
rect 1849 1866 1883 1867
rect 1917 1866 1951 1867
rect 1985 1866 2019 1900
rect 2053 1866 2087 1900
rect 2125 1867 2155 1900
rect 2197 1867 2223 1900
rect 2269 1867 2291 1900
rect 2465 1900 2503 1901
rect 2537 1900 2575 1901
rect 2609 1900 2647 1901
rect 2681 1900 2719 1901
rect 2753 1900 2791 1901
rect 2825 1900 2863 1901
rect 2897 1900 2935 1901
rect 2969 1900 3007 1901
rect 3041 1900 3079 1901
rect 3113 1900 3151 1901
rect 2484 1867 2503 1900
rect 2552 1867 2575 1900
rect 2620 1867 2647 1900
rect 2688 1867 2719 1900
rect 2121 1866 2155 1867
rect 2189 1866 2223 1867
rect 2257 1866 2291 1867
rect 2325 1866 2341 1867
rect 2434 1866 2450 1867
rect 2484 1866 2518 1867
rect 2552 1866 2586 1867
rect 2620 1866 2654 1867
rect 2688 1866 2722 1867
rect 2756 1866 2790 1900
rect 2825 1867 2858 1900
rect 2897 1867 2926 1900
rect 2969 1867 2994 1900
rect 3041 1867 3062 1900
rect 3113 1867 3130 1900
rect 3185 1867 3368 1901
rect 2824 1866 2858 1867
rect 2892 1866 2926 1867
rect 2960 1866 2994 1867
rect 3028 1866 3062 1867
rect 3096 1866 3130 1867
rect 3164 1866 3368 1867
rect -454 1794 -420 1818
rect -454 1728 -420 1760
rect -454 1656 -420 1688
rect -454 1578 -420 1616
rect -454 1506 -420 1544
rect -454 1434 -420 1472
rect -454 1362 -420 1400
rect -454 1290 -420 1328
rect -454 1218 -420 1256
rect -358 1806 -324 1822
rect -358 1738 -324 1772
rect -358 1670 -324 1704
rect -358 1602 -324 1636
rect -358 1534 -324 1568
rect -358 1466 -324 1500
rect -202 1806 -168 1822
rect -202 1738 -168 1772
rect -202 1670 -168 1704
rect -202 1602 -168 1636
rect -202 1534 -168 1568
rect -202 1494 -168 1500
rect -46 1806 -12 1822
rect -46 1738 -12 1772
rect -46 1670 -12 1704
rect -46 1602 -12 1636
rect -46 1534 -12 1568
rect -202 1466 -164 1494
rect -358 1398 -324 1432
rect -358 1330 -324 1364
rect -358 1246 -324 1296
rect -168 1460 -164 1466
rect -46 1466 -12 1500
rect -202 1398 -168 1432
rect -202 1330 -168 1364
rect -202 1280 -168 1296
rect -46 1398 -12 1432
rect -46 1330 -12 1364
rect 110 1806 144 1822
rect 110 1738 144 1772
rect 110 1670 144 1704
rect 110 1602 144 1636
rect 110 1534 144 1568
rect 110 1466 144 1500
rect 110 1398 144 1432
rect 110 1330 144 1364
rect -46 1246 -12 1296
rect 266 1806 300 1822
rect 266 1738 300 1772
rect 494 1806 766 1822
rect 494 1772 732 1806
rect 494 1738 766 1772
rect 266 1670 300 1704
rect 266 1602 300 1636
rect 376 1652 410 1690
rect 494 1704 732 1738
rect 494 1670 766 1704
rect 494 1636 732 1670
rect 494 1620 766 1636
rect 266 1534 300 1568
rect 266 1466 300 1500
rect 266 1398 300 1432
rect 266 1330 300 1364
rect 144 1296 148 1321
rect 110 1287 148 1296
rect 110 1280 144 1287
rect 266 1246 300 1296
rect 494 1321 600 1620
rect 800 1421 851 1866
rect 888 1806 922 1822
rect 968 1816 1098 1866
rect 968 1782 982 1816
rect 1016 1782 1054 1816
rect 1088 1782 1098 1816
rect 1133 1806 1189 1822
rect 888 1738 922 1772
rect 888 1670 922 1690
rect 970 1421 1066 1782
rect 1133 1772 1144 1806
rect 1178 1772 1189 1806
rect 1224 1816 1354 1866
rect 1224 1782 1236 1816
rect 1270 1782 1308 1816
rect 1342 1782 1354 1816
rect 1400 1806 1434 1822
rect 1133 1738 1189 1772
rect 1133 1704 1144 1738
rect 1178 1704 1189 1738
rect 1133 1670 1189 1704
rect 1133 1636 1144 1670
rect 1178 1636 1189 1670
rect 1133 1494 1189 1636
rect 1138 1460 1176 1494
rect 1248 1421 1353 1782
rect 1510 1800 1548 1816
rect 1510 1782 1518 1800
rect 2370 1800 2408 1820
rect 2370 1786 2374 1800
rect 1400 1738 1434 1772
rect 1400 1670 1434 1690
rect 1518 1732 1552 1766
rect 1518 1664 1552 1698
rect 1518 1614 1552 1630
rect 3230 1800 3264 1816
rect 2374 1732 2408 1766
rect 3301 1784 3368 1866
rect 4100 1820 4186 1910
rect 4114 1786 4152 1820
rect 3230 1732 3264 1766
rect 3305 1750 3321 1784
rect 3355 1750 3395 1784
rect 3429 1750 3469 1784
rect 3503 1750 3544 1784
rect 3578 1750 3619 1784
rect 3653 1750 3694 1784
rect 3728 1750 3769 1784
rect 3803 1750 3844 1784
rect 3878 1750 3919 1784
rect 3953 1750 3994 1784
rect 4028 1750 4044 1784
rect 2374 1664 2408 1698
rect 2374 1614 2408 1630
rect 4100 1664 4186 1786
rect 4134 1630 4186 1664
rect 4100 1613 4186 1630
rect 677 1387 693 1421
rect 727 1387 827 1421
rect 861 1387 877 1421
rect 677 1369 877 1387
rect 933 1387 949 1421
rect 983 1387 1027 1421
rect 1061 1387 1105 1421
rect 1139 1387 1183 1421
rect 1217 1387 1261 1421
rect 1295 1387 1339 1421
rect 1373 1387 1389 1421
rect 933 1369 1389 1387
rect 528 1287 566 1321
rect 729 1287 767 1321
rect 732 1277 766 1287
rect -358 1238 300 1246
rect -324 1204 -286 1238
rect -252 1204 -214 1238
rect -180 1204 -142 1238
rect -108 1204 -70 1238
rect -36 1204 2 1238
rect 36 1204 74 1238
rect 108 1204 146 1238
rect 180 1204 218 1238
rect 252 1212 300 1238
rect 512 1228 546 1252
rect -454 1147 -420 1184
rect -287 1124 -271 1158
rect -234 1124 -203 1158
rect -159 1124 -135 1158
rect -84 1124 -67 1158
rect -9 1124 1 1158
rect 66 1124 69 1158
rect 103 1124 108 1158
rect 171 1124 184 1158
rect 239 1124 260 1158
rect 294 1124 336 1158
rect 370 1124 412 1158
rect 446 1124 462 1158
rect -454 1090 -420 1113
rect -454 1078 -334 1090
rect -420 1042 -368 1078
rect -454 1032 -368 1042
rect -454 1006 -334 1032
rect -420 972 -368 1006
rect -420 971 -334 972
rect -454 952 -334 971
rect -454 934 -368 952
rect -420 900 -368 934
rect -454 894 -334 900
rect -454 863 -420 894
rect -454 792 -420 829
rect -454 721 -420 758
rect -454 650 -420 687
rect -454 592 -420 616
rect -382 854 -310 860
rect -382 820 -368 854
rect -334 820 -310 854
rect -382 782 -310 820
rect -382 748 -368 782
rect -334 748 -310 782
rect -484 480 -450 518
rect -484 439 -450 446
rect -484 408 -446 439
rect -450 405 -446 408
rect -484 371 -480 374
rect -484 337 -446 371
rect -484 303 -480 337
rect -484 269 -446 303
rect -484 236 -480 269
rect -480 201 -446 235
rect -480 133 -446 167
rect -480 65 -446 99
rect -480 -3 -446 31
rect -480 -71 -446 -37
rect -480 -139 -446 -105
rect -480 -207 -446 -173
rect -480 -275 -446 -241
rect -480 -394 -446 -309
rect -382 158 -310 748
rect -276 386 -242 1124
rect -192 1078 -158 1084
rect -192 1006 -158 1026
rect -192 934 -158 946
rect -192 820 -158 866
rect -192 741 -158 786
rect -192 662 -158 707
rect -192 604 -158 628
rect -276 318 -242 352
rect -276 268 -242 284
rect -200 552 -134 564
rect -200 518 -184 552
rect -150 518 -134 552
rect -200 480 -134 518
rect -200 446 -184 480
rect -150 446 -134 480
rect -200 408 -134 446
rect -200 374 -184 408
rect -150 374 -134 408
rect -382 124 -364 158
rect -330 124 -310 158
rect -382 90 -310 124
rect -382 56 -364 90
rect -330 56 -310 90
rect -382 22 -310 56
rect -382 -12 -364 22
rect -330 -12 -310 22
rect -382 -46 -310 -12
rect -382 -80 -364 -46
rect -330 -80 -310 -46
rect -382 -114 -310 -80
rect -382 -148 -364 -114
rect -330 -148 -310 -114
rect -382 -182 -310 -148
rect -382 -216 -364 -182
rect -330 -216 -310 -182
rect -382 -250 -310 -216
rect -382 -284 -364 -250
rect -330 -284 -310 -250
rect -382 -318 -310 -284
rect -382 -352 -364 -318
rect -330 -352 -310 -318
rect -382 -368 -310 -352
rect -200 158 -134 374
rect -100 386 -66 1124
rect -16 1078 18 1084
rect -16 1006 18 1026
rect -16 952 18 972
rect -16 894 18 900
rect -100 318 -66 352
rect -100 268 -66 284
rect -32 854 42 860
rect -32 820 -16 854
rect 18 820 42 854
rect -32 782 42 820
rect -32 748 -16 782
rect 18 748 42 782
rect -200 124 -188 158
rect -154 124 -134 158
rect -200 90 -134 124
rect -200 56 -188 90
rect -154 56 -134 90
rect -200 22 -134 56
rect -200 -12 -188 22
rect -154 -12 -134 22
rect -200 -46 -134 -12
rect -200 -80 -188 -46
rect -154 -80 -134 -46
rect -200 -114 -134 -80
rect -200 -148 -188 -114
rect -154 -148 -134 -114
rect -200 -182 -134 -148
rect -200 -216 -188 -182
rect -154 -216 -134 -182
rect -200 -250 -134 -216
rect -200 -284 -188 -250
rect -154 -284 -134 -250
rect -200 -318 -134 -284
rect -200 -352 -188 -318
rect -154 -352 -134 -318
rect -200 -368 -134 -352
rect -32 158 42 748
rect 76 386 110 1124
rect 160 1078 194 1084
rect 160 1006 194 1026
rect 160 934 194 946
rect 160 820 194 866
rect 160 741 194 786
rect 160 662 194 707
rect 160 604 194 628
rect 76 318 110 352
rect 76 268 110 284
rect 152 552 218 564
rect 152 518 168 552
rect 202 518 218 552
rect 152 480 218 518
rect 152 446 168 480
rect 202 446 218 480
rect 152 408 218 446
rect 152 374 168 408
rect 202 374 218 408
rect -32 124 -12 158
rect 22 124 42 158
rect -32 90 42 124
rect -32 56 -12 90
rect 22 56 42 90
rect -32 22 42 56
rect -32 -12 -12 22
rect 22 -12 42 22
rect -32 -46 42 -12
rect -32 -80 -12 -46
rect 22 -80 42 -46
rect -32 -114 42 -80
rect -32 -148 -12 -114
rect 22 -148 42 -114
rect -32 -182 42 -148
rect -32 -216 -12 -182
rect 22 -216 42 -182
rect -32 -250 42 -216
rect -32 -284 -12 -250
rect 22 -284 42 -250
rect -32 -318 42 -284
rect -32 -352 -12 -318
rect 22 -352 42 -318
rect -32 -368 42 -352
rect 152 158 218 374
rect 252 386 286 1124
rect 336 1078 370 1090
rect 336 1006 370 1032
rect 336 952 370 972
rect 336 894 370 900
rect 252 318 286 352
rect 252 268 286 284
rect 320 854 394 860
rect 320 820 336 854
rect 370 820 394 854
rect 320 782 394 820
rect 320 748 336 782
rect 370 748 394 782
rect 152 124 164 158
rect 198 124 218 158
rect 152 90 218 124
rect 152 56 164 90
rect 198 56 218 90
rect 152 22 218 56
rect 152 -12 164 22
rect 198 -12 218 22
rect 152 -46 218 -12
rect 152 -80 164 -46
rect 198 -80 218 -46
rect 152 -114 218 -80
rect 152 -148 164 -114
rect 198 -148 218 -114
rect 152 -182 218 -148
rect 152 -216 164 -182
rect 198 -216 218 -182
rect 152 -250 218 -216
rect 152 -284 164 -250
rect 198 -284 218 -250
rect 152 -318 218 -284
rect 152 -352 164 -318
rect 198 -352 218 -318
rect 152 -368 218 -352
rect 320 158 394 748
rect 428 386 462 1124
rect 512 1157 546 1194
rect 512 1086 546 1123
rect 732 1209 766 1243
rect 732 1141 766 1175
rect 732 1091 766 1107
rect 888 1277 922 1293
rect 1146 1287 1184 1321
rect 888 1209 922 1243
rect 888 1147 922 1175
rect 512 1015 546 1052
rect 888 1075 922 1107
rect 1144 1277 1178 1287
rect 1144 1209 1178 1243
rect 1144 1141 1178 1175
rect 1144 1091 1178 1107
rect 1400 1277 1434 1293
rect 1400 1209 1434 1243
rect 1400 1147 1434 1175
rect 888 1010 922 1041
rect 1400 1075 1434 1107
rect 1400 1010 1434 1041
rect 1677 1010 1684 1252
rect 546 1002 580 1010
rect 1022 1002 1057 1010
rect 1091 1002 1126 1010
rect 1160 1002 1195 1010
rect 1229 1002 1264 1010
rect 1298 1002 1333 1010
rect 1367 1002 1402 1010
rect 1436 1002 1471 1010
rect 1505 1002 1540 1010
rect 1574 1002 1609 1010
rect 512 944 516 981
rect 512 896 516 910
rect 1229 976 1237 1002
rect 1298 976 1310 1002
rect 1367 976 1383 1002
rect 1436 976 1456 1002
rect 1505 976 1529 1002
rect 1574 976 1602 1002
rect 1643 976 1684 1010
rect 1198 968 1237 976
rect 1271 968 1310 976
rect 1344 968 1383 976
rect 1417 968 1456 976
rect 1490 968 1529 976
rect 1563 968 1602 976
rect 1636 968 1684 976
rect 1198 942 1684 968
rect 1229 930 1264 942
rect 1298 930 1333 942
rect 1367 930 1402 942
rect 1436 930 1471 942
rect 1505 930 1540 942
rect 1574 930 1609 942
rect 1229 908 1237 930
rect 1298 908 1310 930
rect 1367 908 1383 930
rect 1436 908 1456 930
rect 1505 908 1529 930
rect 1574 908 1602 930
rect 1643 908 1684 942
rect 1198 896 1237 908
rect 1271 896 1310 908
rect 1344 896 1383 908
rect 1417 896 1456 908
rect 1490 896 1529 908
rect 1563 896 1602 908
rect 1636 896 1684 908
rect 512 873 580 896
rect 546 840 580 873
rect 1022 874 1684 896
rect 1022 840 1057 874
rect 1091 840 1126 874
rect 1160 840 1195 874
rect 1229 840 1264 874
rect 1298 840 1333 874
rect 1367 840 1402 874
rect 1436 840 1471 874
rect 1505 840 1540 874
rect 1574 840 1609 874
rect 1643 840 1684 874
rect 512 802 546 839
rect 512 732 546 768
rect 512 662 546 698
rect 512 604 546 628
rect 428 318 462 352
rect 428 268 462 284
rect 500 552 675 564
rect 500 518 506 552
rect 540 518 630 552
rect 664 518 675 552
rect 500 480 675 518
rect 500 446 506 480
rect 540 446 630 480
rect 664 446 675 480
rect 500 408 675 446
rect 500 374 506 408
rect 540 374 630 408
rect 664 406 675 408
rect 500 372 632 374
rect 666 372 675 406
rect 500 338 675 372
rect 500 304 632 338
rect 666 304 675 338
rect 500 270 675 304
rect 320 124 340 158
rect 374 124 394 158
rect 320 90 394 124
rect 320 56 340 90
rect 374 56 394 90
rect 320 22 394 56
rect 320 -12 340 22
rect 374 -12 394 22
rect 320 -46 394 -12
rect 320 -80 340 -46
rect 374 -80 394 -46
rect 320 -114 394 -80
rect 320 -148 340 -114
rect 374 -148 394 -114
rect 320 -182 394 -148
rect 320 -216 340 -182
rect 374 -216 394 -182
rect 320 -250 394 -216
rect 320 -284 340 -250
rect 374 -284 394 -250
rect 320 -318 394 -284
rect 320 -352 340 -318
rect 374 -352 394 -318
rect 320 -368 394 -352
rect 500 236 632 270
rect 666 236 675 270
rect 500 202 675 236
rect 500 168 632 202
rect 666 168 675 202
rect 500 158 675 168
rect 500 124 516 158
rect 550 134 675 158
rect 550 124 632 134
rect 500 100 632 124
rect 666 100 675 134
rect 500 90 675 100
rect 500 56 516 90
rect 550 66 675 90
rect 550 56 632 66
rect 500 32 632 56
rect 666 32 675 66
rect 500 22 675 32
rect 500 -12 516 22
rect 550 -2 675 22
rect 550 -12 632 -2
rect 500 -36 632 -12
rect 666 -36 675 -2
rect 500 -46 675 -36
rect 500 -80 516 -46
rect 550 -70 675 -46
rect 550 -80 632 -70
rect 500 -104 632 -80
rect 666 -104 675 -70
rect 500 -114 675 -104
rect 500 -148 516 -114
rect 550 -138 675 -114
rect 550 -148 632 -138
rect 500 -172 632 -148
rect 666 -172 675 -138
rect 500 -182 675 -172
rect 500 -216 516 -182
rect 550 -206 675 -182
rect 550 -216 632 -206
rect 500 -240 632 -216
rect 666 -240 675 -206
rect 500 -250 675 -240
rect 500 -284 516 -250
rect 550 -274 675 -250
rect 550 -284 632 -274
rect 500 -308 632 -284
rect 666 -308 675 -274
rect 500 -318 675 -308
rect 500 -352 516 -318
rect 550 -352 675 -318
rect 500 -394 675 -352
<< viali >>
rect -299 1900 -265 1901
rect -227 1900 -193 1901
rect -155 1900 -121 1901
rect -83 1900 -49 1901
rect -11 1900 23 1901
rect 61 1900 95 1901
rect 133 1900 167 1901
rect 205 1900 239 1901
rect 1587 1900 1621 1901
rect 1659 1900 1693 1901
rect 1731 1900 1765 1901
rect 1803 1900 1837 1901
rect 1875 1900 1909 1901
rect 1947 1900 1981 1901
rect 2019 1900 2053 1901
rect 2091 1900 2125 1901
rect 2163 1900 2197 1901
rect 2235 1900 2269 1901
rect 2307 1900 2341 1901
rect -299 1867 -282 1900
rect -282 1867 -265 1900
rect -227 1867 -214 1900
rect -214 1867 -193 1900
rect -155 1867 -146 1900
rect -146 1867 -121 1900
rect -83 1867 -78 1900
rect -78 1867 -49 1900
rect -11 1867 -10 1900
rect -10 1867 23 1900
rect 61 1867 92 1900
rect 92 1867 95 1900
rect 133 1867 160 1900
rect 160 1867 167 1900
rect 205 1867 228 1900
rect 228 1867 239 1900
rect 1587 1867 1611 1900
rect 1611 1867 1621 1900
rect 1659 1867 1679 1900
rect 1679 1867 1693 1900
rect 1731 1867 1747 1900
rect 1747 1867 1765 1900
rect 1803 1867 1815 1900
rect 1815 1867 1837 1900
rect 1875 1867 1883 1900
rect 1883 1867 1909 1900
rect 1947 1867 1951 1900
rect 1951 1867 1981 1900
rect 2019 1867 2053 1900
rect 2091 1867 2121 1900
rect 2121 1867 2125 1900
rect 2163 1867 2189 1900
rect 2189 1867 2197 1900
rect 2235 1867 2257 1900
rect 2257 1867 2269 1900
rect 2307 1867 2325 1900
rect 2325 1867 2341 1900
rect 2431 1900 2465 1901
rect 2503 1900 2537 1901
rect 2575 1900 2609 1901
rect 2647 1900 2681 1901
rect 2719 1900 2753 1901
rect 2791 1900 2825 1901
rect 2863 1900 2897 1901
rect 2935 1900 2969 1901
rect 3007 1900 3041 1901
rect 3079 1900 3113 1901
rect 3151 1900 3185 1901
rect 2431 1867 2450 1900
rect 2450 1867 2465 1900
rect 2503 1867 2518 1900
rect 2518 1867 2537 1900
rect 2575 1867 2586 1900
rect 2586 1867 2609 1900
rect 2647 1867 2654 1900
rect 2654 1867 2681 1900
rect 2719 1867 2722 1900
rect 2722 1867 2753 1900
rect 2791 1867 2824 1900
rect 2824 1867 2825 1900
rect 2863 1867 2892 1900
rect 2892 1867 2897 1900
rect 2935 1867 2960 1900
rect 2960 1867 2969 1900
rect 3007 1867 3028 1900
rect 3028 1867 3041 1900
rect 3079 1867 3096 1900
rect 3096 1867 3113 1900
rect 3151 1867 3164 1900
rect 3164 1867 3185 1900
rect -454 1722 -420 1728
rect -454 1694 -420 1722
rect -454 1650 -420 1656
rect -454 1622 -420 1650
rect -236 1460 -202 1494
rect -164 1460 -130 1494
rect 76 1287 110 1321
rect 376 1690 410 1724
rect 376 1618 410 1652
rect 148 1287 182 1321
rect 982 1782 1016 1816
rect 1054 1782 1088 1816
rect 888 1704 922 1724
rect 888 1690 922 1704
rect 888 1636 922 1652
rect 888 1618 922 1636
rect 1236 1782 1270 1816
rect 1308 1782 1342 1816
rect 1104 1460 1138 1494
rect 1176 1460 1210 1494
rect 1476 1782 1510 1816
rect 1548 1800 1582 1816
rect 1548 1782 1552 1800
rect 1552 1782 1582 1800
rect 2336 1786 2370 1820
rect 1400 1704 1434 1724
rect 1400 1690 1434 1704
rect 1400 1636 1434 1652
rect 1400 1618 1434 1636
rect 2408 1786 2442 1820
rect 4080 1786 4114 1820
rect 4152 1786 4186 1820
rect 3158 1698 3230 1720
rect 3230 1698 3264 1720
rect 3158 1664 3264 1698
rect 3158 1630 3230 1664
rect 3230 1630 3264 1664
rect 3158 1614 3264 1630
rect 494 1287 528 1321
rect 566 1287 600 1321
rect 695 1287 729 1321
rect 767 1287 801 1321
rect -358 1204 -324 1238
rect -286 1204 -252 1238
rect -214 1204 -180 1238
rect -142 1204 -108 1238
rect -70 1204 -36 1238
rect 2 1204 36 1238
rect 74 1204 108 1238
rect 146 1204 180 1238
rect 218 1204 252 1238
rect -268 1124 -237 1158
rect -237 1124 -234 1158
rect -193 1124 -169 1158
rect -169 1124 -159 1158
rect -118 1124 -101 1158
rect -101 1124 -84 1158
rect -43 1124 -33 1158
rect -33 1124 -9 1158
rect 32 1124 35 1158
rect 35 1124 66 1158
rect 108 1124 137 1158
rect 137 1124 142 1158
rect 184 1124 205 1158
rect 205 1124 218 1158
rect 260 1124 294 1158
rect 336 1124 370 1158
rect 412 1124 446 1158
rect -454 1076 -420 1078
rect -454 1044 -420 1076
rect -368 1066 -334 1078
rect -368 1044 -334 1066
rect -454 1005 -420 1006
rect -454 972 -420 1005
rect -368 972 -334 1006
rect -454 900 -420 934
rect -368 918 -334 934
rect -368 900 -334 918
rect -368 820 -334 854
rect -368 748 -334 782
rect -484 518 -450 552
rect -484 446 -450 480
rect -484 405 -450 408
rect -484 374 -480 405
rect -480 374 -450 405
rect -192 1060 -158 1078
rect -192 1044 -158 1060
rect -192 980 -158 1006
rect -192 972 -158 980
rect -192 900 -158 934
rect -184 518 -150 552
rect -184 446 -150 480
rect -184 374 -150 408
rect -16 1060 18 1078
rect -16 1044 18 1060
rect -16 972 18 1006
rect -16 918 18 934
rect -16 900 18 918
rect -16 820 18 854
rect -16 748 18 782
rect 160 1060 194 1078
rect 160 1044 194 1060
rect 160 980 194 1006
rect 160 972 194 980
rect 160 900 194 934
rect 168 518 202 552
rect 168 446 202 480
rect 168 374 202 408
rect 336 1066 370 1078
rect 336 1044 370 1066
rect 336 972 370 1006
rect 336 918 370 934
rect 336 900 370 918
rect 336 820 370 854
rect 336 748 370 782
rect 1112 1287 1146 1321
rect 1184 1287 1218 1321
rect 888 1141 922 1147
rect 888 1113 922 1141
rect 1400 1141 1434 1147
rect 1400 1113 1434 1141
rect 888 1041 922 1075
rect 1400 1041 1434 1075
rect 516 981 546 1002
rect 546 981 580 1002
rect 516 944 580 981
rect 516 910 546 944
rect 546 910 580 944
rect 516 896 580 910
rect 580 896 1022 1002
rect 1022 976 1057 1002
rect 1057 976 1091 1002
rect 1091 976 1126 1002
rect 1126 976 1160 1002
rect 1160 976 1195 1002
rect 1195 976 1198 1002
rect 1237 976 1264 1002
rect 1264 976 1271 1002
rect 1310 976 1333 1002
rect 1333 976 1344 1002
rect 1383 976 1402 1002
rect 1402 976 1417 1002
rect 1456 976 1471 1002
rect 1471 976 1490 1002
rect 1529 976 1540 1002
rect 1540 976 1563 1002
rect 1602 976 1609 1002
rect 1609 976 1636 1002
rect 1022 942 1198 976
rect 1237 968 1271 976
rect 1310 968 1344 976
rect 1383 968 1417 976
rect 1456 968 1490 976
rect 1529 968 1563 976
rect 1602 968 1636 976
rect 1022 908 1057 942
rect 1057 908 1091 942
rect 1091 908 1126 942
rect 1126 908 1160 942
rect 1160 908 1195 942
rect 1195 908 1198 942
rect 1237 908 1264 930
rect 1264 908 1271 930
rect 1310 908 1333 930
rect 1333 908 1344 930
rect 1383 908 1402 930
rect 1402 908 1417 930
rect 1456 908 1471 930
rect 1471 908 1490 930
rect 1529 908 1540 930
rect 1540 908 1563 930
rect 1602 908 1609 930
rect 1609 908 1636 930
rect 1022 896 1198 908
rect 1237 896 1271 908
rect 1310 896 1344 908
rect 1383 896 1417 908
rect 1456 896 1490 908
rect 1529 896 1563 908
rect 1602 896 1636 908
rect 506 518 540 552
rect 630 518 664 552
rect 506 446 540 480
rect 630 446 664 480
rect 506 374 540 408
rect 630 406 664 408
rect 630 374 632 406
rect 632 374 664 406
<< metal1 >>
rect -827 1861 -821 1913
rect -769 1861 -757 1913
rect -705 1901 2353 1913
rect -705 1867 -299 1901
rect -265 1867 -227 1901
rect -193 1867 -155 1901
rect -121 1867 -83 1901
rect -49 1867 -11 1901
rect 23 1867 61 1901
rect 95 1867 133 1901
rect 167 1867 205 1901
rect 239 1867 1587 1901
rect 1621 1867 1659 1901
rect 1693 1867 1731 1901
rect 1765 1867 1803 1901
rect 1837 1867 1875 1901
rect 1909 1867 1947 1901
rect 1981 1867 2019 1901
rect 2053 1867 2091 1901
rect 2125 1867 2163 1901
rect 2197 1867 2235 1901
rect 2269 1867 2307 1901
rect 2341 1867 2353 1901
rect -705 1861 2353 1867
rect 2408 1861 2414 1913
rect 2466 1861 2478 1913
rect 2530 1901 3197 1913
rect 2537 1867 2575 1901
rect 2609 1867 2647 1901
rect 2681 1867 2719 1901
rect 2753 1867 2791 1901
rect 2825 1867 2863 1901
rect 2897 1867 2935 1901
rect 2969 1867 3007 1901
rect 3041 1867 3079 1901
rect 3113 1867 3151 1901
rect 3185 1867 3197 1901
rect 2530 1861 3197 1867
rect 970 1816 1354 1822
rect 970 1782 982 1816
rect 1016 1782 1054 1816
rect 1088 1782 1236 1816
rect 1270 1782 1308 1816
rect 1342 1782 1354 1816
rect 970 1776 1354 1782
rect 1464 1776 1470 1828
rect 1522 1776 1534 1828
rect 1586 1776 1594 1828
rect 2324 1820 4198 1826
rect 2324 1786 2336 1820
rect 2370 1786 2408 1820
rect 2442 1786 4080 1820
rect 4114 1786 4152 1820
rect 4186 1786 4198 1820
rect 2324 1780 4198 1786
rect -520 1728 3426 1748
rect -520 1694 -454 1728
rect -420 1724 3426 1728
rect -420 1694 376 1724
rect -520 1690 376 1694
rect 410 1690 888 1724
rect 922 1690 1400 1724
rect 1434 1720 3426 1724
rect 1434 1690 3158 1720
rect -520 1656 3158 1690
rect -520 1622 -454 1656
rect -420 1652 3158 1656
rect -420 1622 376 1652
rect -520 1618 376 1622
rect 410 1618 888 1652
rect 922 1618 1400 1652
rect 1434 1618 3158 1652
rect -520 1614 3158 1618
rect 3264 1614 3426 1720
rect -520 1602 3426 1614
rect -248 1494 1516 1500
rect -248 1460 -236 1494
rect -202 1460 -164 1494
rect -130 1460 1104 1494
rect 1138 1460 1176 1494
rect 1210 1460 1516 1494
rect -248 1454 1516 1460
tri 1455 1428 1481 1454 ne
tri 1450 1327 1481 1358 se
rect 1481 1327 1516 1454
rect 64 1321 825 1327
rect 64 1287 76 1321
rect 110 1287 148 1321
rect 182 1287 494 1321
rect 528 1287 566 1321
rect 600 1287 695 1321
rect 729 1287 767 1321
rect 801 1287 825 1321
rect 64 1281 825 1287
rect 1098 1321 1516 1327
rect 1098 1287 1112 1321
rect 1146 1287 1184 1321
rect 1218 1287 1516 1321
rect 1098 1281 1516 1287
rect -751 1240 -699 1246
tri -699 1238 -691 1246 sw
rect -370 1238 1470 1250
rect -699 1204 -691 1238
tri -691 1204 -657 1238 sw
rect -370 1204 -358 1238
rect -324 1204 -286 1238
rect -252 1204 -214 1238
rect -180 1204 -142 1238
rect -108 1204 -70 1238
rect -36 1204 2 1238
rect 36 1204 74 1238
rect 108 1204 146 1238
rect 180 1204 218 1238
rect 252 1204 1470 1238
rect -699 1198 -657 1204
tri -657 1198 -651 1204 sw
rect -370 1198 1470 1204
rect 1522 1198 1534 1250
rect 1586 1198 1592 1250
rect 2408 1240 2460 1246
rect -699 1189 -651 1198
tri -651 1189 -642 1198 sw
rect -699 1188 -642 1189
rect -751 1176 -642 1188
rect -699 1170 -642 1176
tri -642 1170 -623 1189 sw
tri 2389 1170 2408 1189 se
rect 2408 1176 2460 1188
rect -699 1158 458 1170
tri 2383 1164 2389 1170 se
rect 2389 1164 2408 1170
rect -699 1124 -268 1158
rect -234 1124 -193 1158
rect -159 1124 -118 1158
rect -84 1124 -43 1158
rect -9 1124 32 1158
rect 66 1124 108 1158
rect 142 1124 184 1158
rect 218 1124 260 1158
rect 294 1124 336 1158
rect 370 1124 412 1158
rect 446 1124 458 1158
rect -751 1118 458 1124
rect 882 1147 1440 1159
rect 882 1113 888 1147
rect 922 1113 1400 1147
rect 1434 1113 1440 1147
rect 1527 1124 2408 1164
rect 1527 1118 2460 1124
rect -520 1078 545 1090
rect -520 1044 -454 1078
rect -420 1044 -368 1078
rect -334 1044 -192 1078
rect -158 1044 -16 1078
rect 18 1044 160 1078
rect 194 1044 336 1078
rect 370 1075 545 1078
tri 545 1075 560 1090 sw
tri 877 1075 882 1080 se
rect 882 1075 1440 1113
rect 370 1044 560 1075
rect -520 1041 560 1044
tri 560 1041 594 1075 sw
tri 858 1056 877 1075 se
rect 877 1056 888 1075
tri 843 1041 858 1056 se
rect 858 1041 888 1056
rect 922 1041 1400 1075
rect 1434 1041 1440 1075
tri 1642 1056 1676 1090 se
rect 1676 1056 3426 1090
rect -520 1010 594 1041
tri 594 1010 625 1041 sw
tri 812 1010 843 1041 se
rect 843 1010 1440 1041
tri 1440 1010 1486 1056 sw
tri 1596 1010 1642 1056 se
rect 1642 1010 3426 1056
rect -520 1006 3426 1010
rect -520 972 -454 1006
rect -420 972 -368 1006
rect -334 972 -192 1006
rect -158 972 -16 1006
rect 18 972 160 1006
rect 194 972 336 1006
rect 370 1002 3426 1006
rect 370 972 516 1002
rect -520 934 516 972
rect -520 900 -454 934
rect -420 900 -368 934
rect -334 900 -192 934
rect -158 900 -16 934
rect 18 900 160 934
rect 194 900 336 934
rect 370 900 516 934
rect -520 896 516 900
rect 1198 968 1237 1002
rect 1271 968 1310 1002
rect 1344 968 1383 1002
rect 1417 968 1456 1002
rect 1490 968 1529 1002
rect 1563 968 1602 1002
rect 1636 968 3426 1002
rect 1198 930 3426 968
rect 1198 896 1237 930
rect 1271 896 1310 930
rect 1344 896 1383 930
rect 1417 896 1456 930
rect 1490 896 1529 930
rect 1563 896 1602 930
rect 1636 896 3426 930
rect -520 888 3426 896
rect -380 854 1470 860
rect -380 820 -368 854
rect -334 820 -16 854
rect 18 820 336 854
rect 370 820 1470 854
rect -380 808 1470 820
rect 1522 808 1534 860
rect 1586 808 1592 860
rect -380 782 -282 808
tri -282 782 -256 808 nw
tri -94 782 -68 808 ne
rect -68 782 70 808
tri 70 782 96 808 nw
tri 258 782 284 808 ne
rect 284 782 382 808
rect -380 748 -368 782
rect -334 748 -316 782
tri -316 748 -282 782 nw
tri -68 748 -34 782 ne
rect -34 748 -16 782
rect 18 748 36 782
tri 36 748 70 782 nw
tri 284 748 318 782 ne
rect 318 748 336 782
rect 370 748 382 782
rect -380 742 -322 748
tri -322 742 -316 748 nw
tri -34 742 -28 748 ne
rect -28 742 30 748
tri 30 742 36 748 nw
tri 318 742 324 748 ne
rect 324 742 382 748
tri 382 742 448 808 nw
rect -520 552 3426 564
rect -520 518 -484 552
rect -450 518 -184 552
rect -150 518 168 552
rect 202 518 506 552
rect 540 518 630 552
rect 664 518 3426 552
rect -520 480 3426 518
rect -520 446 -484 480
rect -450 446 -184 480
rect -150 446 168 480
rect 202 446 506 480
rect 540 446 630 480
rect 664 446 3426 480
rect -520 408 3426 446
rect -520 374 -484 408
rect -450 374 -184 408
rect -150 374 168 408
rect 202 374 506 408
rect 540 374 630 408
rect 664 374 3426 408
rect -520 362 3426 374
<< via1 >>
rect -821 1861 -769 1913
rect -757 1861 -705 1913
rect 2414 1901 2466 1913
rect 2414 1867 2431 1901
rect 2431 1867 2465 1901
rect 2465 1867 2466 1901
rect 2414 1861 2466 1867
rect 2478 1901 2530 1913
rect 2478 1867 2503 1901
rect 2503 1867 2530 1901
rect 2478 1861 2530 1867
rect 1470 1816 1522 1828
rect 1470 1782 1476 1816
rect 1476 1782 1510 1816
rect 1510 1782 1522 1816
rect 1470 1776 1522 1782
rect 1534 1816 1586 1828
rect 1534 1782 1548 1816
rect 1548 1782 1582 1816
rect 1582 1782 1586 1816
rect 1534 1776 1586 1782
rect -751 1188 -699 1240
rect 1470 1198 1522 1250
rect 1534 1198 1586 1250
rect -751 1124 -699 1176
rect 2408 1188 2460 1240
rect 2408 1124 2460 1176
rect 1470 808 1522 860
rect 1534 808 1586 860
<< metal2 >>
rect -827 1861 -821 1913
rect -769 1861 -757 1913
rect -705 1861 -699 1913
rect -827 1240 -699 1861
rect 2408 1861 2414 1913
rect 2466 1861 2478 1913
rect 2530 1861 2536 1913
rect -827 1188 -751 1240
rect -827 1176 -699 1188
rect -827 1124 -751 1176
rect -827 1118 -699 1124
rect 1464 1776 1470 1828
rect 1522 1776 1534 1828
rect 1586 1776 1592 1828
rect 1464 1250 1592 1776
rect 1464 1198 1470 1250
rect 1522 1198 1534 1250
rect 1586 1198 1592 1250
rect 1464 860 1592 1198
rect 2408 1240 2460 1861
tri 2460 1836 2485 1861 nw
rect 2408 1176 2460 1188
rect 2408 1118 2460 1124
rect 1464 808 1470 860
rect 1522 808 1534 860
rect 1586 808 1592 860
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1640697850
transform 1 0 1464 0 -1 860
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1640697850
transform 0 1 -751 1 0 1118
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1640697850
transform 1 0 -827 0 -1 1913
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1640697850
transform 0 -1 2460 -1 0 1246
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_4
timestamp 1640697850
transform -1 0 2536 0 1 1861
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_5
timestamp 1640697850
transform 1 0 1464 0 -1 1250
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_6
timestamp 1640697850
transform -1 0 1592 0 1 1776
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808294  sky130_fd_pr__via_pol1__example_55959141808294_0
timestamp 1640697850
transform 0 -1 244 -1 0 1916
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808294  sky130_fd_pr__via_pol1__example_55959141808294_1
timestamp 1640697850
transform 0 -1 255 -1 0 1174
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_0
timestamp 1640697850
transform 0 -1 2341 1 0 1850
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_1
timestamp 1640697850
transform 0 -1 3180 1 0 1850
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1640697850
transform -1 0 -226 0 -1 402
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1640697850
transform -1 0 -50 0 -1 402
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_2
timestamp 1640697850
transform -1 0 126 0 -1 402
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_3
timestamp 1640697850
transform -1 0 302 0 -1 402
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_4
timestamp 1640697850
transform -1 0 478 0 -1 402
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_0
timestamp 1640697850
transform 1 0 336 0 -1 854
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_1
timestamp 1640697850
transform 1 0 -368 0 -1 854
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_2
timestamp 1640697850
transform 1 0 -16 0 -1 854
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_0
timestamp 1640697850
transform 0 1 3158 -1 0 1720
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808357  sky130_fd_pr__via_l1m1__example_55959141808357_0
timestamp 1640697850
transform 1 0 -358 0 1 1204
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_0
timestamp 1640697850
transform 1 0 -299 0 1 1867
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808326  sky130_fd_pr__via_l1m1__example_55959141808326_0
timestamp 1640697850
transform -1 0 3185 0 1 1867
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808326  sky130_fd_pr__via_l1m1__example_55959141808326_1
timestamp 1640697850
transform -1 0 2341 0 1 1867
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1640697850
transform 0 -1 922 -1 0 1147
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1640697850
transform -1 0 1218 0 1 1287
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1640697850
transform -1 0 801 0 1 1287
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1640697850
transform -1 0 182 0 1 1287
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1640697850
transform 0 -1 1434 -1 0 1724
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1640697850
transform 0 -1 922 -1 0 1724
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1640697850
transform -1 0 1088 0 1 1782
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1640697850
transform 0 1 -454 -1 0 1728
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1640697850
transform -1 0 1342 0 1 1782
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1640697850
transform -1 0 1582 0 1 1782
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1640697850
transform -1 0 -130 0 1 1460
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1640697850
transform -1 0 1210 0 1 1460
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_12
timestamp 1640697850
transform 0 -1 410 -1 0 1724
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_13
timestamp 1640697850
transform -1 0 600 0 1 1287
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_14
timestamp 1640697850
transform 0 -1 1434 -1 0 1147
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1640697850
transform 0 1 -454 -1 0 1078
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1640697850
transform 0 1 -368 -1 0 1078
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_2
timestamp 1640697850
transform 0 1 -16 -1 0 1078
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_3
timestamp 1640697850
transform 0 1 336 -1 0 1078
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_4
timestamp 1640697850
transform 0 1 160 -1 0 1078
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_5
timestamp 1640697850
transform 0 1 -192 -1 0 1078
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_6
timestamp 1640697850
transform 0 1 -484 -1 0 552
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_7
timestamp 1640697850
transform 0 1 -184 -1 0 552
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_8
timestamp 1640697850
transform 0 1 168 -1 0 552
box 0 0 1 1
use sky130_fd_pr__pfet_01v8__example_55959141808359  sky130_fd_pr__pfet_01v8__example_55959141808359_0
timestamp 1640697850
transform -1 0 3219 0 1 1618
box -28 0 1684 97
use sky130_fd_pr__pfet_01v8__example_55959141808355  sky130_fd_pr__pfet_01v8__example_55959141808355_0
timestamp 1640697850
transform 1 0 -1 0 -1 1818
box -28 0 284 267
use sky130_fd_pr__pfet_01v8__example_55959141808355  sky130_fd_pr__pfet_01v8__example_55959141808355_1
timestamp 1640697850
transform -1 0 -57 0 -1 1818
box -28 0 284 267
use sky130_fd_pr__pfet_01v8__example_55959141808358  sky130_fd_pr__pfet_01v8__example_55959141808358_0
timestamp 1640697850
transform 1 0 3289 0 1 1618
box -42 0 828 29
use sky130_fd_pr__pfet_01v8__example_55959141808353  sky130_fd_pr__pfet_01v8__example_55959141808353_0
timestamp 1640697850
transform -1 0 1133 0 -1 1289
box -28 0 228 97
use sky130_fd_pr__pfet_01v8__example_55959141808353  sky130_fd_pr__pfet_01v8__example_55959141808353_1
timestamp 1640697850
transform 1 0 1189 0 -1 1289
box -28 0 228 97
use sky130_fd_pr__pfet_01v8__example_55959141808353  sky130_fd_pr__pfet_01v8__example_55959141808353_2
timestamp 1640697850
transform -1 0 1133 0 -1 1818
box -28 0 228 97
use sky130_fd_pr__pfet_01v8__example_55959141808353  sky130_fd_pr__pfet_01v8__example_55959141808353_3
timestamp 1640697850
transform 1 0 1189 0 -1 1818
box -28 0 228 97
use sky130_fd_pr__pfet_01v8__example_55959141808352  sky130_fd_pr__pfet_01v8__example_55959141808352_0
timestamp 1640697850
transform 1 0 777 0 -1 1289
box -28 0 128 97
use sky130_fd_pr__pfet_01v8__example_55959141808352  sky130_fd_pr__pfet_01v8__example_55959141808352_1
timestamp 1640697850
transform 1 0 777 0 -1 1818
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808351  sky130_fd_pr__nfet_01v8__example_55959141808351_0
timestamp 1640697850
transform -1 0 505 0 1 -364
box -28 0 852 267
<< labels >>
flabel locali s 726 1373 772 1419 3 FreeSans 300 180 0 0 EN_FAST_N[0]
port 1 nsew
flabel metal1 s 3386 1602 3426 1748 7 FreeSans 300 180 0 0 VCC_IO
port 2 nsew
flabel metal1 s 3386 362 3426 564 7 FreeSans 300 180 0 0 VGND_IO
port 3 nsew
flabel metal1 s -520 1602 -480 1748 3 FreeSans 300 180 0 0 VCC_IO
port 2 nsew
flabel metal1 s -520 362 -480 564 3 FreeSans 300 180 0 0 VGND_IO
port 3 nsew
flabel metal1 s -520 888 -480 1090 3 FreeSans 300 180 0 0 VCC_IO
port 2 nsew
flabel metal1 s 3386 888 3426 1090 7 FreeSans 300 180 0 0 VCC_IO
port 2 nsew
flabel metal1 s -311 1861 -265 1913 3 FreeSans 300 180 0 0 DRVLO_H_N
port 4 nsew
flabel metal1 s 1030 1776 1078 1822 7 FreeSans 300 180 0 0 EN_FAST_N[1]
port 5 nsew
flabel metal1 s 1528 1118 1574 1164 7 FreeSans 300 180 0 0 PDEN_H_N
port 6 nsew
flabel metal1 s 505 1198 552 1250 7 FreeSans 300 180 0 0 PD_H
port 7 nsew
flabel comment s 2630 1917 2630 1917 0 FreeSans 300 0 0 0 PDEN_H_N
flabel comment s 3094 1686 3094 1686 0 FreeSans 300 0 0 0 VCC_IO
flabel comment s 45 1149 45 1149 3 FreeSans 300 180 0 0 DRVLO_H_N
flabel comment s 349 1562 349 1562 0 FreeSans 300 0 0 0 INTNR0
flabel comment s 518 1484 518 1484 0 FreeSans 300 0 0 0 INTNR1
flabel comment s -82 1232 -82 1232 0 FreeSans 300 0 0 0 PD_H
flabel comment s 16 844 16 844 0 FreeSans 300 0 0 0 PD_H
flabel comment s 1947 1924 1947 1924 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 1327 1917 1327 1917 0 FreeSans 300 0 0 0 EN_FAST_N[1]
flabel comment s 2386 1810 2386 1810 0 FreeSans 300 90 0 0 INT_SLOW
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 37044282
string GDS_START 37015112
<< end >>
