magic
tech sky130A
magscale 1 2
timestamp 1640697850
<< labels >>
flabel comment s 62 25 62 25 2 FreeSans 50 0 0 0 EM1O
flabel comment s 50 27 50 27 0 FreeSans 50 0 0 0 A
flabel comment s 86 27 86 27 0 FreeSans 50 0 0 0 B
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 39963454
string GDS_START 39962686
<< end >>
