magic
tech sky130A
magscale 1 2
timestamp 1640697850
use sky130_fd_pr__hvdfl1sd2__example_55959141808143  sky130_fd_pr__hvdfl1sd2__example_55959141808143_0
timestamp 1640697850
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808102  sky130_fd_pr__hvdfl1sd__example_55959141808102_0
timestamp 1640697850
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808102  sky130_fd_pr__hvdfl1sd__example_55959141808102_1
timestamp 1640697850
transform 1 0 296 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 324 267 324 267 0 FreeSans 300 0 0 0 S
flabel comment s 148 267 148 267 0 FreeSans 300 0 0 0 D
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 36848516
string GDS_START 36846816
<< end >>
