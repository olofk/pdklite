magic
tech sky130A
magscale 1 2
timestamp 1619729480
<< checkpaint >>
rect -1260 -853 16260 41260
<< metal3 >>
rect 106 11282 112 11346
rect 176 11282 193 11346
rect 257 11282 274 11346
rect 338 11282 355 11346
rect 419 11282 436 11346
rect 500 11282 517 11346
rect 581 11282 598 11346
rect 662 11282 679 11346
rect 743 11282 760 11346
rect 824 11282 841 11346
rect 905 11282 922 11346
rect 986 11282 1003 11346
rect 1067 11282 1084 11346
rect 1148 11282 1165 11346
rect 1229 11282 1246 11346
rect 1310 11282 1327 11346
rect 1391 11282 1408 11346
rect 1472 11282 1489 11346
rect 1553 11282 1570 11346
rect 1634 11282 1651 11346
rect 1715 11282 1732 11346
rect 1796 11282 1813 11346
rect 1877 11282 1894 11346
rect 1958 11282 1975 11346
rect 2039 11282 2056 11346
rect 2120 11282 2137 11346
rect 2201 11282 2218 11346
rect 2282 11282 2299 11346
rect 2363 11282 2380 11346
rect 2444 11282 2461 11346
rect 2525 11282 2542 11346
rect 2606 11282 2623 11346
rect 2687 11282 2704 11346
rect 2768 11282 2785 11346
rect 2849 11282 2866 11346
rect 2930 11282 2947 11346
rect 3011 11282 3028 11346
rect 3092 11282 3109 11346
rect 3173 11282 3190 11346
rect 3254 11282 3271 11346
rect 3335 11282 3352 11346
rect 3416 11282 3433 11346
rect 3497 11282 3514 11346
rect 3578 11282 3595 11346
rect 3659 11282 3676 11346
rect 3740 11282 3757 11346
rect 3821 11282 3838 11346
rect 3902 11282 3919 11346
rect 3983 11282 4000 11346
rect 4064 11282 4081 11346
rect 4145 11282 4162 11346
rect 4226 11282 4243 11346
rect 4307 11282 4324 11346
rect 4388 11282 4405 11346
rect 4469 11282 4486 11346
rect 4550 11282 4567 11346
rect 4631 11282 4648 11346
rect 4712 11282 4729 11346
rect 4793 11282 4809 11346
rect 4873 11282 4879 11346
rect 10078 11282 10084 11346
rect 10148 11282 10165 11346
rect 10229 11282 10246 11346
rect 10310 11282 10327 11346
rect 10391 11282 10408 11346
rect 10472 11282 10489 11346
rect 10553 11282 10570 11346
rect 10634 11282 10651 11346
rect 10715 11282 10732 11346
rect 10796 11282 10813 11346
rect 10877 11282 10894 11346
rect 10958 11282 10975 11346
rect 11039 11282 11056 11346
rect 11120 11282 11137 11346
rect 11201 11282 11218 11346
rect 11282 11282 11299 11346
rect 11363 11282 11380 11346
rect 11444 11282 11461 11346
rect 11525 11282 11542 11346
rect 11606 11282 11623 11346
rect 11687 11282 11704 11346
rect 11768 11282 11785 11346
rect 11849 11282 11866 11346
rect 11930 11282 11947 11346
rect 12011 11282 12028 11346
rect 12092 11282 12109 11346
rect 12173 11282 12190 11346
rect 12254 11282 12271 11346
rect 12335 11282 12352 11346
rect 12416 11282 12433 11346
rect 12497 11282 12514 11346
rect 12578 11282 12595 11346
rect 12659 11282 12676 11346
rect 12740 11282 12757 11346
rect 12821 11282 12838 11346
rect 12902 11282 12919 11346
rect 12983 11282 13000 11346
rect 13064 11282 13081 11346
rect 13145 11282 13162 11346
rect 13226 11282 13243 11346
rect 13307 11282 13324 11346
rect 13388 11282 13405 11346
rect 13469 11282 13486 11346
rect 13550 11282 13567 11346
rect 13631 11282 13648 11346
rect 13712 11282 13729 11346
rect 13793 11282 13810 11346
rect 13874 11282 13891 11346
rect 13955 11282 13972 11346
rect 14036 11282 14053 11346
rect 14117 11282 14134 11346
rect 14198 11282 14215 11346
rect 14279 11282 14296 11346
rect 14360 11282 14378 11346
rect 14442 11282 14460 11346
rect 14524 11282 14542 11346
rect 14606 11282 14624 11346
rect 14688 11282 14706 11346
rect 14770 11282 14788 11346
rect 14852 11282 14858 11346
rect 99 10563 4879 10564
rect 99 10499 105 10563
rect 169 10499 187 10563
rect 251 10499 269 10563
rect 333 10499 351 10563
rect 415 10499 433 10563
rect 497 10499 515 10563
rect 579 10499 597 10563
rect 661 10499 678 10563
rect 742 10499 759 10563
rect 823 10499 840 10563
rect 904 10499 921 10563
rect 985 10499 1002 10563
rect 1066 10499 1083 10563
rect 1147 10499 1164 10563
rect 1228 10499 1245 10563
rect 1309 10499 1326 10563
rect 1390 10499 1407 10563
rect 1471 10499 1488 10563
rect 1552 10499 1569 10563
rect 1633 10499 1650 10563
rect 1714 10499 1731 10563
rect 1795 10499 1812 10563
rect 1876 10499 1893 10563
rect 1957 10499 1974 10563
rect 2038 10499 2055 10563
rect 2119 10499 2136 10563
rect 2200 10499 2217 10563
rect 2281 10499 2298 10563
rect 2362 10499 2379 10563
rect 2443 10499 2460 10563
rect 2524 10499 2541 10563
rect 2605 10499 2622 10563
rect 2686 10499 2703 10563
rect 2767 10499 2784 10563
rect 2848 10499 2865 10563
rect 2929 10499 2946 10563
rect 3010 10499 3027 10563
rect 3091 10499 3108 10563
rect 3172 10499 3189 10563
rect 3253 10499 3270 10563
rect 3334 10499 3351 10563
rect 3415 10499 3432 10563
rect 3496 10499 3513 10563
rect 3577 10499 3594 10563
rect 3658 10499 3675 10563
rect 3739 10499 3756 10563
rect 3820 10499 3837 10563
rect 3901 10499 3918 10563
rect 3982 10499 3999 10563
rect 4063 10499 4080 10563
rect 4144 10499 4161 10563
rect 4225 10499 4242 10563
rect 4306 10499 4323 10563
rect 4387 10499 4404 10563
rect 4468 10499 4485 10563
rect 4549 10499 4566 10563
rect 4630 10499 4647 10563
rect 4711 10499 4728 10563
rect 4792 10499 4809 10563
rect 4873 10499 4879 10563
rect 99 10479 4879 10499
rect 99 10415 105 10479
rect 169 10415 187 10479
rect 251 10415 269 10479
rect 333 10415 351 10479
rect 415 10415 433 10479
rect 497 10415 515 10479
rect 579 10415 597 10479
rect 661 10415 678 10479
rect 742 10415 759 10479
rect 823 10415 840 10479
rect 904 10415 921 10479
rect 985 10415 1002 10479
rect 1066 10415 1083 10479
rect 1147 10415 1164 10479
rect 1228 10415 1245 10479
rect 1309 10415 1326 10479
rect 1390 10415 1407 10479
rect 1471 10415 1488 10479
rect 1552 10415 1569 10479
rect 1633 10415 1650 10479
rect 1714 10415 1731 10479
rect 1795 10415 1812 10479
rect 1876 10415 1893 10479
rect 1957 10415 1974 10479
rect 2038 10415 2055 10479
rect 2119 10415 2136 10479
rect 2200 10415 2217 10479
rect 2281 10415 2298 10479
rect 2362 10415 2379 10479
rect 2443 10415 2460 10479
rect 2524 10415 2541 10479
rect 2605 10415 2622 10479
rect 2686 10415 2703 10479
rect 2767 10415 2784 10479
rect 2848 10415 2865 10479
rect 2929 10415 2946 10479
rect 3010 10415 3027 10479
rect 3091 10415 3108 10479
rect 3172 10415 3189 10479
rect 3253 10415 3270 10479
rect 3334 10415 3351 10479
rect 3415 10415 3432 10479
rect 3496 10415 3513 10479
rect 3577 10415 3594 10479
rect 3658 10415 3675 10479
rect 3739 10415 3756 10479
rect 3820 10415 3837 10479
rect 3901 10415 3918 10479
rect 3982 10415 3999 10479
rect 4063 10415 4080 10479
rect 4144 10415 4161 10479
rect 4225 10415 4242 10479
rect 4306 10415 4323 10479
rect 4387 10415 4404 10479
rect 4468 10415 4485 10479
rect 4549 10415 4566 10479
rect 4630 10415 4647 10479
rect 4711 10415 4728 10479
rect 4792 10415 4809 10479
rect 4873 10415 4879 10479
rect 99 10395 4879 10415
rect 99 10331 105 10395
rect 169 10331 187 10395
rect 251 10331 269 10395
rect 333 10331 351 10395
rect 415 10331 433 10395
rect 497 10331 515 10395
rect 579 10331 597 10395
rect 661 10331 678 10395
rect 742 10331 759 10395
rect 823 10331 840 10395
rect 904 10331 921 10395
rect 985 10331 1002 10395
rect 1066 10331 1083 10395
rect 1147 10331 1164 10395
rect 1228 10331 1245 10395
rect 1309 10331 1326 10395
rect 1390 10331 1407 10395
rect 1471 10331 1488 10395
rect 1552 10331 1569 10395
rect 1633 10331 1650 10395
rect 1714 10331 1731 10395
rect 1795 10331 1812 10395
rect 1876 10331 1893 10395
rect 1957 10331 1974 10395
rect 2038 10331 2055 10395
rect 2119 10331 2136 10395
rect 2200 10331 2217 10395
rect 2281 10331 2298 10395
rect 2362 10331 2379 10395
rect 2443 10331 2460 10395
rect 2524 10331 2541 10395
rect 2605 10331 2622 10395
rect 2686 10331 2703 10395
rect 2767 10331 2784 10395
rect 2848 10331 2865 10395
rect 2929 10331 2946 10395
rect 3010 10331 3027 10395
rect 3091 10331 3108 10395
rect 3172 10331 3189 10395
rect 3253 10331 3270 10395
rect 3334 10331 3351 10395
rect 3415 10331 3432 10395
rect 3496 10331 3513 10395
rect 3577 10331 3594 10395
rect 3658 10331 3675 10395
rect 3739 10331 3756 10395
rect 3820 10331 3837 10395
rect 3901 10331 3918 10395
rect 3982 10331 3999 10395
rect 4063 10331 4080 10395
rect 4144 10331 4161 10395
rect 4225 10331 4242 10395
rect 4306 10331 4323 10395
rect 4387 10331 4404 10395
rect 4468 10331 4485 10395
rect 4549 10331 4566 10395
rect 4630 10331 4647 10395
rect 4711 10331 4728 10395
rect 4792 10331 4809 10395
rect 4873 10331 4879 10395
rect 99 10330 4879 10331
rect 10078 10563 14858 10564
rect 10078 10499 10084 10563
rect 10148 10499 10166 10563
rect 10230 10499 10248 10563
rect 10312 10499 10330 10563
rect 10394 10499 10412 10563
rect 10476 10499 10494 10563
rect 10558 10499 10576 10563
rect 10640 10499 10657 10563
rect 10721 10499 10738 10563
rect 10802 10499 10819 10563
rect 10883 10499 10900 10563
rect 10964 10499 10981 10563
rect 11045 10499 11062 10563
rect 11126 10499 11143 10563
rect 11207 10499 11224 10563
rect 11288 10499 11305 10563
rect 11369 10499 11386 10563
rect 11450 10499 11467 10563
rect 11531 10499 11548 10563
rect 11612 10499 11629 10563
rect 11693 10499 11710 10563
rect 11774 10499 11791 10563
rect 11855 10499 11872 10563
rect 11936 10499 11953 10563
rect 12017 10499 12034 10563
rect 12098 10499 12115 10563
rect 12179 10499 12196 10563
rect 12260 10499 12277 10563
rect 12341 10499 12358 10563
rect 12422 10499 12439 10563
rect 12503 10499 12520 10563
rect 12584 10499 12601 10563
rect 12665 10499 12682 10563
rect 12746 10499 12763 10563
rect 12827 10499 12844 10563
rect 12908 10499 12925 10563
rect 12989 10499 13006 10563
rect 13070 10499 13087 10563
rect 13151 10499 13168 10563
rect 13232 10499 13249 10563
rect 13313 10499 13330 10563
rect 13394 10499 13411 10563
rect 13475 10499 13492 10563
rect 13556 10499 13573 10563
rect 13637 10499 13654 10563
rect 13718 10499 13735 10563
rect 13799 10499 13816 10563
rect 13880 10499 13897 10563
rect 13961 10499 13978 10563
rect 14042 10499 14059 10563
rect 14123 10499 14140 10563
rect 14204 10499 14221 10563
rect 14285 10499 14302 10563
rect 14366 10499 14383 10563
rect 14447 10499 14464 10563
rect 14528 10499 14545 10563
rect 14609 10499 14626 10563
rect 14690 10499 14707 10563
rect 14771 10499 14788 10563
rect 14852 10499 14858 10563
rect 10078 10479 14858 10499
rect 10078 10415 10084 10479
rect 10148 10415 10166 10479
rect 10230 10415 10248 10479
rect 10312 10415 10330 10479
rect 10394 10415 10412 10479
rect 10476 10415 10494 10479
rect 10558 10415 10576 10479
rect 10640 10415 10657 10479
rect 10721 10415 10738 10479
rect 10802 10415 10819 10479
rect 10883 10415 10900 10479
rect 10964 10415 10981 10479
rect 11045 10415 11062 10479
rect 11126 10415 11143 10479
rect 11207 10415 11224 10479
rect 11288 10415 11305 10479
rect 11369 10415 11386 10479
rect 11450 10415 11467 10479
rect 11531 10415 11548 10479
rect 11612 10415 11629 10479
rect 11693 10415 11710 10479
rect 11774 10415 11791 10479
rect 11855 10415 11872 10479
rect 11936 10415 11953 10479
rect 12017 10415 12034 10479
rect 12098 10415 12115 10479
rect 12179 10415 12196 10479
rect 12260 10415 12277 10479
rect 12341 10415 12358 10479
rect 12422 10415 12439 10479
rect 12503 10415 12520 10479
rect 12584 10415 12601 10479
rect 12665 10415 12682 10479
rect 12746 10415 12763 10479
rect 12827 10415 12844 10479
rect 12908 10415 12925 10479
rect 12989 10415 13006 10479
rect 13070 10415 13087 10479
rect 13151 10415 13168 10479
rect 13232 10415 13249 10479
rect 13313 10415 13330 10479
rect 13394 10415 13411 10479
rect 13475 10415 13492 10479
rect 13556 10415 13573 10479
rect 13637 10415 13654 10479
rect 13718 10415 13735 10479
rect 13799 10415 13816 10479
rect 13880 10415 13897 10479
rect 13961 10415 13978 10479
rect 14042 10415 14059 10479
rect 14123 10415 14140 10479
rect 14204 10415 14221 10479
rect 14285 10415 14302 10479
rect 14366 10415 14383 10479
rect 14447 10415 14464 10479
rect 14528 10415 14545 10479
rect 14609 10415 14626 10479
rect 14690 10415 14707 10479
rect 14771 10415 14788 10479
rect 14852 10415 14858 10479
rect 10078 10395 14858 10415
rect 10078 10331 10084 10395
rect 10148 10331 10166 10395
rect 10230 10331 10248 10395
rect 10312 10331 10330 10395
rect 10394 10331 10412 10395
rect 10476 10331 10494 10395
rect 10558 10331 10576 10395
rect 10640 10331 10657 10395
rect 10721 10331 10738 10395
rect 10802 10331 10819 10395
rect 10883 10331 10900 10395
rect 10964 10331 10981 10395
rect 11045 10331 11062 10395
rect 11126 10331 11143 10395
rect 11207 10331 11224 10395
rect 11288 10331 11305 10395
rect 11369 10331 11386 10395
rect 11450 10331 11467 10395
rect 11531 10331 11548 10395
rect 11612 10331 11629 10395
rect 11693 10331 11710 10395
rect 11774 10331 11791 10395
rect 11855 10331 11872 10395
rect 11936 10331 11953 10395
rect 12017 10331 12034 10395
rect 12098 10331 12115 10395
rect 12179 10331 12196 10395
rect 12260 10331 12277 10395
rect 12341 10331 12358 10395
rect 12422 10331 12439 10395
rect 12503 10331 12520 10395
rect 12584 10331 12601 10395
rect 12665 10331 12682 10395
rect 12746 10331 12763 10395
rect 12827 10331 12844 10395
rect 12908 10331 12925 10395
rect 12989 10331 13006 10395
rect 13070 10331 13087 10395
rect 13151 10331 13168 10395
rect 13232 10331 13249 10395
rect 13313 10331 13330 10395
rect 13394 10331 13411 10395
rect 13475 10331 13492 10395
rect 13556 10331 13573 10395
rect 13637 10331 13654 10395
rect 13718 10331 13735 10395
rect 13799 10331 13816 10395
rect 13880 10331 13897 10395
rect 13961 10331 13978 10395
rect 14042 10331 14059 10395
rect 14123 10331 14140 10395
rect 14204 10331 14221 10395
rect 14285 10331 14302 10395
rect 14366 10331 14383 10395
rect 14447 10331 14464 10395
rect 14528 10331 14545 10395
rect 14609 10331 14626 10395
rect 14690 10331 14707 10395
rect 14771 10331 14788 10395
rect 14852 10331 14858 10395
rect 10078 10330 14858 10331
rect 106 9548 112 9612
rect 176 9548 193 9612
rect 257 9548 274 9612
rect 338 9548 355 9612
rect 419 9548 436 9612
rect 500 9548 517 9612
rect 581 9548 598 9612
rect 662 9548 679 9612
rect 743 9548 760 9612
rect 824 9548 841 9612
rect 905 9548 922 9612
rect 986 9548 1003 9612
rect 1067 9548 1084 9612
rect 1148 9548 1165 9612
rect 1229 9548 1246 9612
rect 1310 9548 1327 9612
rect 1391 9548 1408 9612
rect 1472 9548 1489 9612
rect 1553 9548 1570 9612
rect 1634 9548 1651 9612
rect 1715 9548 1732 9612
rect 1796 9548 1813 9612
rect 1877 9548 1894 9612
rect 1958 9548 1975 9612
rect 2039 9548 2056 9612
rect 2120 9548 2137 9612
rect 2201 9548 2218 9612
rect 2282 9548 2299 9612
rect 2363 9548 2380 9612
rect 2444 9548 2461 9612
rect 2525 9548 2542 9612
rect 2606 9548 2623 9612
rect 2687 9548 2704 9612
rect 2768 9548 2785 9612
rect 2849 9548 2866 9612
rect 2930 9548 2947 9612
rect 3011 9548 3028 9612
rect 3092 9548 3109 9612
rect 3173 9548 3190 9612
rect 3254 9548 3271 9612
rect 3335 9548 3352 9612
rect 3416 9548 3433 9612
rect 3497 9548 3514 9612
rect 3578 9548 3595 9612
rect 3659 9548 3676 9612
rect 3740 9548 3757 9612
rect 3821 9548 3838 9612
rect 3902 9548 3919 9612
rect 3983 9548 4000 9612
rect 4064 9548 4081 9612
rect 4145 9548 4162 9612
rect 4226 9548 4243 9612
rect 4307 9548 4324 9612
rect 4388 9548 4405 9612
rect 4469 9548 4486 9612
rect 4550 9548 4567 9612
rect 4631 9548 4648 9612
rect 4712 9548 4729 9612
rect 4793 9548 4809 9612
rect 4873 9548 4879 9612
rect 10078 9548 10084 9612
rect 10148 9548 10165 9612
rect 10229 9548 10246 9612
rect 10310 9548 10327 9612
rect 10391 9548 10408 9612
rect 10472 9548 10489 9612
rect 10553 9548 10570 9612
rect 10634 9548 10651 9612
rect 10715 9548 10732 9612
rect 10796 9548 10813 9612
rect 10877 9548 10894 9612
rect 10958 9548 10975 9612
rect 11039 9548 11056 9612
rect 11120 9548 11137 9612
rect 11201 9548 11218 9612
rect 11282 9548 11299 9612
rect 11363 9548 11380 9612
rect 11444 9548 11461 9612
rect 11525 9548 11542 9612
rect 11606 9548 11623 9612
rect 11687 9548 11704 9612
rect 11768 9548 11785 9612
rect 11849 9548 11866 9612
rect 11930 9548 11947 9612
rect 12011 9548 12028 9612
rect 12092 9548 12109 9612
rect 12173 9548 12190 9612
rect 12254 9548 12271 9612
rect 12335 9548 12352 9612
rect 12416 9548 12433 9612
rect 12497 9548 12514 9612
rect 12578 9548 12595 9612
rect 12659 9548 12676 9612
rect 12740 9548 12757 9612
rect 12821 9548 12838 9612
rect 12902 9548 12919 9612
rect 12983 9548 13000 9612
rect 13064 9548 13081 9612
rect 13145 9548 13162 9612
rect 13226 9548 13243 9612
rect 13307 9548 13324 9612
rect 13388 9548 13405 9612
rect 13469 9548 13486 9612
rect 13550 9548 13567 9612
rect 13631 9548 13648 9612
rect 13712 9548 13729 9612
rect 13793 9548 13810 9612
rect 13874 9548 13891 9612
rect 13955 9548 13972 9612
rect 14036 9548 14053 9612
rect 14117 9548 14134 9612
rect 14198 9548 14215 9612
rect 14279 9548 14296 9612
rect 14360 9548 14378 9612
rect 14442 9548 14460 9612
rect 14524 9548 14542 9612
rect 14606 9548 14624 9612
rect 14688 9548 14706 9612
rect 14770 9548 14788 9612
rect 14852 9548 14858 9612
rect 194 8032 4879 8036
rect 194 7968 200 8032
rect 264 7968 281 8032
rect 345 7968 362 8032
rect 426 7968 443 8032
rect 507 7968 524 8032
rect 588 7968 605 8032
rect 669 7968 686 8032
rect 750 7968 767 8032
rect 831 7968 848 8032
rect 912 7968 929 8032
rect 993 7968 1010 8032
rect 1074 7968 1091 8032
rect 1155 7968 1172 8032
rect 1236 7968 1253 8032
rect 1317 7968 1334 8032
rect 1398 7968 1415 8032
rect 1479 7968 1496 8032
rect 1560 7968 1577 8032
rect 1641 7968 1658 8032
rect 1722 7968 1739 8032
rect 1803 7968 1820 8032
rect 1884 7968 1901 8032
rect 1965 7968 1982 8032
rect 2046 7968 2063 8032
rect 2127 7968 2144 8032
rect 2208 7968 2225 8032
rect 2289 7968 2306 8032
rect 2370 7968 2387 8032
rect 2451 7968 2468 8032
rect 2532 7968 2549 8032
rect 2613 7968 2630 8032
rect 2694 7968 2711 8032
rect 2775 7968 2792 8032
rect 2856 7968 2873 8032
rect 2937 7968 2954 8032
rect 3018 7968 3035 8032
rect 3099 7968 3116 8032
rect 3180 7968 3197 8032
rect 3261 7968 3278 8032
rect 3342 7968 3359 8032
rect 3423 7968 3440 8032
rect 3504 7968 3521 8032
rect 3585 7968 3602 8032
rect 3666 7968 3683 8032
rect 3747 7968 3764 8032
rect 3828 7968 3845 8032
rect 3909 7968 3926 8032
rect 3990 7968 4007 8032
rect 4071 7968 4088 8032
rect 4152 7968 4169 8032
rect 4233 7968 4249 8032
rect 4313 7968 4329 8032
rect 4393 7968 4409 8032
rect 4473 7968 4489 8032
rect 4553 7968 4569 8032
rect 4633 7968 4649 8032
rect 4713 7968 4729 8032
rect 4793 7968 4809 8032
rect 4873 7968 4879 8032
rect 194 7944 4879 7968
rect 194 7880 200 7944
rect 264 7880 281 7944
rect 345 7880 362 7944
rect 426 7880 443 7944
rect 507 7880 524 7944
rect 588 7880 605 7944
rect 669 7880 686 7944
rect 750 7880 767 7944
rect 831 7880 848 7944
rect 912 7880 929 7944
rect 993 7880 1010 7944
rect 1074 7880 1091 7944
rect 1155 7880 1172 7944
rect 1236 7880 1253 7944
rect 1317 7880 1334 7944
rect 1398 7880 1415 7944
rect 1479 7880 1496 7944
rect 1560 7880 1577 7944
rect 1641 7880 1658 7944
rect 1722 7880 1739 7944
rect 1803 7880 1820 7944
rect 1884 7880 1901 7944
rect 1965 7880 1982 7944
rect 2046 7880 2063 7944
rect 2127 7880 2144 7944
rect 2208 7880 2225 7944
rect 2289 7880 2306 7944
rect 2370 7880 2387 7944
rect 2451 7880 2468 7944
rect 2532 7880 2549 7944
rect 2613 7880 2630 7944
rect 2694 7880 2711 7944
rect 2775 7880 2792 7944
rect 2856 7880 2873 7944
rect 2937 7880 2954 7944
rect 3018 7880 3035 7944
rect 3099 7880 3116 7944
rect 3180 7880 3197 7944
rect 3261 7880 3278 7944
rect 3342 7880 3359 7944
rect 3423 7880 3440 7944
rect 3504 7880 3521 7944
rect 3585 7880 3602 7944
rect 3666 7880 3683 7944
rect 3747 7880 3764 7944
rect 3828 7880 3845 7944
rect 3909 7880 3926 7944
rect 3990 7880 4007 7944
rect 4071 7880 4088 7944
rect 4152 7880 4169 7944
rect 4233 7880 4249 7944
rect 4313 7880 4329 7944
rect 4393 7880 4409 7944
rect 4473 7880 4489 7944
rect 4553 7880 4569 7944
rect 4633 7880 4649 7944
rect 4713 7880 4729 7944
rect 4793 7880 4809 7944
rect 4873 7880 4879 7944
rect 194 7856 4879 7880
rect 194 7792 200 7856
rect 264 7792 281 7856
rect 345 7792 362 7856
rect 426 7792 443 7856
rect 507 7792 524 7856
rect 588 7792 605 7856
rect 669 7792 686 7856
rect 750 7792 767 7856
rect 831 7792 848 7856
rect 912 7792 929 7856
rect 993 7792 1010 7856
rect 1074 7792 1091 7856
rect 1155 7792 1172 7856
rect 1236 7792 1253 7856
rect 1317 7792 1334 7856
rect 1398 7792 1415 7856
rect 1479 7792 1496 7856
rect 1560 7792 1577 7856
rect 1641 7792 1658 7856
rect 1722 7792 1739 7856
rect 1803 7792 1820 7856
rect 1884 7792 1901 7856
rect 1965 7792 1982 7856
rect 2046 7792 2063 7856
rect 2127 7792 2144 7856
rect 2208 7792 2225 7856
rect 2289 7792 2306 7856
rect 2370 7792 2387 7856
rect 2451 7792 2468 7856
rect 2532 7792 2549 7856
rect 2613 7792 2630 7856
rect 2694 7792 2711 7856
rect 2775 7792 2792 7856
rect 2856 7792 2873 7856
rect 2937 7792 2954 7856
rect 3018 7792 3035 7856
rect 3099 7792 3116 7856
rect 3180 7792 3197 7856
rect 3261 7792 3278 7856
rect 3342 7792 3359 7856
rect 3423 7792 3440 7856
rect 3504 7792 3521 7856
rect 3585 7792 3602 7856
rect 3666 7792 3683 7856
rect 3747 7792 3764 7856
rect 3828 7792 3845 7856
rect 3909 7792 3926 7856
rect 3990 7792 4007 7856
rect 4071 7792 4088 7856
rect 4152 7792 4169 7856
rect 4233 7792 4249 7856
rect 4313 7792 4329 7856
rect 4393 7792 4409 7856
rect 4473 7792 4489 7856
rect 4553 7792 4569 7856
rect 4633 7792 4649 7856
rect 4713 7792 4729 7856
rect 4793 7792 4809 7856
rect 4873 7792 4879 7856
rect 194 7768 4879 7792
rect 194 7704 200 7768
rect 264 7704 281 7768
rect 345 7704 362 7768
rect 426 7704 443 7768
rect 507 7704 524 7768
rect 588 7704 605 7768
rect 669 7704 686 7768
rect 750 7704 767 7768
rect 831 7704 848 7768
rect 912 7704 929 7768
rect 993 7704 1010 7768
rect 1074 7704 1091 7768
rect 1155 7704 1172 7768
rect 1236 7704 1253 7768
rect 1317 7704 1334 7768
rect 1398 7704 1415 7768
rect 1479 7704 1496 7768
rect 1560 7704 1577 7768
rect 1641 7704 1658 7768
rect 1722 7704 1739 7768
rect 1803 7704 1820 7768
rect 1884 7704 1901 7768
rect 1965 7704 1982 7768
rect 2046 7704 2063 7768
rect 2127 7704 2144 7768
rect 2208 7704 2225 7768
rect 2289 7704 2306 7768
rect 2370 7704 2387 7768
rect 2451 7704 2468 7768
rect 2532 7704 2549 7768
rect 2613 7704 2630 7768
rect 2694 7704 2711 7768
rect 2775 7704 2792 7768
rect 2856 7704 2873 7768
rect 2937 7704 2954 7768
rect 3018 7704 3035 7768
rect 3099 7704 3116 7768
rect 3180 7704 3197 7768
rect 3261 7704 3278 7768
rect 3342 7704 3359 7768
rect 3423 7704 3440 7768
rect 3504 7704 3521 7768
rect 3585 7704 3602 7768
rect 3666 7704 3683 7768
rect 3747 7704 3764 7768
rect 3828 7704 3845 7768
rect 3909 7704 3926 7768
rect 3990 7704 4007 7768
rect 4071 7704 4088 7768
rect 4152 7704 4169 7768
rect 4233 7704 4249 7768
rect 4313 7704 4329 7768
rect 4393 7704 4409 7768
rect 4473 7704 4489 7768
rect 4553 7704 4569 7768
rect 4633 7704 4649 7768
rect 4713 7704 4729 7768
rect 4793 7704 4809 7768
rect 4873 7704 4879 7768
rect 194 7680 4879 7704
rect 194 7616 200 7680
rect 264 7616 281 7680
rect 345 7616 362 7680
rect 426 7616 443 7680
rect 507 7616 524 7680
rect 588 7616 605 7680
rect 669 7616 686 7680
rect 750 7616 767 7680
rect 831 7616 848 7680
rect 912 7616 929 7680
rect 993 7616 1010 7680
rect 1074 7616 1091 7680
rect 1155 7616 1172 7680
rect 1236 7616 1253 7680
rect 1317 7616 1334 7680
rect 1398 7616 1415 7680
rect 1479 7616 1496 7680
rect 1560 7616 1577 7680
rect 1641 7616 1658 7680
rect 1722 7616 1739 7680
rect 1803 7616 1820 7680
rect 1884 7616 1901 7680
rect 1965 7616 1982 7680
rect 2046 7616 2063 7680
rect 2127 7616 2144 7680
rect 2208 7616 2225 7680
rect 2289 7616 2306 7680
rect 2370 7616 2387 7680
rect 2451 7616 2468 7680
rect 2532 7616 2549 7680
rect 2613 7616 2630 7680
rect 2694 7616 2711 7680
rect 2775 7616 2792 7680
rect 2856 7616 2873 7680
rect 2937 7616 2954 7680
rect 3018 7616 3035 7680
rect 3099 7616 3116 7680
rect 3180 7616 3197 7680
rect 3261 7616 3278 7680
rect 3342 7616 3359 7680
rect 3423 7616 3440 7680
rect 3504 7616 3521 7680
rect 3585 7616 3602 7680
rect 3666 7616 3683 7680
rect 3747 7616 3764 7680
rect 3828 7616 3845 7680
rect 3909 7616 3926 7680
rect 3990 7616 4007 7680
rect 4071 7616 4088 7680
rect 4152 7616 4169 7680
rect 4233 7616 4249 7680
rect 4313 7616 4329 7680
rect 4393 7616 4409 7680
rect 4473 7616 4489 7680
rect 4553 7616 4569 7680
rect 4633 7616 4649 7680
rect 4713 7616 4729 7680
rect 4793 7616 4809 7680
rect 4873 7616 4879 7680
rect 194 7592 4879 7616
rect 194 7528 200 7592
rect 264 7528 281 7592
rect 345 7528 362 7592
rect 426 7528 443 7592
rect 507 7528 524 7592
rect 588 7528 605 7592
rect 669 7528 686 7592
rect 750 7528 767 7592
rect 831 7528 848 7592
rect 912 7528 929 7592
rect 993 7528 1010 7592
rect 1074 7528 1091 7592
rect 1155 7528 1172 7592
rect 1236 7528 1253 7592
rect 1317 7528 1334 7592
rect 1398 7528 1415 7592
rect 1479 7528 1496 7592
rect 1560 7528 1577 7592
rect 1641 7528 1658 7592
rect 1722 7528 1739 7592
rect 1803 7528 1820 7592
rect 1884 7528 1901 7592
rect 1965 7528 1982 7592
rect 2046 7528 2063 7592
rect 2127 7528 2144 7592
rect 2208 7528 2225 7592
rect 2289 7528 2306 7592
rect 2370 7528 2387 7592
rect 2451 7528 2468 7592
rect 2532 7528 2549 7592
rect 2613 7528 2630 7592
rect 2694 7528 2711 7592
rect 2775 7528 2792 7592
rect 2856 7528 2873 7592
rect 2937 7528 2954 7592
rect 3018 7528 3035 7592
rect 3099 7528 3116 7592
rect 3180 7528 3197 7592
rect 3261 7528 3278 7592
rect 3342 7528 3359 7592
rect 3423 7528 3440 7592
rect 3504 7528 3521 7592
rect 3585 7528 3602 7592
rect 3666 7528 3683 7592
rect 3747 7528 3764 7592
rect 3828 7528 3845 7592
rect 3909 7528 3926 7592
rect 3990 7528 4007 7592
rect 4071 7528 4088 7592
rect 4152 7528 4169 7592
rect 4233 7528 4249 7592
rect 4313 7528 4329 7592
rect 4393 7528 4409 7592
rect 4473 7528 4489 7592
rect 4553 7528 4569 7592
rect 4633 7528 4649 7592
rect 4713 7528 4729 7592
rect 4793 7528 4809 7592
rect 4873 7528 4879 7592
rect 194 7504 4879 7528
rect 194 7440 200 7504
rect 264 7440 281 7504
rect 345 7440 362 7504
rect 426 7440 443 7504
rect 507 7440 524 7504
rect 588 7440 605 7504
rect 669 7440 686 7504
rect 750 7440 767 7504
rect 831 7440 848 7504
rect 912 7440 929 7504
rect 993 7440 1010 7504
rect 1074 7440 1091 7504
rect 1155 7440 1172 7504
rect 1236 7440 1253 7504
rect 1317 7440 1334 7504
rect 1398 7440 1415 7504
rect 1479 7440 1496 7504
rect 1560 7440 1577 7504
rect 1641 7440 1658 7504
rect 1722 7440 1739 7504
rect 1803 7440 1820 7504
rect 1884 7440 1901 7504
rect 1965 7440 1982 7504
rect 2046 7440 2063 7504
rect 2127 7440 2144 7504
rect 2208 7440 2225 7504
rect 2289 7440 2306 7504
rect 2370 7440 2387 7504
rect 2451 7440 2468 7504
rect 2532 7440 2549 7504
rect 2613 7440 2630 7504
rect 2694 7440 2711 7504
rect 2775 7440 2792 7504
rect 2856 7440 2873 7504
rect 2937 7440 2954 7504
rect 3018 7440 3035 7504
rect 3099 7440 3116 7504
rect 3180 7440 3197 7504
rect 3261 7440 3278 7504
rect 3342 7440 3359 7504
rect 3423 7440 3440 7504
rect 3504 7440 3521 7504
rect 3585 7440 3602 7504
rect 3666 7440 3683 7504
rect 3747 7440 3764 7504
rect 3828 7440 3845 7504
rect 3909 7440 3926 7504
rect 3990 7440 4007 7504
rect 4071 7440 4088 7504
rect 4152 7440 4169 7504
rect 4233 7440 4249 7504
rect 4313 7440 4329 7504
rect 4393 7440 4409 7504
rect 4473 7440 4489 7504
rect 4553 7440 4569 7504
rect 4633 7440 4649 7504
rect 4713 7440 4729 7504
rect 4793 7440 4809 7504
rect 4873 7440 4879 7504
rect 194 7416 4879 7440
rect 194 7352 200 7416
rect 264 7352 281 7416
rect 345 7352 362 7416
rect 426 7352 443 7416
rect 507 7352 524 7416
rect 588 7352 605 7416
rect 669 7352 686 7416
rect 750 7352 767 7416
rect 831 7352 848 7416
rect 912 7352 929 7416
rect 993 7352 1010 7416
rect 1074 7352 1091 7416
rect 1155 7352 1172 7416
rect 1236 7352 1253 7416
rect 1317 7352 1334 7416
rect 1398 7352 1415 7416
rect 1479 7352 1496 7416
rect 1560 7352 1577 7416
rect 1641 7352 1658 7416
rect 1722 7352 1739 7416
rect 1803 7352 1820 7416
rect 1884 7352 1901 7416
rect 1965 7352 1982 7416
rect 2046 7352 2063 7416
rect 2127 7352 2144 7416
rect 2208 7352 2225 7416
rect 2289 7352 2306 7416
rect 2370 7352 2387 7416
rect 2451 7352 2468 7416
rect 2532 7352 2549 7416
rect 2613 7352 2630 7416
rect 2694 7352 2711 7416
rect 2775 7352 2792 7416
rect 2856 7352 2873 7416
rect 2937 7352 2954 7416
rect 3018 7352 3035 7416
rect 3099 7352 3116 7416
rect 3180 7352 3197 7416
rect 3261 7352 3278 7416
rect 3342 7352 3359 7416
rect 3423 7352 3440 7416
rect 3504 7352 3521 7416
rect 3585 7352 3602 7416
rect 3666 7352 3683 7416
rect 3747 7352 3764 7416
rect 3828 7352 3845 7416
rect 3909 7352 3926 7416
rect 3990 7352 4007 7416
rect 4071 7352 4088 7416
rect 4152 7352 4169 7416
rect 4233 7352 4249 7416
rect 4313 7352 4329 7416
rect 4393 7352 4409 7416
rect 4473 7352 4489 7416
rect 4553 7352 4569 7416
rect 4633 7352 4649 7416
rect 4713 7352 4729 7416
rect 4793 7352 4809 7416
rect 4873 7352 4879 7416
rect 194 7348 4879 7352
rect 10078 8032 14858 8036
rect 10078 7968 10084 8032
rect 10148 7968 10166 8032
rect 10230 7968 10248 8032
rect 10312 7968 10330 8032
rect 10394 7968 10412 8032
rect 10476 7968 10494 8032
rect 10558 7968 10576 8032
rect 10640 7968 10657 8032
rect 10721 7968 10738 8032
rect 10802 7968 10819 8032
rect 10883 7968 10900 8032
rect 10964 7968 10981 8032
rect 11045 7968 11062 8032
rect 11126 7968 11143 8032
rect 11207 7968 11224 8032
rect 11288 7968 11305 8032
rect 11369 7968 11386 8032
rect 11450 7968 11467 8032
rect 11531 7968 11548 8032
rect 11612 7968 11629 8032
rect 11693 7968 11710 8032
rect 11774 7968 11791 8032
rect 11855 7968 11872 8032
rect 11936 7968 11953 8032
rect 12017 7968 12034 8032
rect 12098 7968 12115 8032
rect 12179 7968 12196 8032
rect 12260 7968 12277 8032
rect 12341 7968 12358 8032
rect 12422 7968 12439 8032
rect 12503 7968 12520 8032
rect 12584 7968 12601 8032
rect 12665 7968 12682 8032
rect 12746 7968 12763 8032
rect 12827 7968 12844 8032
rect 12908 7968 12925 8032
rect 12989 7968 13006 8032
rect 13070 7968 13087 8032
rect 13151 7968 13168 8032
rect 13232 7968 13249 8032
rect 13313 7968 13330 8032
rect 13394 7968 13411 8032
rect 13475 7968 13492 8032
rect 13556 7968 13573 8032
rect 13637 7968 13654 8032
rect 13718 7968 13735 8032
rect 13799 7968 13816 8032
rect 13880 7968 13897 8032
rect 13961 7968 13978 8032
rect 14042 7968 14059 8032
rect 14123 7968 14140 8032
rect 14204 7968 14221 8032
rect 14285 7968 14302 8032
rect 14366 7968 14383 8032
rect 14447 7968 14464 8032
rect 14528 7968 14545 8032
rect 14609 7968 14626 8032
rect 14690 7968 14707 8032
rect 14771 7968 14788 8032
rect 14852 7968 14858 8032
rect 10078 7944 14858 7968
rect 10078 7880 10084 7944
rect 10148 7880 10166 7944
rect 10230 7880 10248 7944
rect 10312 7880 10330 7944
rect 10394 7880 10412 7944
rect 10476 7880 10494 7944
rect 10558 7880 10576 7944
rect 10640 7880 10657 7944
rect 10721 7880 10738 7944
rect 10802 7880 10819 7944
rect 10883 7880 10900 7944
rect 10964 7880 10981 7944
rect 11045 7880 11062 7944
rect 11126 7880 11143 7944
rect 11207 7880 11224 7944
rect 11288 7880 11305 7944
rect 11369 7880 11386 7944
rect 11450 7880 11467 7944
rect 11531 7880 11548 7944
rect 11612 7880 11629 7944
rect 11693 7880 11710 7944
rect 11774 7880 11791 7944
rect 11855 7880 11872 7944
rect 11936 7880 11953 7944
rect 12017 7880 12034 7944
rect 12098 7880 12115 7944
rect 12179 7880 12196 7944
rect 12260 7880 12277 7944
rect 12341 7880 12358 7944
rect 12422 7880 12439 7944
rect 12503 7880 12520 7944
rect 12584 7880 12601 7944
rect 12665 7880 12682 7944
rect 12746 7880 12763 7944
rect 12827 7880 12844 7944
rect 12908 7880 12925 7944
rect 12989 7880 13006 7944
rect 13070 7880 13087 7944
rect 13151 7880 13168 7944
rect 13232 7880 13249 7944
rect 13313 7880 13330 7944
rect 13394 7880 13411 7944
rect 13475 7880 13492 7944
rect 13556 7880 13573 7944
rect 13637 7880 13654 7944
rect 13718 7880 13735 7944
rect 13799 7880 13816 7944
rect 13880 7880 13897 7944
rect 13961 7880 13978 7944
rect 14042 7880 14059 7944
rect 14123 7880 14140 7944
rect 14204 7880 14221 7944
rect 14285 7880 14302 7944
rect 14366 7880 14383 7944
rect 14447 7880 14464 7944
rect 14528 7880 14545 7944
rect 14609 7880 14626 7944
rect 14690 7880 14707 7944
rect 14771 7880 14788 7944
rect 14852 7880 14858 7944
rect 10078 7856 14858 7880
rect 10078 7792 10084 7856
rect 10148 7792 10166 7856
rect 10230 7792 10248 7856
rect 10312 7792 10330 7856
rect 10394 7792 10412 7856
rect 10476 7792 10494 7856
rect 10558 7792 10576 7856
rect 10640 7792 10657 7856
rect 10721 7792 10738 7856
rect 10802 7792 10819 7856
rect 10883 7792 10900 7856
rect 10964 7792 10981 7856
rect 11045 7792 11062 7856
rect 11126 7792 11143 7856
rect 11207 7792 11224 7856
rect 11288 7792 11305 7856
rect 11369 7792 11386 7856
rect 11450 7792 11467 7856
rect 11531 7792 11548 7856
rect 11612 7792 11629 7856
rect 11693 7792 11710 7856
rect 11774 7792 11791 7856
rect 11855 7792 11872 7856
rect 11936 7792 11953 7856
rect 12017 7792 12034 7856
rect 12098 7792 12115 7856
rect 12179 7792 12196 7856
rect 12260 7792 12277 7856
rect 12341 7792 12358 7856
rect 12422 7792 12439 7856
rect 12503 7792 12520 7856
rect 12584 7792 12601 7856
rect 12665 7792 12682 7856
rect 12746 7792 12763 7856
rect 12827 7792 12844 7856
rect 12908 7792 12925 7856
rect 12989 7792 13006 7856
rect 13070 7792 13087 7856
rect 13151 7792 13168 7856
rect 13232 7792 13249 7856
rect 13313 7792 13330 7856
rect 13394 7792 13411 7856
rect 13475 7792 13492 7856
rect 13556 7792 13573 7856
rect 13637 7792 13654 7856
rect 13718 7792 13735 7856
rect 13799 7792 13816 7856
rect 13880 7792 13897 7856
rect 13961 7792 13978 7856
rect 14042 7792 14059 7856
rect 14123 7792 14140 7856
rect 14204 7792 14221 7856
rect 14285 7792 14302 7856
rect 14366 7792 14383 7856
rect 14447 7792 14464 7856
rect 14528 7792 14545 7856
rect 14609 7792 14626 7856
rect 14690 7792 14707 7856
rect 14771 7792 14788 7856
rect 14852 7792 14858 7856
rect 10078 7768 14858 7792
rect 10078 7704 10084 7768
rect 10148 7704 10166 7768
rect 10230 7704 10248 7768
rect 10312 7704 10330 7768
rect 10394 7704 10412 7768
rect 10476 7704 10494 7768
rect 10558 7704 10576 7768
rect 10640 7704 10657 7768
rect 10721 7704 10738 7768
rect 10802 7704 10819 7768
rect 10883 7704 10900 7768
rect 10964 7704 10981 7768
rect 11045 7704 11062 7768
rect 11126 7704 11143 7768
rect 11207 7704 11224 7768
rect 11288 7704 11305 7768
rect 11369 7704 11386 7768
rect 11450 7704 11467 7768
rect 11531 7704 11548 7768
rect 11612 7704 11629 7768
rect 11693 7704 11710 7768
rect 11774 7704 11791 7768
rect 11855 7704 11872 7768
rect 11936 7704 11953 7768
rect 12017 7704 12034 7768
rect 12098 7704 12115 7768
rect 12179 7704 12196 7768
rect 12260 7704 12277 7768
rect 12341 7704 12358 7768
rect 12422 7704 12439 7768
rect 12503 7704 12520 7768
rect 12584 7704 12601 7768
rect 12665 7704 12682 7768
rect 12746 7704 12763 7768
rect 12827 7704 12844 7768
rect 12908 7704 12925 7768
rect 12989 7704 13006 7768
rect 13070 7704 13087 7768
rect 13151 7704 13168 7768
rect 13232 7704 13249 7768
rect 13313 7704 13330 7768
rect 13394 7704 13411 7768
rect 13475 7704 13492 7768
rect 13556 7704 13573 7768
rect 13637 7704 13654 7768
rect 13718 7704 13735 7768
rect 13799 7704 13816 7768
rect 13880 7704 13897 7768
rect 13961 7704 13978 7768
rect 14042 7704 14059 7768
rect 14123 7704 14140 7768
rect 14204 7704 14221 7768
rect 14285 7704 14302 7768
rect 14366 7704 14383 7768
rect 14447 7704 14464 7768
rect 14528 7704 14545 7768
rect 14609 7704 14626 7768
rect 14690 7704 14707 7768
rect 14771 7704 14788 7768
rect 14852 7704 14858 7768
rect 10078 7680 14858 7704
rect 10078 7616 10084 7680
rect 10148 7616 10166 7680
rect 10230 7616 10248 7680
rect 10312 7616 10330 7680
rect 10394 7616 10412 7680
rect 10476 7616 10494 7680
rect 10558 7616 10576 7680
rect 10640 7616 10657 7680
rect 10721 7616 10738 7680
rect 10802 7616 10819 7680
rect 10883 7616 10900 7680
rect 10964 7616 10981 7680
rect 11045 7616 11062 7680
rect 11126 7616 11143 7680
rect 11207 7616 11224 7680
rect 11288 7616 11305 7680
rect 11369 7616 11386 7680
rect 11450 7616 11467 7680
rect 11531 7616 11548 7680
rect 11612 7616 11629 7680
rect 11693 7616 11710 7680
rect 11774 7616 11791 7680
rect 11855 7616 11872 7680
rect 11936 7616 11953 7680
rect 12017 7616 12034 7680
rect 12098 7616 12115 7680
rect 12179 7616 12196 7680
rect 12260 7616 12277 7680
rect 12341 7616 12358 7680
rect 12422 7616 12439 7680
rect 12503 7616 12520 7680
rect 12584 7616 12601 7680
rect 12665 7616 12682 7680
rect 12746 7616 12763 7680
rect 12827 7616 12844 7680
rect 12908 7616 12925 7680
rect 12989 7616 13006 7680
rect 13070 7616 13087 7680
rect 13151 7616 13168 7680
rect 13232 7616 13249 7680
rect 13313 7616 13330 7680
rect 13394 7616 13411 7680
rect 13475 7616 13492 7680
rect 13556 7616 13573 7680
rect 13637 7616 13654 7680
rect 13718 7616 13735 7680
rect 13799 7616 13816 7680
rect 13880 7616 13897 7680
rect 13961 7616 13978 7680
rect 14042 7616 14059 7680
rect 14123 7616 14140 7680
rect 14204 7616 14221 7680
rect 14285 7616 14302 7680
rect 14366 7616 14383 7680
rect 14447 7616 14464 7680
rect 14528 7616 14545 7680
rect 14609 7616 14626 7680
rect 14690 7616 14707 7680
rect 14771 7616 14788 7680
rect 14852 7616 14858 7680
rect 10078 7592 14858 7616
rect 10078 7528 10084 7592
rect 10148 7528 10166 7592
rect 10230 7528 10248 7592
rect 10312 7528 10330 7592
rect 10394 7528 10412 7592
rect 10476 7528 10494 7592
rect 10558 7528 10576 7592
rect 10640 7528 10657 7592
rect 10721 7528 10738 7592
rect 10802 7528 10819 7592
rect 10883 7528 10900 7592
rect 10964 7528 10981 7592
rect 11045 7528 11062 7592
rect 11126 7528 11143 7592
rect 11207 7528 11224 7592
rect 11288 7528 11305 7592
rect 11369 7528 11386 7592
rect 11450 7528 11467 7592
rect 11531 7528 11548 7592
rect 11612 7528 11629 7592
rect 11693 7528 11710 7592
rect 11774 7528 11791 7592
rect 11855 7528 11872 7592
rect 11936 7528 11953 7592
rect 12017 7528 12034 7592
rect 12098 7528 12115 7592
rect 12179 7528 12196 7592
rect 12260 7528 12277 7592
rect 12341 7528 12358 7592
rect 12422 7528 12439 7592
rect 12503 7528 12520 7592
rect 12584 7528 12601 7592
rect 12665 7528 12682 7592
rect 12746 7528 12763 7592
rect 12827 7528 12844 7592
rect 12908 7528 12925 7592
rect 12989 7528 13006 7592
rect 13070 7528 13087 7592
rect 13151 7528 13168 7592
rect 13232 7528 13249 7592
rect 13313 7528 13330 7592
rect 13394 7528 13411 7592
rect 13475 7528 13492 7592
rect 13556 7528 13573 7592
rect 13637 7528 13654 7592
rect 13718 7528 13735 7592
rect 13799 7528 13816 7592
rect 13880 7528 13897 7592
rect 13961 7528 13978 7592
rect 14042 7528 14059 7592
rect 14123 7528 14140 7592
rect 14204 7528 14221 7592
rect 14285 7528 14302 7592
rect 14366 7528 14383 7592
rect 14447 7528 14464 7592
rect 14528 7528 14545 7592
rect 14609 7528 14626 7592
rect 14690 7528 14707 7592
rect 14771 7528 14788 7592
rect 14852 7528 14858 7592
rect 10078 7504 14858 7528
rect 10078 7440 10084 7504
rect 10148 7440 10166 7504
rect 10230 7440 10248 7504
rect 10312 7440 10330 7504
rect 10394 7440 10412 7504
rect 10476 7440 10494 7504
rect 10558 7440 10576 7504
rect 10640 7440 10657 7504
rect 10721 7440 10738 7504
rect 10802 7440 10819 7504
rect 10883 7440 10900 7504
rect 10964 7440 10981 7504
rect 11045 7440 11062 7504
rect 11126 7440 11143 7504
rect 11207 7440 11224 7504
rect 11288 7440 11305 7504
rect 11369 7440 11386 7504
rect 11450 7440 11467 7504
rect 11531 7440 11548 7504
rect 11612 7440 11629 7504
rect 11693 7440 11710 7504
rect 11774 7440 11791 7504
rect 11855 7440 11872 7504
rect 11936 7440 11953 7504
rect 12017 7440 12034 7504
rect 12098 7440 12115 7504
rect 12179 7440 12196 7504
rect 12260 7440 12277 7504
rect 12341 7440 12358 7504
rect 12422 7440 12439 7504
rect 12503 7440 12520 7504
rect 12584 7440 12601 7504
rect 12665 7440 12682 7504
rect 12746 7440 12763 7504
rect 12827 7440 12844 7504
rect 12908 7440 12925 7504
rect 12989 7440 13006 7504
rect 13070 7440 13087 7504
rect 13151 7440 13168 7504
rect 13232 7440 13249 7504
rect 13313 7440 13330 7504
rect 13394 7440 13411 7504
rect 13475 7440 13492 7504
rect 13556 7440 13573 7504
rect 13637 7440 13654 7504
rect 13718 7440 13735 7504
rect 13799 7440 13816 7504
rect 13880 7440 13897 7504
rect 13961 7440 13978 7504
rect 14042 7440 14059 7504
rect 14123 7440 14140 7504
rect 14204 7440 14221 7504
rect 14285 7440 14302 7504
rect 14366 7440 14383 7504
rect 14447 7440 14464 7504
rect 14528 7440 14545 7504
rect 14609 7440 14626 7504
rect 14690 7440 14707 7504
rect 14771 7440 14788 7504
rect 14852 7440 14858 7504
rect 10078 7416 14858 7440
rect 10078 7352 10084 7416
rect 10148 7352 10166 7416
rect 10230 7352 10248 7416
rect 10312 7352 10330 7416
rect 10394 7352 10412 7416
rect 10476 7352 10494 7416
rect 10558 7352 10576 7416
rect 10640 7352 10657 7416
rect 10721 7352 10738 7416
rect 10802 7352 10819 7416
rect 10883 7352 10900 7416
rect 10964 7352 10981 7416
rect 11045 7352 11062 7416
rect 11126 7352 11143 7416
rect 11207 7352 11224 7416
rect 11288 7352 11305 7416
rect 11369 7352 11386 7416
rect 11450 7352 11467 7416
rect 11531 7352 11548 7416
rect 11612 7352 11629 7416
rect 11693 7352 11710 7416
rect 11774 7352 11791 7416
rect 11855 7352 11872 7416
rect 11936 7352 11953 7416
rect 12017 7352 12034 7416
rect 12098 7352 12115 7416
rect 12179 7352 12196 7416
rect 12260 7352 12277 7416
rect 12341 7352 12358 7416
rect 12422 7352 12439 7416
rect 12503 7352 12520 7416
rect 12584 7352 12601 7416
rect 12665 7352 12682 7416
rect 12746 7352 12763 7416
rect 12827 7352 12844 7416
rect 12908 7352 12925 7416
rect 12989 7352 13006 7416
rect 13070 7352 13087 7416
rect 13151 7352 13168 7416
rect 13232 7352 13249 7416
rect 13313 7352 13330 7416
rect 13394 7352 13411 7416
rect 13475 7352 13492 7416
rect 13556 7352 13573 7416
rect 13637 7352 13654 7416
rect 13718 7352 13735 7416
rect 13799 7352 13816 7416
rect 13880 7352 13897 7416
rect 13961 7352 13978 7416
rect 14042 7352 14059 7416
rect 14123 7352 14140 7416
rect 14204 7352 14221 7416
rect 14285 7352 14302 7416
rect 14366 7352 14383 7416
rect 14447 7352 14464 7416
rect 14528 7352 14545 7416
rect 14609 7352 14626 7416
rect 14690 7352 14707 7416
rect 14771 7352 14788 7416
rect 14852 7352 14858 7416
rect 10078 7348 14858 7352
<< via3 >>
rect 112 11282 176 11346
rect 193 11282 257 11346
rect 274 11282 338 11346
rect 355 11282 419 11346
rect 436 11282 500 11346
rect 517 11282 581 11346
rect 598 11282 662 11346
rect 679 11282 743 11346
rect 760 11282 824 11346
rect 841 11282 905 11346
rect 922 11282 986 11346
rect 1003 11282 1067 11346
rect 1084 11282 1148 11346
rect 1165 11282 1229 11346
rect 1246 11282 1310 11346
rect 1327 11282 1391 11346
rect 1408 11282 1472 11346
rect 1489 11282 1553 11346
rect 1570 11282 1634 11346
rect 1651 11282 1715 11346
rect 1732 11282 1796 11346
rect 1813 11282 1877 11346
rect 1894 11282 1958 11346
rect 1975 11282 2039 11346
rect 2056 11282 2120 11346
rect 2137 11282 2201 11346
rect 2218 11282 2282 11346
rect 2299 11282 2363 11346
rect 2380 11282 2444 11346
rect 2461 11282 2525 11346
rect 2542 11282 2606 11346
rect 2623 11282 2687 11346
rect 2704 11282 2768 11346
rect 2785 11282 2849 11346
rect 2866 11282 2930 11346
rect 2947 11282 3011 11346
rect 3028 11282 3092 11346
rect 3109 11282 3173 11346
rect 3190 11282 3254 11346
rect 3271 11282 3335 11346
rect 3352 11282 3416 11346
rect 3433 11282 3497 11346
rect 3514 11282 3578 11346
rect 3595 11282 3659 11346
rect 3676 11282 3740 11346
rect 3757 11282 3821 11346
rect 3838 11282 3902 11346
rect 3919 11282 3983 11346
rect 4000 11282 4064 11346
rect 4081 11282 4145 11346
rect 4162 11282 4226 11346
rect 4243 11282 4307 11346
rect 4324 11282 4388 11346
rect 4405 11282 4469 11346
rect 4486 11282 4550 11346
rect 4567 11282 4631 11346
rect 4648 11282 4712 11346
rect 4729 11282 4793 11346
rect 4809 11282 4873 11346
rect 10084 11282 10148 11346
rect 10165 11282 10229 11346
rect 10246 11282 10310 11346
rect 10327 11282 10391 11346
rect 10408 11282 10472 11346
rect 10489 11282 10553 11346
rect 10570 11282 10634 11346
rect 10651 11282 10715 11346
rect 10732 11282 10796 11346
rect 10813 11282 10877 11346
rect 10894 11282 10958 11346
rect 10975 11282 11039 11346
rect 11056 11282 11120 11346
rect 11137 11282 11201 11346
rect 11218 11282 11282 11346
rect 11299 11282 11363 11346
rect 11380 11282 11444 11346
rect 11461 11282 11525 11346
rect 11542 11282 11606 11346
rect 11623 11282 11687 11346
rect 11704 11282 11768 11346
rect 11785 11282 11849 11346
rect 11866 11282 11930 11346
rect 11947 11282 12011 11346
rect 12028 11282 12092 11346
rect 12109 11282 12173 11346
rect 12190 11282 12254 11346
rect 12271 11282 12335 11346
rect 12352 11282 12416 11346
rect 12433 11282 12497 11346
rect 12514 11282 12578 11346
rect 12595 11282 12659 11346
rect 12676 11282 12740 11346
rect 12757 11282 12821 11346
rect 12838 11282 12902 11346
rect 12919 11282 12983 11346
rect 13000 11282 13064 11346
rect 13081 11282 13145 11346
rect 13162 11282 13226 11346
rect 13243 11282 13307 11346
rect 13324 11282 13388 11346
rect 13405 11282 13469 11346
rect 13486 11282 13550 11346
rect 13567 11282 13631 11346
rect 13648 11282 13712 11346
rect 13729 11282 13793 11346
rect 13810 11282 13874 11346
rect 13891 11282 13955 11346
rect 13972 11282 14036 11346
rect 14053 11282 14117 11346
rect 14134 11282 14198 11346
rect 14215 11282 14279 11346
rect 14296 11282 14360 11346
rect 14378 11282 14442 11346
rect 14460 11282 14524 11346
rect 14542 11282 14606 11346
rect 14624 11282 14688 11346
rect 14706 11282 14770 11346
rect 14788 11282 14852 11346
rect 105 10499 169 10563
rect 187 10499 251 10563
rect 269 10499 333 10563
rect 351 10499 415 10563
rect 433 10499 497 10563
rect 515 10499 579 10563
rect 597 10499 661 10563
rect 678 10499 742 10563
rect 759 10499 823 10563
rect 840 10499 904 10563
rect 921 10499 985 10563
rect 1002 10499 1066 10563
rect 1083 10499 1147 10563
rect 1164 10499 1228 10563
rect 1245 10499 1309 10563
rect 1326 10499 1390 10563
rect 1407 10499 1471 10563
rect 1488 10499 1552 10563
rect 1569 10499 1633 10563
rect 1650 10499 1714 10563
rect 1731 10499 1795 10563
rect 1812 10499 1876 10563
rect 1893 10499 1957 10563
rect 1974 10499 2038 10563
rect 2055 10499 2119 10563
rect 2136 10499 2200 10563
rect 2217 10499 2281 10563
rect 2298 10499 2362 10563
rect 2379 10499 2443 10563
rect 2460 10499 2524 10563
rect 2541 10499 2605 10563
rect 2622 10499 2686 10563
rect 2703 10499 2767 10563
rect 2784 10499 2848 10563
rect 2865 10499 2929 10563
rect 2946 10499 3010 10563
rect 3027 10499 3091 10563
rect 3108 10499 3172 10563
rect 3189 10499 3253 10563
rect 3270 10499 3334 10563
rect 3351 10499 3415 10563
rect 3432 10499 3496 10563
rect 3513 10499 3577 10563
rect 3594 10499 3658 10563
rect 3675 10499 3739 10563
rect 3756 10499 3820 10563
rect 3837 10499 3901 10563
rect 3918 10499 3982 10563
rect 3999 10499 4063 10563
rect 4080 10499 4144 10563
rect 4161 10499 4225 10563
rect 4242 10499 4306 10563
rect 4323 10499 4387 10563
rect 4404 10499 4468 10563
rect 4485 10499 4549 10563
rect 4566 10499 4630 10563
rect 4647 10499 4711 10563
rect 4728 10499 4792 10563
rect 4809 10499 4873 10563
rect 105 10415 169 10479
rect 187 10415 251 10479
rect 269 10415 333 10479
rect 351 10415 415 10479
rect 433 10415 497 10479
rect 515 10415 579 10479
rect 597 10415 661 10479
rect 678 10415 742 10479
rect 759 10415 823 10479
rect 840 10415 904 10479
rect 921 10415 985 10479
rect 1002 10415 1066 10479
rect 1083 10415 1147 10479
rect 1164 10415 1228 10479
rect 1245 10415 1309 10479
rect 1326 10415 1390 10479
rect 1407 10415 1471 10479
rect 1488 10415 1552 10479
rect 1569 10415 1633 10479
rect 1650 10415 1714 10479
rect 1731 10415 1795 10479
rect 1812 10415 1876 10479
rect 1893 10415 1957 10479
rect 1974 10415 2038 10479
rect 2055 10415 2119 10479
rect 2136 10415 2200 10479
rect 2217 10415 2281 10479
rect 2298 10415 2362 10479
rect 2379 10415 2443 10479
rect 2460 10415 2524 10479
rect 2541 10415 2605 10479
rect 2622 10415 2686 10479
rect 2703 10415 2767 10479
rect 2784 10415 2848 10479
rect 2865 10415 2929 10479
rect 2946 10415 3010 10479
rect 3027 10415 3091 10479
rect 3108 10415 3172 10479
rect 3189 10415 3253 10479
rect 3270 10415 3334 10479
rect 3351 10415 3415 10479
rect 3432 10415 3496 10479
rect 3513 10415 3577 10479
rect 3594 10415 3658 10479
rect 3675 10415 3739 10479
rect 3756 10415 3820 10479
rect 3837 10415 3901 10479
rect 3918 10415 3982 10479
rect 3999 10415 4063 10479
rect 4080 10415 4144 10479
rect 4161 10415 4225 10479
rect 4242 10415 4306 10479
rect 4323 10415 4387 10479
rect 4404 10415 4468 10479
rect 4485 10415 4549 10479
rect 4566 10415 4630 10479
rect 4647 10415 4711 10479
rect 4728 10415 4792 10479
rect 4809 10415 4873 10479
rect 105 10331 169 10395
rect 187 10331 251 10395
rect 269 10331 333 10395
rect 351 10331 415 10395
rect 433 10331 497 10395
rect 515 10331 579 10395
rect 597 10331 661 10395
rect 678 10331 742 10395
rect 759 10331 823 10395
rect 840 10331 904 10395
rect 921 10331 985 10395
rect 1002 10331 1066 10395
rect 1083 10331 1147 10395
rect 1164 10331 1228 10395
rect 1245 10331 1309 10395
rect 1326 10331 1390 10395
rect 1407 10331 1471 10395
rect 1488 10331 1552 10395
rect 1569 10331 1633 10395
rect 1650 10331 1714 10395
rect 1731 10331 1795 10395
rect 1812 10331 1876 10395
rect 1893 10331 1957 10395
rect 1974 10331 2038 10395
rect 2055 10331 2119 10395
rect 2136 10331 2200 10395
rect 2217 10331 2281 10395
rect 2298 10331 2362 10395
rect 2379 10331 2443 10395
rect 2460 10331 2524 10395
rect 2541 10331 2605 10395
rect 2622 10331 2686 10395
rect 2703 10331 2767 10395
rect 2784 10331 2848 10395
rect 2865 10331 2929 10395
rect 2946 10331 3010 10395
rect 3027 10331 3091 10395
rect 3108 10331 3172 10395
rect 3189 10331 3253 10395
rect 3270 10331 3334 10395
rect 3351 10331 3415 10395
rect 3432 10331 3496 10395
rect 3513 10331 3577 10395
rect 3594 10331 3658 10395
rect 3675 10331 3739 10395
rect 3756 10331 3820 10395
rect 3837 10331 3901 10395
rect 3918 10331 3982 10395
rect 3999 10331 4063 10395
rect 4080 10331 4144 10395
rect 4161 10331 4225 10395
rect 4242 10331 4306 10395
rect 4323 10331 4387 10395
rect 4404 10331 4468 10395
rect 4485 10331 4549 10395
rect 4566 10331 4630 10395
rect 4647 10331 4711 10395
rect 4728 10331 4792 10395
rect 4809 10331 4873 10395
rect 10084 10499 10148 10563
rect 10166 10499 10230 10563
rect 10248 10499 10312 10563
rect 10330 10499 10394 10563
rect 10412 10499 10476 10563
rect 10494 10499 10558 10563
rect 10576 10499 10640 10563
rect 10657 10499 10721 10563
rect 10738 10499 10802 10563
rect 10819 10499 10883 10563
rect 10900 10499 10964 10563
rect 10981 10499 11045 10563
rect 11062 10499 11126 10563
rect 11143 10499 11207 10563
rect 11224 10499 11288 10563
rect 11305 10499 11369 10563
rect 11386 10499 11450 10563
rect 11467 10499 11531 10563
rect 11548 10499 11612 10563
rect 11629 10499 11693 10563
rect 11710 10499 11774 10563
rect 11791 10499 11855 10563
rect 11872 10499 11936 10563
rect 11953 10499 12017 10563
rect 12034 10499 12098 10563
rect 12115 10499 12179 10563
rect 12196 10499 12260 10563
rect 12277 10499 12341 10563
rect 12358 10499 12422 10563
rect 12439 10499 12503 10563
rect 12520 10499 12584 10563
rect 12601 10499 12665 10563
rect 12682 10499 12746 10563
rect 12763 10499 12827 10563
rect 12844 10499 12908 10563
rect 12925 10499 12989 10563
rect 13006 10499 13070 10563
rect 13087 10499 13151 10563
rect 13168 10499 13232 10563
rect 13249 10499 13313 10563
rect 13330 10499 13394 10563
rect 13411 10499 13475 10563
rect 13492 10499 13556 10563
rect 13573 10499 13637 10563
rect 13654 10499 13718 10563
rect 13735 10499 13799 10563
rect 13816 10499 13880 10563
rect 13897 10499 13961 10563
rect 13978 10499 14042 10563
rect 14059 10499 14123 10563
rect 14140 10499 14204 10563
rect 14221 10499 14285 10563
rect 14302 10499 14366 10563
rect 14383 10499 14447 10563
rect 14464 10499 14528 10563
rect 14545 10499 14609 10563
rect 14626 10499 14690 10563
rect 14707 10499 14771 10563
rect 14788 10499 14852 10563
rect 10084 10415 10148 10479
rect 10166 10415 10230 10479
rect 10248 10415 10312 10479
rect 10330 10415 10394 10479
rect 10412 10415 10476 10479
rect 10494 10415 10558 10479
rect 10576 10415 10640 10479
rect 10657 10415 10721 10479
rect 10738 10415 10802 10479
rect 10819 10415 10883 10479
rect 10900 10415 10964 10479
rect 10981 10415 11045 10479
rect 11062 10415 11126 10479
rect 11143 10415 11207 10479
rect 11224 10415 11288 10479
rect 11305 10415 11369 10479
rect 11386 10415 11450 10479
rect 11467 10415 11531 10479
rect 11548 10415 11612 10479
rect 11629 10415 11693 10479
rect 11710 10415 11774 10479
rect 11791 10415 11855 10479
rect 11872 10415 11936 10479
rect 11953 10415 12017 10479
rect 12034 10415 12098 10479
rect 12115 10415 12179 10479
rect 12196 10415 12260 10479
rect 12277 10415 12341 10479
rect 12358 10415 12422 10479
rect 12439 10415 12503 10479
rect 12520 10415 12584 10479
rect 12601 10415 12665 10479
rect 12682 10415 12746 10479
rect 12763 10415 12827 10479
rect 12844 10415 12908 10479
rect 12925 10415 12989 10479
rect 13006 10415 13070 10479
rect 13087 10415 13151 10479
rect 13168 10415 13232 10479
rect 13249 10415 13313 10479
rect 13330 10415 13394 10479
rect 13411 10415 13475 10479
rect 13492 10415 13556 10479
rect 13573 10415 13637 10479
rect 13654 10415 13718 10479
rect 13735 10415 13799 10479
rect 13816 10415 13880 10479
rect 13897 10415 13961 10479
rect 13978 10415 14042 10479
rect 14059 10415 14123 10479
rect 14140 10415 14204 10479
rect 14221 10415 14285 10479
rect 14302 10415 14366 10479
rect 14383 10415 14447 10479
rect 14464 10415 14528 10479
rect 14545 10415 14609 10479
rect 14626 10415 14690 10479
rect 14707 10415 14771 10479
rect 14788 10415 14852 10479
rect 10084 10331 10148 10395
rect 10166 10331 10230 10395
rect 10248 10331 10312 10395
rect 10330 10331 10394 10395
rect 10412 10331 10476 10395
rect 10494 10331 10558 10395
rect 10576 10331 10640 10395
rect 10657 10331 10721 10395
rect 10738 10331 10802 10395
rect 10819 10331 10883 10395
rect 10900 10331 10964 10395
rect 10981 10331 11045 10395
rect 11062 10331 11126 10395
rect 11143 10331 11207 10395
rect 11224 10331 11288 10395
rect 11305 10331 11369 10395
rect 11386 10331 11450 10395
rect 11467 10331 11531 10395
rect 11548 10331 11612 10395
rect 11629 10331 11693 10395
rect 11710 10331 11774 10395
rect 11791 10331 11855 10395
rect 11872 10331 11936 10395
rect 11953 10331 12017 10395
rect 12034 10331 12098 10395
rect 12115 10331 12179 10395
rect 12196 10331 12260 10395
rect 12277 10331 12341 10395
rect 12358 10331 12422 10395
rect 12439 10331 12503 10395
rect 12520 10331 12584 10395
rect 12601 10331 12665 10395
rect 12682 10331 12746 10395
rect 12763 10331 12827 10395
rect 12844 10331 12908 10395
rect 12925 10331 12989 10395
rect 13006 10331 13070 10395
rect 13087 10331 13151 10395
rect 13168 10331 13232 10395
rect 13249 10331 13313 10395
rect 13330 10331 13394 10395
rect 13411 10331 13475 10395
rect 13492 10331 13556 10395
rect 13573 10331 13637 10395
rect 13654 10331 13718 10395
rect 13735 10331 13799 10395
rect 13816 10331 13880 10395
rect 13897 10331 13961 10395
rect 13978 10331 14042 10395
rect 14059 10331 14123 10395
rect 14140 10331 14204 10395
rect 14221 10331 14285 10395
rect 14302 10331 14366 10395
rect 14383 10331 14447 10395
rect 14464 10331 14528 10395
rect 14545 10331 14609 10395
rect 14626 10331 14690 10395
rect 14707 10331 14771 10395
rect 14788 10331 14852 10395
rect 112 9548 176 9612
rect 193 9548 257 9612
rect 274 9548 338 9612
rect 355 9548 419 9612
rect 436 9548 500 9612
rect 517 9548 581 9612
rect 598 9548 662 9612
rect 679 9548 743 9612
rect 760 9548 824 9612
rect 841 9548 905 9612
rect 922 9548 986 9612
rect 1003 9548 1067 9612
rect 1084 9548 1148 9612
rect 1165 9548 1229 9612
rect 1246 9548 1310 9612
rect 1327 9548 1391 9612
rect 1408 9548 1472 9612
rect 1489 9548 1553 9612
rect 1570 9548 1634 9612
rect 1651 9548 1715 9612
rect 1732 9548 1796 9612
rect 1813 9548 1877 9612
rect 1894 9548 1958 9612
rect 1975 9548 2039 9612
rect 2056 9548 2120 9612
rect 2137 9548 2201 9612
rect 2218 9548 2282 9612
rect 2299 9548 2363 9612
rect 2380 9548 2444 9612
rect 2461 9548 2525 9612
rect 2542 9548 2606 9612
rect 2623 9548 2687 9612
rect 2704 9548 2768 9612
rect 2785 9548 2849 9612
rect 2866 9548 2930 9612
rect 2947 9548 3011 9612
rect 3028 9548 3092 9612
rect 3109 9548 3173 9612
rect 3190 9548 3254 9612
rect 3271 9548 3335 9612
rect 3352 9548 3416 9612
rect 3433 9548 3497 9612
rect 3514 9548 3578 9612
rect 3595 9548 3659 9612
rect 3676 9548 3740 9612
rect 3757 9548 3821 9612
rect 3838 9548 3902 9612
rect 3919 9548 3983 9612
rect 4000 9548 4064 9612
rect 4081 9548 4145 9612
rect 4162 9548 4226 9612
rect 4243 9548 4307 9612
rect 4324 9548 4388 9612
rect 4405 9548 4469 9612
rect 4486 9548 4550 9612
rect 4567 9548 4631 9612
rect 4648 9548 4712 9612
rect 4729 9548 4793 9612
rect 4809 9548 4873 9612
rect 10084 9548 10148 9612
rect 10165 9548 10229 9612
rect 10246 9548 10310 9612
rect 10327 9548 10391 9612
rect 10408 9548 10472 9612
rect 10489 9548 10553 9612
rect 10570 9548 10634 9612
rect 10651 9548 10715 9612
rect 10732 9548 10796 9612
rect 10813 9548 10877 9612
rect 10894 9548 10958 9612
rect 10975 9548 11039 9612
rect 11056 9548 11120 9612
rect 11137 9548 11201 9612
rect 11218 9548 11282 9612
rect 11299 9548 11363 9612
rect 11380 9548 11444 9612
rect 11461 9548 11525 9612
rect 11542 9548 11606 9612
rect 11623 9548 11687 9612
rect 11704 9548 11768 9612
rect 11785 9548 11849 9612
rect 11866 9548 11930 9612
rect 11947 9548 12011 9612
rect 12028 9548 12092 9612
rect 12109 9548 12173 9612
rect 12190 9548 12254 9612
rect 12271 9548 12335 9612
rect 12352 9548 12416 9612
rect 12433 9548 12497 9612
rect 12514 9548 12578 9612
rect 12595 9548 12659 9612
rect 12676 9548 12740 9612
rect 12757 9548 12821 9612
rect 12838 9548 12902 9612
rect 12919 9548 12983 9612
rect 13000 9548 13064 9612
rect 13081 9548 13145 9612
rect 13162 9548 13226 9612
rect 13243 9548 13307 9612
rect 13324 9548 13388 9612
rect 13405 9548 13469 9612
rect 13486 9548 13550 9612
rect 13567 9548 13631 9612
rect 13648 9548 13712 9612
rect 13729 9548 13793 9612
rect 13810 9548 13874 9612
rect 13891 9548 13955 9612
rect 13972 9548 14036 9612
rect 14053 9548 14117 9612
rect 14134 9548 14198 9612
rect 14215 9548 14279 9612
rect 14296 9548 14360 9612
rect 14378 9548 14442 9612
rect 14460 9548 14524 9612
rect 14542 9548 14606 9612
rect 14624 9548 14688 9612
rect 14706 9548 14770 9612
rect 14788 9548 14852 9612
rect 200 7968 264 8032
rect 281 7968 345 8032
rect 362 7968 426 8032
rect 443 7968 507 8032
rect 524 7968 588 8032
rect 605 7968 669 8032
rect 686 7968 750 8032
rect 767 7968 831 8032
rect 848 7968 912 8032
rect 929 7968 993 8032
rect 1010 7968 1074 8032
rect 1091 7968 1155 8032
rect 1172 7968 1236 8032
rect 1253 7968 1317 8032
rect 1334 7968 1398 8032
rect 1415 7968 1479 8032
rect 1496 7968 1560 8032
rect 1577 7968 1641 8032
rect 1658 7968 1722 8032
rect 1739 7968 1803 8032
rect 1820 7968 1884 8032
rect 1901 7968 1965 8032
rect 1982 7968 2046 8032
rect 2063 7968 2127 8032
rect 2144 7968 2208 8032
rect 2225 7968 2289 8032
rect 2306 7968 2370 8032
rect 2387 7968 2451 8032
rect 2468 7968 2532 8032
rect 2549 7968 2613 8032
rect 2630 7968 2694 8032
rect 2711 7968 2775 8032
rect 2792 7968 2856 8032
rect 2873 7968 2937 8032
rect 2954 7968 3018 8032
rect 3035 7968 3099 8032
rect 3116 7968 3180 8032
rect 3197 7968 3261 8032
rect 3278 7968 3342 8032
rect 3359 7968 3423 8032
rect 3440 7968 3504 8032
rect 3521 7968 3585 8032
rect 3602 7968 3666 8032
rect 3683 7968 3747 8032
rect 3764 7968 3828 8032
rect 3845 7968 3909 8032
rect 3926 7968 3990 8032
rect 4007 7968 4071 8032
rect 4088 7968 4152 8032
rect 4169 7968 4233 8032
rect 4249 7968 4313 8032
rect 4329 7968 4393 8032
rect 4409 7968 4473 8032
rect 4489 7968 4553 8032
rect 4569 7968 4633 8032
rect 4649 7968 4713 8032
rect 4729 7968 4793 8032
rect 4809 7968 4873 8032
rect 200 7880 264 7944
rect 281 7880 345 7944
rect 362 7880 426 7944
rect 443 7880 507 7944
rect 524 7880 588 7944
rect 605 7880 669 7944
rect 686 7880 750 7944
rect 767 7880 831 7944
rect 848 7880 912 7944
rect 929 7880 993 7944
rect 1010 7880 1074 7944
rect 1091 7880 1155 7944
rect 1172 7880 1236 7944
rect 1253 7880 1317 7944
rect 1334 7880 1398 7944
rect 1415 7880 1479 7944
rect 1496 7880 1560 7944
rect 1577 7880 1641 7944
rect 1658 7880 1722 7944
rect 1739 7880 1803 7944
rect 1820 7880 1884 7944
rect 1901 7880 1965 7944
rect 1982 7880 2046 7944
rect 2063 7880 2127 7944
rect 2144 7880 2208 7944
rect 2225 7880 2289 7944
rect 2306 7880 2370 7944
rect 2387 7880 2451 7944
rect 2468 7880 2532 7944
rect 2549 7880 2613 7944
rect 2630 7880 2694 7944
rect 2711 7880 2775 7944
rect 2792 7880 2856 7944
rect 2873 7880 2937 7944
rect 2954 7880 3018 7944
rect 3035 7880 3099 7944
rect 3116 7880 3180 7944
rect 3197 7880 3261 7944
rect 3278 7880 3342 7944
rect 3359 7880 3423 7944
rect 3440 7880 3504 7944
rect 3521 7880 3585 7944
rect 3602 7880 3666 7944
rect 3683 7880 3747 7944
rect 3764 7880 3828 7944
rect 3845 7880 3909 7944
rect 3926 7880 3990 7944
rect 4007 7880 4071 7944
rect 4088 7880 4152 7944
rect 4169 7880 4233 7944
rect 4249 7880 4313 7944
rect 4329 7880 4393 7944
rect 4409 7880 4473 7944
rect 4489 7880 4553 7944
rect 4569 7880 4633 7944
rect 4649 7880 4713 7944
rect 4729 7880 4793 7944
rect 4809 7880 4873 7944
rect 200 7792 264 7856
rect 281 7792 345 7856
rect 362 7792 426 7856
rect 443 7792 507 7856
rect 524 7792 588 7856
rect 605 7792 669 7856
rect 686 7792 750 7856
rect 767 7792 831 7856
rect 848 7792 912 7856
rect 929 7792 993 7856
rect 1010 7792 1074 7856
rect 1091 7792 1155 7856
rect 1172 7792 1236 7856
rect 1253 7792 1317 7856
rect 1334 7792 1398 7856
rect 1415 7792 1479 7856
rect 1496 7792 1560 7856
rect 1577 7792 1641 7856
rect 1658 7792 1722 7856
rect 1739 7792 1803 7856
rect 1820 7792 1884 7856
rect 1901 7792 1965 7856
rect 1982 7792 2046 7856
rect 2063 7792 2127 7856
rect 2144 7792 2208 7856
rect 2225 7792 2289 7856
rect 2306 7792 2370 7856
rect 2387 7792 2451 7856
rect 2468 7792 2532 7856
rect 2549 7792 2613 7856
rect 2630 7792 2694 7856
rect 2711 7792 2775 7856
rect 2792 7792 2856 7856
rect 2873 7792 2937 7856
rect 2954 7792 3018 7856
rect 3035 7792 3099 7856
rect 3116 7792 3180 7856
rect 3197 7792 3261 7856
rect 3278 7792 3342 7856
rect 3359 7792 3423 7856
rect 3440 7792 3504 7856
rect 3521 7792 3585 7856
rect 3602 7792 3666 7856
rect 3683 7792 3747 7856
rect 3764 7792 3828 7856
rect 3845 7792 3909 7856
rect 3926 7792 3990 7856
rect 4007 7792 4071 7856
rect 4088 7792 4152 7856
rect 4169 7792 4233 7856
rect 4249 7792 4313 7856
rect 4329 7792 4393 7856
rect 4409 7792 4473 7856
rect 4489 7792 4553 7856
rect 4569 7792 4633 7856
rect 4649 7792 4713 7856
rect 4729 7792 4793 7856
rect 4809 7792 4873 7856
rect 200 7704 264 7768
rect 281 7704 345 7768
rect 362 7704 426 7768
rect 443 7704 507 7768
rect 524 7704 588 7768
rect 605 7704 669 7768
rect 686 7704 750 7768
rect 767 7704 831 7768
rect 848 7704 912 7768
rect 929 7704 993 7768
rect 1010 7704 1074 7768
rect 1091 7704 1155 7768
rect 1172 7704 1236 7768
rect 1253 7704 1317 7768
rect 1334 7704 1398 7768
rect 1415 7704 1479 7768
rect 1496 7704 1560 7768
rect 1577 7704 1641 7768
rect 1658 7704 1722 7768
rect 1739 7704 1803 7768
rect 1820 7704 1884 7768
rect 1901 7704 1965 7768
rect 1982 7704 2046 7768
rect 2063 7704 2127 7768
rect 2144 7704 2208 7768
rect 2225 7704 2289 7768
rect 2306 7704 2370 7768
rect 2387 7704 2451 7768
rect 2468 7704 2532 7768
rect 2549 7704 2613 7768
rect 2630 7704 2694 7768
rect 2711 7704 2775 7768
rect 2792 7704 2856 7768
rect 2873 7704 2937 7768
rect 2954 7704 3018 7768
rect 3035 7704 3099 7768
rect 3116 7704 3180 7768
rect 3197 7704 3261 7768
rect 3278 7704 3342 7768
rect 3359 7704 3423 7768
rect 3440 7704 3504 7768
rect 3521 7704 3585 7768
rect 3602 7704 3666 7768
rect 3683 7704 3747 7768
rect 3764 7704 3828 7768
rect 3845 7704 3909 7768
rect 3926 7704 3990 7768
rect 4007 7704 4071 7768
rect 4088 7704 4152 7768
rect 4169 7704 4233 7768
rect 4249 7704 4313 7768
rect 4329 7704 4393 7768
rect 4409 7704 4473 7768
rect 4489 7704 4553 7768
rect 4569 7704 4633 7768
rect 4649 7704 4713 7768
rect 4729 7704 4793 7768
rect 4809 7704 4873 7768
rect 200 7616 264 7680
rect 281 7616 345 7680
rect 362 7616 426 7680
rect 443 7616 507 7680
rect 524 7616 588 7680
rect 605 7616 669 7680
rect 686 7616 750 7680
rect 767 7616 831 7680
rect 848 7616 912 7680
rect 929 7616 993 7680
rect 1010 7616 1074 7680
rect 1091 7616 1155 7680
rect 1172 7616 1236 7680
rect 1253 7616 1317 7680
rect 1334 7616 1398 7680
rect 1415 7616 1479 7680
rect 1496 7616 1560 7680
rect 1577 7616 1641 7680
rect 1658 7616 1722 7680
rect 1739 7616 1803 7680
rect 1820 7616 1884 7680
rect 1901 7616 1965 7680
rect 1982 7616 2046 7680
rect 2063 7616 2127 7680
rect 2144 7616 2208 7680
rect 2225 7616 2289 7680
rect 2306 7616 2370 7680
rect 2387 7616 2451 7680
rect 2468 7616 2532 7680
rect 2549 7616 2613 7680
rect 2630 7616 2694 7680
rect 2711 7616 2775 7680
rect 2792 7616 2856 7680
rect 2873 7616 2937 7680
rect 2954 7616 3018 7680
rect 3035 7616 3099 7680
rect 3116 7616 3180 7680
rect 3197 7616 3261 7680
rect 3278 7616 3342 7680
rect 3359 7616 3423 7680
rect 3440 7616 3504 7680
rect 3521 7616 3585 7680
rect 3602 7616 3666 7680
rect 3683 7616 3747 7680
rect 3764 7616 3828 7680
rect 3845 7616 3909 7680
rect 3926 7616 3990 7680
rect 4007 7616 4071 7680
rect 4088 7616 4152 7680
rect 4169 7616 4233 7680
rect 4249 7616 4313 7680
rect 4329 7616 4393 7680
rect 4409 7616 4473 7680
rect 4489 7616 4553 7680
rect 4569 7616 4633 7680
rect 4649 7616 4713 7680
rect 4729 7616 4793 7680
rect 4809 7616 4873 7680
rect 200 7528 264 7592
rect 281 7528 345 7592
rect 362 7528 426 7592
rect 443 7528 507 7592
rect 524 7528 588 7592
rect 605 7528 669 7592
rect 686 7528 750 7592
rect 767 7528 831 7592
rect 848 7528 912 7592
rect 929 7528 993 7592
rect 1010 7528 1074 7592
rect 1091 7528 1155 7592
rect 1172 7528 1236 7592
rect 1253 7528 1317 7592
rect 1334 7528 1398 7592
rect 1415 7528 1479 7592
rect 1496 7528 1560 7592
rect 1577 7528 1641 7592
rect 1658 7528 1722 7592
rect 1739 7528 1803 7592
rect 1820 7528 1884 7592
rect 1901 7528 1965 7592
rect 1982 7528 2046 7592
rect 2063 7528 2127 7592
rect 2144 7528 2208 7592
rect 2225 7528 2289 7592
rect 2306 7528 2370 7592
rect 2387 7528 2451 7592
rect 2468 7528 2532 7592
rect 2549 7528 2613 7592
rect 2630 7528 2694 7592
rect 2711 7528 2775 7592
rect 2792 7528 2856 7592
rect 2873 7528 2937 7592
rect 2954 7528 3018 7592
rect 3035 7528 3099 7592
rect 3116 7528 3180 7592
rect 3197 7528 3261 7592
rect 3278 7528 3342 7592
rect 3359 7528 3423 7592
rect 3440 7528 3504 7592
rect 3521 7528 3585 7592
rect 3602 7528 3666 7592
rect 3683 7528 3747 7592
rect 3764 7528 3828 7592
rect 3845 7528 3909 7592
rect 3926 7528 3990 7592
rect 4007 7528 4071 7592
rect 4088 7528 4152 7592
rect 4169 7528 4233 7592
rect 4249 7528 4313 7592
rect 4329 7528 4393 7592
rect 4409 7528 4473 7592
rect 4489 7528 4553 7592
rect 4569 7528 4633 7592
rect 4649 7528 4713 7592
rect 4729 7528 4793 7592
rect 4809 7528 4873 7592
rect 200 7440 264 7504
rect 281 7440 345 7504
rect 362 7440 426 7504
rect 443 7440 507 7504
rect 524 7440 588 7504
rect 605 7440 669 7504
rect 686 7440 750 7504
rect 767 7440 831 7504
rect 848 7440 912 7504
rect 929 7440 993 7504
rect 1010 7440 1074 7504
rect 1091 7440 1155 7504
rect 1172 7440 1236 7504
rect 1253 7440 1317 7504
rect 1334 7440 1398 7504
rect 1415 7440 1479 7504
rect 1496 7440 1560 7504
rect 1577 7440 1641 7504
rect 1658 7440 1722 7504
rect 1739 7440 1803 7504
rect 1820 7440 1884 7504
rect 1901 7440 1965 7504
rect 1982 7440 2046 7504
rect 2063 7440 2127 7504
rect 2144 7440 2208 7504
rect 2225 7440 2289 7504
rect 2306 7440 2370 7504
rect 2387 7440 2451 7504
rect 2468 7440 2532 7504
rect 2549 7440 2613 7504
rect 2630 7440 2694 7504
rect 2711 7440 2775 7504
rect 2792 7440 2856 7504
rect 2873 7440 2937 7504
rect 2954 7440 3018 7504
rect 3035 7440 3099 7504
rect 3116 7440 3180 7504
rect 3197 7440 3261 7504
rect 3278 7440 3342 7504
rect 3359 7440 3423 7504
rect 3440 7440 3504 7504
rect 3521 7440 3585 7504
rect 3602 7440 3666 7504
rect 3683 7440 3747 7504
rect 3764 7440 3828 7504
rect 3845 7440 3909 7504
rect 3926 7440 3990 7504
rect 4007 7440 4071 7504
rect 4088 7440 4152 7504
rect 4169 7440 4233 7504
rect 4249 7440 4313 7504
rect 4329 7440 4393 7504
rect 4409 7440 4473 7504
rect 4489 7440 4553 7504
rect 4569 7440 4633 7504
rect 4649 7440 4713 7504
rect 4729 7440 4793 7504
rect 4809 7440 4873 7504
rect 200 7352 264 7416
rect 281 7352 345 7416
rect 362 7352 426 7416
rect 443 7352 507 7416
rect 524 7352 588 7416
rect 605 7352 669 7416
rect 686 7352 750 7416
rect 767 7352 831 7416
rect 848 7352 912 7416
rect 929 7352 993 7416
rect 1010 7352 1074 7416
rect 1091 7352 1155 7416
rect 1172 7352 1236 7416
rect 1253 7352 1317 7416
rect 1334 7352 1398 7416
rect 1415 7352 1479 7416
rect 1496 7352 1560 7416
rect 1577 7352 1641 7416
rect 1658 7352 1722 7416
rect 1739 7352 1803 7416
rect 1820 7352 1884 7416
rect 1901 7352 1965 7416
rect 1982 7352 2046 7416
rect 2063 7352 2127 7416
rect 2144 7352 2208 7416
rect 2225 7352 2289 7416
rect 2306 7352 2370 7416
rect 2387 7352 2451 7416
rect 2468 7352 2532 7416
rect 2549 7352 2613 7416
rect 2630 7352 2694 7416
rect 2711 7352 2775 7416
rect 2792 7352 2856 7416
rect 2873 7352 2937 7416
rect 2954 7352 3018 7416
rect 3035 7352 3099 7416
rect 3116 7352 3180 7416
rect 3197 7352 3261 7416
rect 3278 7352 3342 7416
rect 3359 7352 3423 7416
rect 3440 7352 3504 7416
rect 3521 7352 3585 7416
rect 3602 7352 3666 7416
rect 3683 7352 3747 7416
rect 3764 7352 3828 7416
rect 3845 7352 3909 7416
rect 3926 7352 3990 7416
rect 4007 7352 4071 7416
rect 4088 7352 4152 7416
rect 4169 7352 4233 7416
rect 4249 7352 4313 7416
rect 4329 7352 4393 7416
rect 4409 7352 4473 7416
rect 4489 7352 4553 7416
rect 4569 7352 4633 7416
rect 4649 7352 4713 7416
rect 4729 7352 4793 7416
rect 4809 7352 4873 7416
rect 10084 7968 10148 8032
rect 10166 7968 10230 8032
rect 10248 7968 10312 8032
rect 10330 7968 10394 8032
rect 10412 7968 10476 8032
rect 10494 7968 10558 8032
rect 10576 7968 10640 8032
rect 10657 7968 10721 8032
rect 10738 7968 10802 8032
rect 10819 7968 10883 8032
rect 10900 7968 10964 8032
rect 10981 7968 11045 8032
rect 11062 7968 11126 8032
rect 11143 7968 11207 8032
rect 11224 7968 11288 8032
rect 11305 7968 11369 8032
rect 11386 7968 11450 8032
rect 11467 7968 11531 8032
rect 11548 7968 11612 8032
rect 11629 7968 11693 8032
rect 11710 7968 11774 8032
rect 11791 7968 11855 8032
rect 11872 7968 11936 8032
rect 11953 7968 12017 8032
rect 12034 7968 12098 8032
rect 12115 7968 12179 8032
rect 12196 7968 12260 8032
rect 12277 7968 12341 8032
rect 12358 7968 12422 8032
rect 12439 7968 12503 8032
rect 12520 7968 12584 8032
rect 12601 7968 12665 8032
rect 12682 7968 12746 8032
rect 12763 7968 12827 8032
rect 12844 7968 12908 8032
rect 12925 7968 12989 8032
rect 13006 7968 13070 8032
rect 13087 7968 13151 8032
rect 13168 7968 13232 8032
rect 13249 7968 13313 8032
rect 13330 7968 13394 8032
rect 13411 7968 13475 8032
rect 13492 7968 13556 8032
rect 13573 7968 13637 8032
rect 13654 7968 13718 8032
rect 13735 7968 13799 8032
rect 13816 7968 13880 8032
rect 13897 7968 13961 8032
rect 13978 7968 14042 8032
rect 14059 7968 14123 8032
rect 14140 7968 14204 8032
rect 14221 7968 14285 8032
rect 14302 7968 14366 8032
rect 14383 7968 14447 8032
rect 14464 7968 14528 8032
rect 14545 7968 14609 8032
rect 14626 7968 14690 8032
rect 14707 7968 14771 8032
rect 14788 7968 14852 8032
rect 10084 7880 10148 7944
rect 10166 7880 10230 7944
rect 10248 7880 10312 7944
rect 10330 7880 10394 7944
rect 10412 7880 10476 7944
rect 10494 7880 10558 7944
rect 10576 7880 10640 7944
rect 10657 7880 10721 7944
rect 10738 7880 10802 7944
rect 10819 7880 10883 7944
rect 10900 7880 10964 7944
rect 10981 7880 11045 7944
rect 11062 7880 11126 7944
rect 11143 7880 11207 7944
rect 11224 7880 11288 7944
rect 11305 7880 11369 7944
rect 11386 7880 11450 7944
rect 11467 7880 11531 7944
rect 11548 7880 11612 7944
rect 11629 7880 11693 7944
rect 11710 7880 11774 7944
rect 11791 7880 11855 7944
rect 11872 7880 11936 7944
rect 11953 7880 12017 7944
rect 12034 7880 12098 7944
rect 12115 7880 12179 7944
rect 12196 7880 12260 7944
rect 12277 7880 12341 7944
rect 12358 7880 12422 7944
rect 12439 7880 12503 7944
rect 12520 7880 12584 7944
rect 12601 7880 12665 7944
rect 12682 7880 12746 7944
rect 12763 7880 12827 7944
rect 12844 7880 12908 7944
rect 12925 7880 12989 7944
rect 13006 7880 13070 7944
rect 13087 7880 13151 7944
rect 13168 7880 13232 7944
rect 13249 7880 13313 7944
rect 13330 7880 13394 7944
rect 13411 7880 13475 7944
rect 13492 7880 13556 7944
rect 13573 7880 13637 7944
rect 13654 7880 13718 7944
rect 13735 7880 13799 7944
rect 13816 7880 13880 7944
rect 13897 7880 13961 7944
rect 13978 7880 14042 7944
rect 14059 7880 14123 7944
rect 14140 7880 14204 7944
rect 14221 7880 14285 7944
rect 14302 7880 14366 7944
rect 14383 7880 14447 7944
rect 14464 7880 14528 7944
rect 14545 7880 14609 7944
rect 14626 7880 14690 7944
rect 14707 7880 14771 7944
rect 14788 7880 14852 7944
rect 10084 7792 10148 7856
rect 10166 7792 10230 7856
rect 10248 7792 10312 7856
rect 10330 7792 10394 7856
rect 10412 7792 10476 7856
rect 10494 7792 10558 7856
rect 10576 7792 10640 7856
rect 10657 7792 10721 7856
rect 10738 7792 10802 7856
rect 10819 7792 10883 7856
rect 10900 7792 10964 7856
rect 10981 7792 11045 7856
rect 11062 7792 11126 7856
rect 11143 7792 11207 7856
rect 11224 7792 11288 7856
rect 11305 7792 11369 7856
rect 11386 7792 11450 7856
rect 11467 7792 11531 7856
rect 11548 7792 11612 7856
rect 11629 7792 11693 7856
rect 11710 7792 11774 7856
rect 11791 7792 11855 7856
rect 11872 7792 11936 7856
rect 11953 7792 12017 7856
rect 12034 7792 12098 7856
rect 12115 7792 12179 7856
rect 12196 7792 12260 7856
rect 12277 7792 12341 7856
rect 12358 7792 12422 7856
rect 12439 7792 12503 7856
rect 12520 7792 12584 7856
rect 12601 7792 12665 7856
rect 12682 7792 12746 7856
rect 12763 7792 12827 7856
rect 12844 7792 12908 7856
rect 12925 7792 12989 7856
rect 13006 7792 13070 7856
rect 13087 7792 13151 7856
rect 13168 7792 13232 7856
rect 13249 7792 13313 7856
rect 13330 7792 13394 7856
rect 13411 7792 13475 7856
rect 13492 7792 13556 7856
rect 13573 7792 13637 7856
rect 13654 7792 13718 7856
rect 13735 7792 13799 7856
rect 13816 7792 13880 7856
rect 13897 7792 13961 7856
rect 13978 7792 14042 7856
rect 14059 7792 14123 7856
rect 14140 7792 14204 7856
rect 14221 7792 14285 7856
rect 14302 7792 14366 7856
rect 14383 7792 14447 7856
rect 14464 7792 14528 7856
rect 14545 7792 14609 7856
rect 14626 7792 14690 7856
rect 14707 7792 14771 7856
rect 14788 7792 14852 7856
rect 10084 7704 10148 7768
rect 10166 7704 10230 7768
rect 10248 7704 10312 7768
rect 10330 7704 10394 7768
rect 10412 7704 10476 7768
rect 10494 7704 10558 7768
rect 10576 7704 10640 7768
rect 10657 7704 10721 7768
rect 10738 7704 10802 7768
rect 10819 7704 10883 7768
rect 10900 7704 10964 7768
rect 10981 7704 11045 7768
rect 11062 7704 11126 7768
rect 11143 7704 11207 7768
rect 11224 7704 11288 7768
rect 11305 7704 11369 7768
rect 11386 7704 11450 7768
rect 11467 7704 11531 7768
rect 11548 7704 11612 7768
rect 11629 7704 11693 7768
rect 11710 7704 11774 7768
rect 11791 7704 11855 7768
rect 11872 7704 11936 7768
rect 11953 7704 12017 7768
rect 12034 7704 12098 7768
rect 12115 7704 12179 7768
rect 12196 7704 12260 7768
rect 12277 7704 12341 7768
rect 12358 7704 12422 7768
rect 12439 7704 12503 7768
rect 12520 7704 12584 7768
rect 12601 7704 12665 7768
rect 12682 7704 12746 7768
rect 12763 7704 12827 7768
rect 12844 7704 12908 7768
rect 12925 7704 12989 7768
rect 13006 7704 13070 7768
rect 13087 7704 13151 7768
rect 13168 7704 13232 7768
rect 13249 7704 13313 7768
rect 13330 7704 13394 7768
rect 13411 7704 13475 7768
rect 13492 7704 13556 7768
rect 13573 7704 13637 7768
rect 13654 7704 13718 7768
rect 13735 7704 13799 7768
rect 13816 7704 13880 7768
rect 13897 7704 13961 7768
rect 13978 7704 14042 7768
rect 14059 7704 14123 7768
rect 14140 7704 14204 7768
rect 14221 7704 14285 7768
rect 14302 7704 14366 7768
rect 14383 7704 14447 7768
rect 14464 7704 14528 7768
rect 14545 7704 14609 7768
rect 14626 7704 14690 7768
rect 14707 7704 14771 7768
rect 14788 7704 14852 7768
rect 10084 7616 10148 7680
rect 10166 7616 10230 7680
rect 10248 7616 10312 7680
rect 10330 7616 10394 7680
rect 10412 7616 10476 7680
rect 10494 7616 10558 7680
rect 10576 7616 10640 7680
rect 10657 7616 10721 7680
rect 10738 7616 10802 7680
rect 10819 7616 10883 7680
rect 10900 7616 10964 7680
rect 10981 7616 11045 7680
rect 11062 7616 11126 7680
rect 11143 7616 11207 7680
rect 11224 7616 11288 7680
rect 11305 7616 11369 7680
rect 11386 7616 11450 7680
rect 11467 7616 11531 7680
rect 11548 7616 11612 7680
rect 11629 7616 11693 7680
rect 11710 7616 11774 7680
rect 11791 7616 11855 7680
rect 11872 7616 11936 7680
rect 11953 7616 12017 7680
rect 12034 7616 12098 7680
rect 12115 7616 12179 7680
rect 12196 7616 12260 7680
rect 12277 7616 12341 7680
rect 12358 7616 12422 7680
rect 12439 7616 12503 7680
rect 12520 7616 12584 7680
rect 12601 7616 12665 7680
rect 12682 7616 12746 7680
rect 12763 7616 12827 7680
rect 12844 7616 12908 7680
rect 12925 7616 12989 7680
rect 13006 7616 13070 7680
rect 13087 7616 13151 7680
rect 13168 7616 13232 7680
rect 13249 7616 13313 7680
rect 13330 7616 13394 7680
rect 13411 7616 13475 7680
rect 13492 7616 13556 7680
rect 13573 7616 13637 7680
rect 13654 7616 13718 7680
rect 13735 7616 13799 7680
rect 13816 7616 13880 7680
rect 13897 7616 13961 7680
rect 13978 7616 14042 7680
rect 14059 7616 14123 7680
rect 14140 7616 14204 7680
rect 14221 7616 14285 7680
rect 14302 7616 14366 7680
rect 14383 7616 14447 7680
rect 14464 7616 14528 7680
rect 14545 7616 14609 7680
rect 14626 7616 14690 7680
rect 14707 7616 14771 7680
rect 14788 7616 14852 7680
rect 10084 7528 10148 7592
rect 10166 7528 10230 7592
rect 10248 7528 10312 7592
rect 10330 7528 10394 7592
rect 10412 7528 10476 7592
rect 10494 7528 10558 7592
rect 10576 7528 10640 7592
rect 10657 7528 10721 7592
rect 10738 7528 10802 7592
rect 10819 7528 10883 7592
rect 10900 7528 10964 7592
rect 10981 7528 11045 7592
rect 11062 7528 11126 7592
rect 11143 7528 11207 7592
rect 11224 7528 11288 7592
rect 11305 7528 11369 7592
rect 11386 7528 11450 7592
rect 11467 7528 11531 7592
rect 11548 7528 11612 7592
rect 11629 7528 11693 7592
rect 11710 7528 11774 7592
rect 11791 7528 11855 7592
rect 11872 7528 11936 7592
rect 11953 7528 12017 7592
rect 12034 7528 12098 7592
rect 12115 7528 12179 7592
rect 12196 7528 12260 7592
rect 12277 7528 12341 7592
rect 12358 7528 12422 7592
rect 12439 7528 12503 7592
rect 12520 7528 12584 7592
rect 12601 7528 12665 7592
rect 12682 7528 12746 7592
rect 12763 7528 12827 7592
rect 12844 7528 12908 7592
rect 12925 7528 12989 7592
rect 13006 7528 13070 7592
rect 13087 7528 13151 7592
rect 13168 7528 13232 7592
rect 13249 7528 13313 7592
rect 13330 7528 13394 7592
rect 13411 7528 13475 7592
rect 13492 7528 13556 7592
rect 13573 7528 13637 7592
rect 13654 7528 13718 7592
rect 13735 7528 13799 7592
rect 13816 7528 13880 7592
rect 13897 7528 13961 7592
rect 13978 7528 14042 7592
rect 14059 7528 14123 7592
rect 14140 7528 14204 7592
rect 14221 7528 14285 7592
rect 14302 7528 14366 7592
rect 14383 7528 14447 7592
rect 14464 7528 14528 7592
rect 14545 7528 14609 7592
rect 14626 7528 14690 7592
rect 14707 7528 14771 7592
rect 14788 7528 14852 7592
rect 10084 7440 10148 7504
rect 10166 7440 10230 7504
rect 10248 7440 10312 7504
rect 10330 7440 10394 7504
rect 10412 7440 10476 7504
rect 10494 7440 10558 7504
rect 10576 7440 10640 7504
rect 10657 7440 10721 7504
rect 10738 7440 10802 7504
rect 10819 7440 10883 7504
rect 10900 7440 10964 7504
rect 10981 7440 11045 7504
rect 11062 7440 11126 7504
rect 11143 7440 11207 7504
rect 11224 7440 11288 7504
rect 11305 7440 11369 7504
rect 11386 7440 11450 7504
rect 11467 7440 11531 7504
rect 11548 7440 11612 7504
rect 11629 7440 11693 7504
rect 11710 7440 11774 7504
rect 11791 7440 11855 7504
rect 11872 7440 11936 7504
rect 11953 7440 12017 7504
rect 12034 7440 12098 7504
rect 12115 7440 12179 7504
rect 12196 7440 12260 7504
rect 12277 7440 12341 7504
rect 12358 7440 12422 7504
rect 12439 7440 12503 7504
rect 12520 7440 12584 7504
rect 12601 7440 12665 7504
rect 12682 7440 12746 7504
rect 12763 7440 12827 7504
rect 12844 7440 12908 7504
rect 12925 7440 12989 7504
rect 13006 7440 13070 7504
rect 13087 7440 13151 7504
rect 13168 7440 13232 7504
rect 13249 7440 13313 7504
rect 13330 7440 13394 7504
rect 13411 7440 13475 7504
rect 13492 7440 13556 7504
rect 13573 7440 13637 7504
rect 13654 7440 13718 7504
rect 13735 7440 13799 7504
rect 13816 7440 13880 7504
rect 13897 7440 13961 7504
rect 13978 7440 14042 7504
rect 14059 7440 14123 7504
rect 14140 7440 14204 7504
rect 14221 7440 14285 7504
rect 14302 7440 14366 7504
rect 14383 7440 14447 7504
rect 14464 7440 14528 7504
rect 14545 7440 14609 7504
rect 14626 7440 14690 7504
rect 14707 7440 14771 7504
rect 14788 7440 14852 7504
rect 10084 7352 10148 7416
rect 10166 7352 10230 7416
rect 10248 7352 10312 7416
rect 10330 7352 10394 7416
rect 10412 7352 10476 7416
rect 10494 7352 10558 7416
rect 10576 7352 10640 7416
rect 10657 7352 10721 7416
rect 10738 7352 10802 7416
rect 10819 7352 10883 7416
rect 10900 7352 10964 7416
rect 10981 7352 11045 7416
rect 11062 7352 11126 7416
rect 11143 7352 11207 7416
rect 11224 7352 11288 7416
rect 11305 7352 11369 7416
rect 11386 7352 11450 7416
rect 11467 7352 11531 7416
rect 11548 7352 11612 7416
rect 11629 7352 11693 7416
rect 11710 7352 11774 7416
rect 11791 7352 11855 7416
rect 11872 7352 11936 7416
rect 11953 7352 12017 7416
rect 12034 7352 12098 7416
rect 12115 7352 12179 7416
rect 12196 7352 12260 7416
rect 12277 7352 12341 7416
rect 12358 7352 12422 7416
rect 12439 7352 12503 7416
rect 12520 7352 12584 7416
rect 12601 7352 12665 7416
rect 12682 7352 12746 7416
rect 12763 7352 12827 7416
rect 12844 7352 12908 7416
rect 12925 7352 12989 7416
rect 13006 7352 13070 7416
rect 13087 7352 13151 7416
rect 13168 7352 13232 7416
rect 13249 7352 13313 7416
rect 13330 7352 13394 7416
rect 13411 7352 13475 7416
rect 13492 7352 13556 7416
rect 13573 7352 13637 7416
rect 13654 7352 13718 7416
rect 13735 7352 13799 7416
rect 13816 7352 13880 7416
rect 13897 7352 13961 7416
rect 13978 7352 14042 7416
rect 14059 7352 14123 7416
rect 14140 7352 14204 7416
rect 14221 7352 14285 7416
rect 14302 7352 14366 7416
rect 14383 7352 14447 7416
rect 14464 7352 14528 7416
rect 14545 7352 14609 7416
rect 14626 7352 14690 7416
rect 14707 7352 14771 7416
rect 14788 7352 14852 7416
<< metal4 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 19000
rect 14746 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 11647 254 12537
rect 14746 11647 15000 12537
rect 0 11346 4874 11347
rect 0 11282 112 11346
rect 176 11282 193 11346
rect 257 11282 274 11346
rect 338 11282 355 11346
rect 419 11282 436 11346
rect 500 11282 517 11346
rect 581 11282 598 11346
rect 662 11282 679 11346
rect 743 11282 760 11346
rect 824 11282 841 11346
rect 905 11282 922 11346
rect 986 11282 1003 11346
rect 1067 11282 1084 11346
rect 1148 11282 1165 11346
rect 1229 11282 1246 11346
rect 1310 11282 1327 11346
rect 1391 11282 1408 11346
rect 1472 11282 1489 11346
rect 1553 11282 1570 11346
rect 1634 11282 1651 11346
rect 1715 11282 1732 11346
rect 1796 11282 1813 11346
rect 1877 11282 1894 11346
rect 1958 11282 1975 11346
rect 2039 11282 2056 11346
rect 2120 11282 2137 11346
rect 2201 11282 2218 11346
rect 2282 11282 2299 11346
rect 2363 11282 2380 11346
rect 2444 11282 2461 11346
rect 2525 11282 2542 11346
rect 2606 11282 2623 11346
rect 2687 11282 2704 11346
rect 2768 11282 2785 11346
rect 2849 11282 2866 11346
rect 2930 11282 2947 11346
rect 3011 11282 3028 11346
rect 3092 11282 3109 11346
rect 3173 11282 3190 11346
rect 3254 11282 3271 11346
rect 3335 11282 3352 11346
rect 3416 11282 3433 11346
rect 3497 11282 3514 11346
rect 3578 11282 3595 11346
rect 3659 11282 3676 11346
rect 3740 11282 3757 11346
rect 3821 11282 3838 11346
rect 3902 11282 3919 11346
rect 3983 11282 4000 11346
rect 4064 11282 4081 11346
rect 4145 11282 4162 11346
rect 4226 11282 4243 11346
rect 4307 11282 4324 11346
rect 4388 11282 4405 11346
rect 4469 11282 4486 11346
rect 4550 11282 4567 11346
rect 4631 11282 4648 11346
rect 4712 11282 4729 11346
rect 4793 11282 4809 11346
rect 4873 11282 4874 11346
rect 0 11281 4874 11282
rect 10083 11346 15000 11347
rect 10083 11282 10084 11346
rect 10148 11282 10165 11346
rect 10229 11282 10246 11346
rect 10310 11282 10327 11346
rect 10391 11282 10408 11346
rect 10472 11282 10489 11346
rect 10553 11282 10570 11346
rect 10634 11282 10651 11346
rect 10715 11282 10732 11346
rect 10796 11282 10813 11346
rect 10877 11282 10894 11346
rect 10958 11282 10975 11346
rect 11039 11282 11056 11346
rect 11120 11282 11137 11346
rect 11201 11282 11218 11346
rect 11282 11282 11299 11346
rect 11363 11282 11380 11346
rect 11444 11282 11461 11346
rect 11525 11282 11542 11346
rect 11606 11282 11623 11346
rect 11687 11282 11704 11346
rect 11768 11282 11785 11346
rect 11849 11282 11866 11346
rect 11930 11282 11947 11346
rect 12011 11282 12028 11346
rect 12092 11282 12109 11346
rect 12173 11282 12190 11346
rect 12254 11282 12271 11346
rect 12335 11282 12352 11346
rect 12416 11282 12433 11346
rect 12497 11282 12514 11346
rect 12578 11282 12595 11346
rect 12659 11282 12676 11346
rect 12740 11282 12757 11346
rect 12821 11282 12838 11346
rect 12902 11282 12919 11346
rect 12983 11282 13000 11346
rect 13064 11282 13081 11346
rect 13145 11282 13162 11346
rect 13226 11282 13243 11346
rect 13307 11282 13324 11346
rect 13388 11282 13405 11346
rect 13469 11282 13486 11346
rect 13550 11282 13567 11346
rect 13631 11282 13648 11346
rect 13712 11282 13729 11346
rect 13793 11282 13810 11346
rect 13874 11282 13891 11346
rect 13955 11282 13972 11346
rect 14036 11282 14053 11346
rect 14117 11282 14134 11346
rect 14198 11282 14215 11346
rect 14279 11282 14296 11346
rect 14360 11282 14378 11346
rect 14442 11282 14460 11346
rect 14524 11282 14542 11346
rect 14606 11282 14624 11346
rect 14688 11282 14706 11346
rect 14770 11282 14788 11346
rect 14852 11282 15000 11346
rect 10083 11281 15000 11282
rect 0 10625 254 11221
rect 14746 10625 15000 11221
rect 0 10563 4874 10565
rect 0 10499 105 10563
rect 169 10499 187 10563
rect 251 10499 269 10563
rect 333 10499 351 10563
rect 415 10499 433 10563
rect 497 10499 515 10563
rect 579 10499 597 10563
rect 661 10499 678 10563
rect 742 10499 759 10563
rect 823 10499 840 10563
rect 904 10499 921 10563
rect 985 10499 1002 10563
rect 1066 10499 1083 10563
rect 1147 10499 1164 10563
rect 1228 10499 1245 10563
rect 1309 10499 1326 10563
rect 1390 10499 1407 10563
rect 1471 10499 1488 10563
rect 1552 10499 1569 10563
rect 1633 10499 1650 10563
rect 1714 10499 1731 10563
rect 1795 10499 1812 10563
rect 1876 10499 1893 10563
rect 1957 10499 1974 10563
rect 2038 10499 2055 10563
rect 2119 10499 2136 10563
rect 2200 10499 2217 10563
rect 2281 10499 2298 10563
rect 2362 10499 2379 10563
rect 2443 10499 2460 10563
rect 2524 10499 2541 10563
rect 2605 10499 2622 10563
rect 2686 10499 2703 10563
rect 2767 10499 2784 10563
rect 2848 10499 2865 10563
rect 2929 10499 2946 10563
rect 3010 10499 3027 10563
rect 3091 10499 3108 10563
rect 3172 10499 3189 10563
rect 3253 10499 3270 10563
rect 3334 10499 3351 10563
rect 3415 10499 3432 10563
rect 3496 10499 3513 10563
rect 3577 10499 3594 10563
rect 3658 10499 3675 10563
rect 3739 10499 3756 10563
rect 3820 10499 3837 10563
rect 3901 10499 3918 10563
rect 3982 10499 3999 10563
rect 4063 10499 4080 10563
rect 4144 10499 4161 10563
rect 4225 10499 4242 10563
rect 4306 10499 4323 10563
rect 4387 10499 4404 10563
rect 4468 10499 4485 10563
rect 4549 10499 4566 10563
rect 4630 10499 4647 10563
rect 4711 10499 4728 10563
rect 4792 10499 4809 10563
rect 4873 10499 4874 10563
rect 0 10479 4874 10499
rect 0 10415 105 10479
rect 169 10415 187 10479
rect 251 10415 269 10479
rect 333 10415 351 10479
rect 415 10415 433 10479
rect 497 10415 515 10479
rect 579 10415 597 10479
rect 661 10415 678 10479
rect 742 10415 759 10479
rect 823 10415 840 10479
rect 904 10415 921 10479
rect 985 10415 1002 10479
rect 1066 10415 1083 10479
rect 1147 10415 1164 10479
rect 1228 10415 1245 10479
rect 1309 10415 1326 10479
rect 1390 10415 1407 10479
rect 1471 10415 1488 10479
rect 1552 10415 1569 10479
rect 1633 10415 1650 10479
rect 1714 10415 1731 10479
rect 1795 10415 1812 10479
rect 1876 10415 1893 10479
rect 1957 10415 1974 10479
rect 2038 10415 2055 10479
rect 2119 10415 2136 10479
rect 2200 10415 2217 10479
rect 2281 10415 2298 10479
rect 2362 10415 2379 10479
rect 2443 10415 2460 10479
rect 2524 10415 2541 10479
rect 2605 10415 2622 10479
rect 2686 10415 2703 10479
rect 2767 10415 2784 10479
rect 2848 10415 2865 10479
rect 2929 10415 2946 10479
rect 3010 10415 3027 10479
rect 3091 10415 3108 10479
rect 3172 10415 3189 10479
rect 3253 10415 3270 10479
rect 3334 10415 3351 10479
rect 3415 10415 3432 10479
rect 3496 10415 3513 10479
rect 3577 10415 3594 10479
rect 3658 10415 3675 10479
rect 3739 10415 3756 10479
rect 3820 10415 3837 10479
rect 3901 10415 3918 10479
rect 3982 10415 3999 10479
rect 4063 10415 4080 10479
rect 4144 10415 4161 10479
rect 4225 10415 4242 10479
rect 4306 10415 4323 10479
rect 4387 10415 4404 10479
rect 4468 10415 4485 10479
rect 4549 10415 4566 10479
rect 4630 10415 4647 10479
rect 4711 10415 4728 10479
rect 4792 10415 4809 10479
rect 4873 10415 4874 10479
rect 0 10395 4874 10415
rect 0 10331 105 10395
rect 169 10331 187 10395
rect 251 10331 269 10395
rect 333 10331 351 10395
rect 415 10331 433 10395
rect 497 10331 515 10395
rect 579 10331 597 10395
rect 661 10331 678 10395
rect 742 10331 759 10395
rect 823 10331 840 10395
rect 904 10331 921 10395
rect 985 10331 1002 10395
rect 1066 10331 1083 10395
rect 1147 10331 1164 10395
rect 1228 10331 1245 10395
rect 1309 10331 1326 10395
rect 1390 10331 1407 10395
rect 1471 10331 1488 10395
rect 1552 10331 1569 10395
rect 1633 10331 1650 10395
rect 1714 10331 1731 10395
rect 1795 10331 1812 10395
rect 1876 10331 1893 10395
rect 1957 10331 1974 10395
rect 2038 10331 2055 10395
rect 2119 10331 2136 10395
rect 2200 10331 2217 10395
rect 2281 10331 2298 10395
rect 2362 10331 2379 10395
rect 2443 10331 2460 10395
rect 2524 10331 2541 10395
rect 2605 10331 2622 10395
rect 2686 10331 2703 10395
rect 2767 10331 2784 10395
rect 2848 10331 2865 10395
rect 2929 10331 2946 10395
rect 3010 10331 3027 10395
rect 3091 10331 3108 10395
rect 3172 10331 3189 10395
rect 3253 10331 3270 10395
rect 3334 10331 3351 10395
rect 3415 10331 3432 10395
rect 3496 10331 3513 10395
rect 3577 10331 3594 10395
rect 3658 10331 3675 10395
rect 3739 10331 3756 10395
rect 3820 10331 3837 10395
rect 3901 10331 3918 10395
rect 3982 10331 3999 10395
rect 4063 10331 4080 10395
rect 4144 10331 4161 10395
rect 4225 10331 4242 10395
rect 4306 10331 4323 10395
rect 4387 10331 4404 10395
rect 4468 10331 4485 10395
rect 4549 10331 4566 10395
rect 4630 10331 4647 10395
rect 4711 10331 4728 10395
rect 4792 10331 4809 10395
rect 4873 10331 4874 10395
rect 0 10329 4874 10331
rect 10083 10563 15000 10565
rect 10083 10499 10084 10563
rect 10148 10499 10166 10563
rect 10230 10499 10248 10563
rect 10312 10499 10330 10563
rect 10394 10499 10412 10563
rect 10476 10499 10494 10563
rect 10558 10499 10576 10563
rect 10640 10499 10657 10563
rect 10721 10499 10738 10563
rect 10802 10499 10819 10563
rect 10883 10499 10900 10563
rect 10964 10499 10981 10563
rect 11045 10499 11062 10563
rect 11126 10499 11143 10563
rect 11207 10499 11224 10563
rect 11288 10499 11305 10563
rect 11369 10499 11386 10563
rect 11450 10499 11467 10563
rect 11531 10499 11548 10563
rect 11612 10499 11629 10563
rect 11693 10499 11710 10563
rect 11774 10499 11791 10563
rect 11855 10499 11872 10563
rect 11936 10499 11953 10563
rect 12017 10499 12034 10563
rect 12098 10499 12115 10563
rect 12179 10499 12196 10563
rect 12260 10499 12277 10563
rect 12341 10499 12358 10563
rect 12422 10499 12439 10563
rect 12503 10499 12520 10563
rect 12584 10499 12601 10563
rect 12665 10499 12682 10563
rect 12746 10499 12763 10563
rect 12827 10499 12844 10563
rect 12908 10499 12925 10563
rect 12989 10499 13006 10563
rect 13070 10499 13087 10563
rect 13151 10499 13168 10563
rect 13232 10499 13249 10563
rect 13313 10499 13330 10563
rect 13394 10499 13411 10563
rect 13475 10499 13492 10563
rect 13556 10499 13573 10563
rect 13637 10499 13654 10563
rect 13718 10499 13735 10563
rect 13799 10499 13816 10563
rect 13880 10499 13897 10563
rect 13961 10499 13978 10563
rect 14042 10499 14059 10563
rect 14123 10499 14140 10563
rect 14204 10499 14221 10563
rect 14285 10499 14302 10563
rect 14366 10499 14383 10563
rect 14447 10499 14464 10563
rect 14528 10499 14545 10563
rect 14609 10499 14626 10563
rect 14690 10499 14707 10563
rect 14771 10499 14788 10563
rect 14852 10499 15000 10563
rect 10083 10479 15000 10499
rect 10083 10415 10084 10479
rect 10148 10415 10166 10479
rect 10230 10415 10248 10479
rect 10312 10415 10330 10479
rect 10394 10415 10412 10479
rect 10476 10415 10494 10479
rect 10558 10415 10576 10479
rect 10640 10415 10657 10479
rect 10721 10415 10738 10479
rect 10802 10415 10819 10479
rect 10883 10415 10900 10479
rect 10964 10415 10981 10479
rect 11045 10415 11062 10479
rect 11126 10415 11143 10479
rect 11207 10415 11224 10479
rect 11288 10415 11305 10479
rect 11369 10415 11386 10479
rect 11450 10415 11467 10479
rect 11531 10415 11548 10479
rect 11612 10415 11629 10479
rect 11693 10415 11710 10479
rect 11774 10415 11791 10479
rect 11855 10415 11872 10479
rect 11936 10415 11953 10479
rect 12017 10415 12034 10479
rect 12098 10415 12115 10479
rect 12179 10415 12196 10479
rect 12260 10415 12277 10479
rect 12341 10415 12358 10479
rect 12422 10415 12439 10479
rect 12503 10415 12520 10479
rect 12584 10415 12601 10479
rect 12665 10415 12682 10479
rect 12746 10415 12763 10479
rect 12827 10415 12844 10479
rect 12908 10415 12925 10479
rect 12989 10415 13006 10479
rect 13070 10415 13087 10479
rect 13151 10415 13168 10479
rect 13232 10415 13249 10479
rect 13313 10415 13330 10479
rect 13394 10415 13411 10479
rect 13475 10415 13492 10479
rect 13556 10415 13573 10479
rect 13637 10415 13654 10479
rect 13718 10415 13735 10479
rect 13799 10415 13816 10479
rect 13880 10415 13897 10479
rect 13961 10415 13978 10479
rect 14042 10415 14059 10479
rect 14123 10415 14140 10479
rect 14204 10415 14221 10479
rect 14285 10415 14302 10479
rect 14366 10415 14383 10479
rect 14447 10415 14464 10479
rect 14528 10415 14545 10479
rect 14609 10415 14626 10479
rect 14690 10415 14707 10479
rect 14771 10415 14788 10479
rect 14852 10415 15000 10479
rect 10083 10395 15000 10415
rect 10083 10331 10084 10395
rect 10148 10331 10166 10395
rect 10230 10331 10248 10395
rect 10312 10331 10330 10395
rect 10394 10331 10412 10395
rect 10476 10331 10494 10395
rect 10558 10331 10576 10395
rect 10640 10331 10657 10395
rect 10721 10331 10738 10395
rect 10802 10331 10819 10395
rect 10883 10331 10900 10395
rect 10964 10331 10981 10395
rect 11045 10331 11062 10395
rect 11126 10331 11143 10395
rect 11207 10331 11224 10395
rect 11288 10331 11305 10395
rect 11369 10331 11386 10395
rect 11450 10331 11467 10395
rect 11531 10331 11548 10395
rect 11612 10331 11629 10395
rect 11693 10331 11710 10395
rect 11774 10331 11791 10395
rect 11855 10331 11872 10395
rect 11936 10331 11953 10395
rect 12017 10331 12034 10395
rect 12098 10331 12115 10395
rect 12179 10331 12196 10395
rect 12260 10331 12277 10395
rect 12341 10331 12358 10395
rect 12422 10331 12439 10395
rect 12503 10331 12520 10395
rect 12584 10331 12601 10395
rect 12665 10331 12682 10395
rect 12746 10331 12763 10395
rect 12827 10331 12844 10395
rect 12908 10331 12925 10395
rect 12989 10331 13006 10395
rect 13070 10331 13087 10395
rect 13151 10331 13168 10395
rect 13232 10331 13249 10395
rect 13313 10331 13330 10395
rect 13394 10331 13411 10395
rect 13475 10331 13492 10395
rect 13556 10331 13573 10395
rect 13637 10331 13654 10395
rect 13718 10331 13735 10395
rect 13799 10331 13816 10395
rect 13880 10331 13897 10395
rect 13961 10331 13978 10395
rect 14042 10331 14059 10395
rect 14123 10331 14140 10395
rect 14204 10331 14221 10395
rect 14285 10331 14302 10395
rect 14366 10331 14383 10395
rect 14447 10331 14464 10395
rect 14528 10331 14545 10395
rect 14609 10331 14626 10395
rect 14690 10331 14707 10395
rect 14771 10331 14788 10395
rect 14852 10331 15000 10395
rect 10083 10329 15000 10331
rect 0 9673 254 10269
rect 14746 9673 15000 10269
rect 0 9612 4874 9613
rect 0 9548 112 9612
rect 176 9548 193 9612
rect 257 9548 274 9612
rect 338 9548 355 9612
rect 419 9548 436 9612
rect 500 9548 517 9612
rect 581 9548 598 9612
rect 662 9548 679 9612
rect 743 9548 760 9612
rect 824 9548 841 9612
rect 905 9548 922 9612
rect 986 9548 1003 9612
rect 1067 9548 1084 9612
rect 1148 9548 1165 9612
rect 1229 9548 1246 9612
rect 1310 9548 1327 9612
rect 1391 9548 1408 9612
rect 1472 9548 1489 9612
rect 1553 9548 1570 9612
rect 1634 9548 1651 9612
rect 1715 9548 1732 9612
rect 1796 9548 1813 9612
rect 1877 9548 1894 9612
rect 1958 9548 1975 9612
rect 2039 9548 2056 9612
rect 2120 9548 2137 9612
rect 2201 9548 2218 9612
rect 2282 9548 2299 9612
rect 2363 9548 2380 9612
rect 2444 9548 2461 9612
rect 2525 9548 2542 9612
rect 2606 9548 2623 9612
rect 2687 9548 2704 9612
rect 2768 9548 2785 9612
rect 2849 9548 2866 9612
rect 2930 9548 2947 9612
rect 3011 9548 3028 9612
rect 3092 9548 3109 9612
rect 3173 9548 3190 9612
rect 3254 9548 3271 9612
rect 3335 9548 3352 9612
rect 3416 9548 3433 9612
rect 3497 9548 3514 9612
rect 3578 9548 3595 9612
rect 3659 9548 3676 9612
rect 3740 9548 3757 9612
rect 3821 9548 3838 9612
rect 3902 9548 3919 9612
rect 3983 9548 4000 9612
rect 4064 9548 4081 9612
rect 4145 9548 4162 9612
rect 4226 9548 4243 9612
rect 4307 9548 4324 9612
rect 4388 9548 4405 9612
rect 4469 9548 4486 9612
rect 4550 9548 4567 9612
rect 4631 9548 4648 9612
rect 4712 9548 4729 9612
rect 4793 9548 4809 9612
rect 4873 9548 4874 9612
rect 0 9547 4874 9548
rect 10083 9612 15000 9613
rect 10083 9548 10084 9612
rect 10148 9548 10165 9612
rect 10229 9548 10246 9612
rect 10310 9548 10327 9612
rect 10391 9548 10408 9612
rect 10472 9548 10489 9612
rect 10553 9548 10570 9612
rect 10634 9548 10651 9612
rect 10715 9548 10732 9612
rect 10796 9548 10813 9612
rect 10877 9548 10894 9612
rect 10958 9548 10975 9612
rect 11039 9548 11056 9612
rect 11120 9548 11137 9612
rect 11201 9548 11218 9612
rect 11282 9548 11299 9612
rect 11363 9548 11380 9612
rect 11444 9548 11461 9612
rect 11525 9548 11542 9612
rect 11606 9548 11623 9612
rect 11687 9548 11704 9612
rect 11768 9548 11785 9612
rect 11849 9548 11866 9612
rect 11930 9548 11947 9612
rect 12011 9548 12028 9612
rect 12092 9548 12109 9612
rect 12173 9548 12190 9612
rect 12254 9548 12271 9612
rect 12335 9548 12352 9612
rect 12416 9548 12433 9612
rect 12497 9548 12514 9612
rect 12578 9548 12595 9612
rect 12659 9548 12676 9612
rect 12740 9548 12757 9612
rect 12821 9548 12838 9612
rect 12902 9548 12919 9612
rect 12983 9548 13000 9612
rect 13064 9548 13081 9612
rect 13145 9548 13162 9612
rect 13226 9548 13243 9612
rect 13307 9548 13324 9612
rect 13388 9548 13405 9612
rect 13469 9548 13486 9612
rect 13550 9548 13567 9612
rect 13631 9548 13648 9612
rect 13712 9548 13729 9612
rect 13793 9548 13810 9612
rect 13874 9548 13891 9612
rect 13955 9548 13972 9612
rect 14036 9548 14053 9612
rect 14117 9548 14134 9612
rect 14198 9548 14215 9612
rect 14279 9548 14296 9612
rect 14360 9548 14378 9612
rect 14442 9548 14460 9612
rect 14524 9548 14542 9612
rect 14606 9548 14624 9612
rect 14688 9548 14706 9612
rect 14770 9548 14788 9612
rect 14852 9548 15000 9612
rect 10083 9547 15000 9548
rect 0 8317 254 9247
rect 14746 8317 15000 9247
rect 0 8032 4874 8037
rect 0 7968 200 8032
rect 264 7968 281 8032
rect 345 7968 362 8032
rect 426 7968 443 8032
rect 507 7968 524 8032
rect 588 7968 605 8032
rect 669 7968 686 8032
rect 750 7968 767 8032
rect 831 7968 848 8032
rect 912 7968 929 8032
rect 993 7968 1010 8032
rect 1074 7968 1091 8032
rect 1155 7968 1172 8032
rect 1236 7968 1253 8032
rect 1317 7968 1334 8032
rect 1398 7968 1415 8032
rect 1479 7968 1496 8032
rect 1560 7968 1577 8032
rect 1641 7968 1658 8032
rect 1722 7968 1739 8032
rect 1803 7968 1820 8032
rect 1884 7968 1901 8032
rect 1965 7968 1982 8032
rect 2046 7968 2063 8032
rect 2127 7968 2144 8032
rect 2208 7968 2225 8032
rect 2289 7968 2306 8032
rect 2370 7968 2387 8032
rect 2451 7968 2468 8032
rect 2532 7968 2549 8032
rect 2613 7968 2630 8032
rect 2694 7968 2711 8032
rect 2775 7968 2792 8032
rect 2856 7968 2873 8032
rect 2937 7968 2954 8032
rect 3018 7968 3035 8032
rect 3099 7968 3116 8032
rect 3180 7968 3197 8032
rect 3261 7968 3278 8032
rect 3342 7968 3359 8032
rect 3423 7968 3440 8032
rect 3504 7968 3521 8032
rect 3585 7968 3602 8032
rect 3666 7968 3683 8032
rect 3747 7968 3764 8032
rect 3828 7968 3845 8032
rect 3909 7968 3926 8032
rect 3990 7968 4007 8032
rect 4071 7968 4088 8032
rect 4152 7968 4169 8032
rect 4233 7968 4249 8032
rect 4313 7968 4329 8032
rect 4393 7968 4409 8032
rect 4473 7968 4489 8032
rect 4553 7968 4569 8032
rect 4633 7968 4649 8032
rect 4713 7968 4729 8032
rect 4793 7968 4809 8032
rect 4873 7968 4874 8032
rect 0 7944 4874 7968
rect 0 7880 200 7944
rect 264 7880 281 7944
rect 345 7880 362 7944
rect 426 7880 443 7944
rect 507 7880 524 7944
rect 588 7880 605 7944
rect 669 7880 686 7944
rect 750 7880 767 7944
rect 831 7880 848 7944
rect 912 7880 929 7944
rect 993 7880 1010 7944
rect 1074 7880 1091 7944
rect 1155 7880 1172 7944
rect 1236 7880 1253 7944
rect 1317 7880 1334 7944
rect 1398 7880 1415 7944
rect 1479 7880 1496 7944
rect 1560 7880 1577 7944
rect 1641 7880 1658 7944
rect 1722 7880 1739 7944
rect 1803 7880 1820 7944
rect 1884 7880 1901 7944
rect 1965 7880 1982 7944
rect 2046 7880 2063 7944
rect 2127 7880 2144 7944
rect 2208 7880 2225 7944
rect 2289 7880 2306 7944
rect 2370 7880 2387 7944
rect 2451 7880 2468 7944
rect 2532 7880 2549 7944
rect 2613 7880 2630 7944
rect 2694 7880 2711 7944
rect 2775 7880 2792 7944
rect 2856 7880 2873 7944
rect 2937 7880 2954 7944
rect 3018 7880 3035 7944
rect 3099 7880 3116 7944
rect 3180 7880 3197 7944
rect 3261 7880 3278 7944
rect 3342 7880 3359 7944
rect 3423 7880 3440 7944
rect 3504 7880 3521 7944
rect 3585 7880 3602 7944
rect 3666 7880 3683 7944
rect 3747 7880 3764 7944
rect 3828 7880 3845 7944
rect 3909 7880 3926 7944
rect 3990 7880 4007 7944
rect 4071 7880 4088 7944
rect 4152 7880 4169 7944
rect 4233 7880 4249 7944
rect 4313 7880 4329 7944
rect 4393 7880 4409 7944
rect 4473 7880 4489 7944
rect 4553 7880 4569 7944
rect 4633 7880 4649 7944
rect 4713 7880 4729 7944
rect 4793 7880 4809 7944
rect 4873 7880 4874 7944
rect 0 7856 4874 7880
rect 0 7792 200 7856
rect 264 7792 281 7856
rect 345 7792 362 7856
rect 426 7792 443 7856
rect 507 7792 524 7856
rect 588 7792 605 7856
rect 669 7792 686 7856
rect 750 7792 767 7856
rect 831 7792 848 7856
rect 912 7792 929 7856
rect 993 7792 1010 7856
rect 1074 7792 1091 7856
rect 1155 7792 1172 7856
rect 1236 7792 1253 7856
rect 1317 7792 1334 7856
rect 1398 7792 1415 7856
rect 1479 7792 1496 7856
rect 1560 7792 1577 7856
rect 1641 7792 1658 7856
rect 1722 7792 1739 7856
rect 1803 7792 1820 7856
rect 1884 7792 1901 7856
rect 1965 7792 1982 7856
rect 2046 7792 2063 7856
rect 2127 7792 2144 7856
rect 2208 7792 2225 7856
rect 2289 7792 2306 7856
rect 2370 7792 2387 7856
rect 2451 7792 2468 7856
rect 2532 7792 2549 7856
rect 2613 7792 2630 7856
rect 2694 7792 2711 7856
rect 2775 7792 2792 7856
rect 2856 7792 2873 7856
rect 2937 7792 2954 7856
rect 3018 7792 3035 7856
rect 3099 7792 3116 7856
rect 3180 7792 3197 7856
rect 3261 7792 3278 7856
rect 3342 7792 3359 7856
rect 3423 7792 3440 7856
rect 3504 7792 3521 7856
rect 3585 7792 3602 7856
rect 3666 7792 3683 7856
rect 3747 7792 3764 7856
rect 3828 7792 3845 7856
rect 3909 7792 3926 7856
rect 3990 7792 4007 7856
rect 4071 7792 4088 7856
rect 4152 7792 4169 7856
rect 4233 7792 4249 7856
rect 4313 7792 4329 7856
rect 4393 7792 4409 7856
rect 4473 7792 4489 7856
rect 4553 7792 4569 7856
rect 4633 7792 4649 7856
rect 4713 7792 4729 7856
rect 4793 7792 4809 7856
rect 4873 7792 4874 7856
rect 0 7768 4874 7792
rect 0 7704 200 7768
rect 264 7704 281 7768
rect 345 7704 362 7768
rect 426 7704 443 7768
rect 507 7704 524 7768
rect 588 7704 605 7768
rect 669 7704 686 7768
rect 750 7704 767 7768
rect 831 7704 848 7768
rect 912 7704 929 7768
rect 993 7704 1010 7768
rect 1074 7704 1091 7768
rect 1155 7704 1172 7768
rect 1236 7704 1253 7768
rect 1317 7704 1334 7768
rect 1398 7704 1415 7768
rect 1479 7704 1496 7768
rect 1560 7704 1577 7768
rect 1641 7704 1658 7768
rect 1722 7704 1739 7768
rect 1803 7704 1820 7768
rect 1884 7704 1901 7768
rect 1965 7704 1982 7768
rect 2046 7704 2063 7768
rect 2127 7704 2144 7768
rect 2208 7704 2225 7768
rect 2289 7704 2306 7768
rect 2370 7704 2387 7768
rect 2451 7704 2468 7768
rect 2532 7704 2549 7768
rect 2613 7704 2630 7768
rect 2694 7704 2711 7768
rect 2775 7704 2792 7768
rect 2856 7704 2873 7768
rect 2937 7704 2954 7768
rect 3018 7704 3035 7768
rect 3099 7704 3116 7768
rect 3180 7704 3197 7768
rect 3261 7704 3278 7768
rect 3342 7704 3359 7768
rect 3423 7704 3440 7768
rect 3504 7704 3521 7768
rect 3585 7704 3602 7768
rect 3666 7704 3683 7768
rect 3747 7704 3764 7768
rect 3828 7704 3845 7768
rect 3909 7704 3926 7768
rect 3990 7704 4007 7768
rect 4071 7704 4088 7768
rect 4152 7704 4169 7768
rect 4233 7704 4249 7768
rect 4313 7704 4329 7768
rect 4393 7704 4409 7768
rect 4473 7704 4489 7768
rect 4553 7704 4569 7768
rect 4633 7704 4649 7768
rect 4713 7704 4729 7768
rect 4793 7704 4809 7768
rect 4873 7704 4874 7768
rect 0 7680 4874 7704
rect 0 7616 200 7680
rect 264 7616 281 7680
rect 345 7616 362 7680
rect 426 7616 443 7680
rect 507 7616 524 7680
rect 588 7616 605 7680
rect 669 7616 686 7680
rect 750 7616 767 7680
rect 831 7616 848 7680
rect 912 7616 929 7680
rect 993 7616 1010 7680
rect 1074 7616 1091 7680
rect 1155 7616 1172 7680
rect 1236 7616 1253 7680
rect 1317 7616 1334 7680
rect 1398 7616 1415 7680
rect 1479 7616 1496 7680
rect 1560 7616 1577 7680
rect 1641 7616 1658 7680
rect 1722 7616 1739 7680
rect 1803 7616 1820 7680
rect 1884 7616 1901 7680
rect 1965 7616 1982 7680
rect 2046 7616 2063 7680
rect 2127 7616 2144 7680
rect 2208 7616 2225 7680
rect 2289 7616 2306 7680
rect 2370 7616 2387 7680
rect 2451 7616 2468 7680
rect 2532 7616 2549 7680
rect 2613 7616 2630 7680
rect 2694 7616 2711 7680
rect 2775 7616 2792 7680
rect 2856 7616 2873 7680
rect 2937 7616 2954 7680
rect 3018 7616 3035 7680
rect 3099 7616 3116 7680
rect 3180 7616 3197 7680
rect 3261 7616 3278 7680
rect 3342 7616 3359 7680
rect 3423 7616 3440 7680
rect 3504 7616 3521 7680
rect 3585 7616 3602 7680
rect 3666 7616 3683 7680
rect 3747 7616 3764 7680
rect 3828 7616 3845 7680
rect 3909 7616 3926 7680
rect 3990 7616 4007 7680
rect 4071 7616 4088 7680
rect 4152 7616 4169 7680
rect 4233 7616 4249 7680
rect 4313 7616 4329 7680
rect 4393 7616 4409 7680
rect 4473 7616 4489 7680
rect 4553 7616 4569 7680
rect 4633 7616 4649 7680
rect 4713 7616 4729 7680
rect 4793 7616 4809 7680
rect 4873 7616 4874 7680
rect 0 7592 4874 7616
rect 0 7528 200 7592
rect 264 7528 281 7592
rect 345 7528 362 7592
rect 426 7528 443 7592
rect 507 7528 524 7592
rect 588 7528 605 7592
rect 669 7528 686 7592
rect 750 7528 767 7592
rect 831 7528 848 7592
rect 912 7528 929 7592
rect 993 7528 1010 7592
rect 1074 7528 1091 7592
rect 1155 7528 1172 7592
rect 1236 7528 1253 7592
rect 1317 7528 1334 7592
rect 1398 7528 1415 7592
rect 1479 7528 1496 7592
rect 1560 7528 1577 7592
rect 1641 7528 1658 7592
rect 1722 7528 1739 7592
rect 1803 7528 1820 7592
rect 1884 7528 1901 7592
rect 1965 7528 1982 7592
rect 2046 7528 2063 7592
rect 2127 7528 2144 7592
rect 2208 7528 2225 7592
rect 2289 7528 2306 7592
rect 2370 7528 2387 7592
rect 2451 7528 2468 7592
rect 2532 7528 2549 7592
rect 2613 7528 2630 7592
rect 2694 7528 2711 7592
rect 2775 7528 2792 7592
rect 2856 7528 2873 7592
rect 2937 7528 2954 7592
rect 3018 7528 3035 7592
rect 3099 7528 3116 7592
rect 3180 7528 3197 7592
rect 3261 7528 3278 7592
rect 3342 7528 3359 7592
rect 3423 7528 3440 7592
rect 3504 7528 3521 7592
rect 3585 7528 3602 7592
rect 3666 7528 3683 7592
rect 3747 7528 3764 7592
rect 3828 7528 3845 7592
rect 3909 7528 3926 7592
rect 3990 7528 4007 7592
rect 4071 7528 4088 7592
rect 4152 7528 4169 7592
rect 4233 7528 4249 7592
rect 4313 7528 4329 7592
rect 4393 7528 4409 7592
rect 4473 7528 4489 7592
rect 4553 7528 4569 7592
rect 4633 7528 4649 7592
rect 4713 7528 4729 7592
rect 4793 7528 4809 7592
rect 4873 7528 4874 7592
rect 0 7504 4874 7528
rect 0 7440 200 7504
rect 264 7440 281 7504
rect 345 7440 362 7504
rect 426 7440 443 7504
rect 507 7440 524 7504
rect 588 7440 605 7504
rect 669 7440 686 7504
rect 750 7440 767 7504
rect 831 7440 848 7504
rect 912 7440 929 7504
rect 993 7440 1010 7504
rect 1074 7440 1091 7504
rect 1155 7440 1172 7504
rect 1236 7440 1253 7504
rect 1317 7440 1334 7504
rect 1398 7440 1415 7504
rect 1479 7440 1496 7504
rect 1560 7440 1577 7504
rect 1641 7440 1658 7504
rect 1722 7440 1739 7504
rect 1803 7440 1820 7504
rect 1884 7440 1901 7504
rect 1965 7440 1982 7504
rect 2046 7440 2063 7504
rect 2127 7440 2144 7504
rect 2208 7440 2225 7504
rect 2289 7440 2306 7504
rect 2370 7440 2387 7504
rect 2451 7440 2468 7504
rect 2532 7440 2549 7504
rect 2613 7440 2630 7504
rect 2694 7440 2711 7504
rect 2775 7440 2792 7504
rect 2856 7440 2873 7504
rect 2937 7440 2954 7504
rect 3018 7440 3035 7504
rect 3099 7440 3116 7504
rect 3180 7440 3197 7504
rect 3261 7440 3278 7504
rect 3342 7440 3359 7504
rect 3423 7440 3440 7504
rect 3504 7440 3521 7504
rect 3585 7440 3602 7504
rect 3666 7440 3683 7504
rect 3747 7440 3764 7504
rect 3828 7440 3845 7504
rect 3909 7440 3926 7504
rect 3990 7440 4007 7504
rect 4071 7440 4088 7504
rect 4152 7440 4169 7504
rect 4233 7440 4249 7504
rect 4313 7440 4329 7504
rect 4393 7440 4409 7504
rect 4473 7440 4489 7504
rect 4553 7440 4569 7504
rect 4633 7440 4649 7504
rect 4713 7440 4729 7504
rect 4793 7440 4809 7504
rect 4873 7440 4874 7504
rect 0 7416 4874 7440
rect 0 7352 200 7416
rect 264 7352 281 7416
rect 345 7352 362 7416
rect 426 7352 443 7416
rect 507 7352 524 7416
rect 588 7352 605 7416
rect 669 7352 686 7416
rect 750 7352 767 7416
rect 831 7352 848 7416
rect 912 7352 929 7416
rect 993 7352 1010 7416
rect 1074 7352 1091 7416
rect 1155 7352 1172 7416
rect 1236 7352 1253 7416
rect 1317 7352 1334 7416
rect 1398 7352 1415 7416
rect 1479 7352 1496 7416
rect 1560 7352 1577 7416
rect 1641 7352 1658 7416
rect 1722 7352 1739 7416
rect 1803 7352 1820 7416
rect 1884 7352 1901 7416
rect 1965 7352 1982 7416
rect 2046 7352 2063 7416
rect 2127 7352 2144 7416
rect 2208 7352 2225 7416
rect 2289 7352 2306 7416
rect 2370 7352 2387 7416
rect 2451 7352 2468 7416
rect 2532 7352 2549 7416
rect 2613 7352 2630 7416
rect 2694 7352 2711 7416
rect 2775 7352 2792 7416
rect 2856 7352 2873 7416
rect 2937 7352 2954 7416
rect 3018 7352 3035 7416
rect 3099 7352 3116 7416
rect 3180 7352 3197 7416
rect 3261 7352 3278 7416
rect 3342 7352 3359 7416
rect 3423 7352 3440 7416
rect 3504 7352 3521 7416
rect 3585 7352 3602 7416
rect 3666 7352 3683 7416
rect 3747 7352 3764 7416
rect 3828 7352 3845 7416
rect 3909 7352 3926 7416
rect 3990 7352 4007 7416
rect 4071 7352 4088 7416
rect 4152 7352 4169 7416
rect 4233 7352 4249 7416
rect 4313 7352 4329 7416
rect 4393 7352 4409 7416
rect 4473 7352 4489 7416
rect 4553 7352 4569 7416
rect 4633 7352 4649 7416
rect 4713 7352 4729 7416
rect 4793 7352 4809 7416
rect 4873 7352 4874 7416
rect 0 7347 4874 7352
rect 10083 8032 15000 8037
rect 10083 7968 10084 8032
rect 10148 7968 10166 8032
rect 10230 7968 10248 8032
rect 10312 7968 10330 8032
rect 10394 7968 10412 8032
rect 10476 7968 10494 8032
rect 10558 7968 10576 8032
rect 10640 7968 10657 8032
rect 10721 7968 10738 8032
rect 10802 7968 10819 8032
rect 10883 7968 10900 8032
rect 10964 7968 10981 8032
rect 11045 7968 11062 8032
rect 11126 7968 11143 8032
rect 11207 7968 11224 8032
rect 11288 7968 11305 8032
rect 11369 7968 11386 8032
rect 11450 7968 11467 8032
rect 11531 7968 11548 8032
rect 11612 7968 11629 8032
rect 11693 7968 11710 8032
rect 11774 7968 11791 8032
rect 11855 7968 11872 8032
rect 11936 7968 11953 8032
rect 12017 7968 12034 8032
rect 12098 7968 12115 8032
rect 12179 7968 12196 8032
rect 12260 7968 12277 8032
rect 12341 7968 12358 8032
rect 12422 7968 12439 8032
rect 12503 7968 12520 8032
rect 12584 7968 12601 8032
rect 12665 7968 12682 8032
rect 12746 7968 12763 8032
rect 12827 7968 12844 8032
rect 12908 7968 12925 8032
rect 12989 7968 13006 8032
rect 13070 7968 13087 8032
rect 13151 7968 13168 8032
rect 13232 7968 13249 8032
rect 13313 7968 13330 8032
rect 13394 7968 13411 8032
rect 13475 7968 13492 8032
rect 13556 7968 13573 8032
rect 13637 7968 13654 8032
rect 13718 7968 13735 8032
rect 13799 7968 13816 8032
rect 13880 7968 13897 8032
rect 13961 7968 13978 8032
rect 14042 7968 14059 8032
rect 14123 7968 14140 8032
rect 14204 7968 14221 8032
rect 14285 7968 14302 8032
rect 14366 7968 14383 8032
rect 14447 7968 14464 8032
rect 14528 7968 14545 8032
rect 14609 7968 14626 8032
rect 14690 7968 14707 8032
rect 14771 7968 14788 8032
rect 14852 7968 15000 8032
rect 10083 7944 15000 7968
rect 10083 7880 10084 7944
rect 10148 7880 10166 7944
rect 10230 7880 10248 7944
rect 10312 7880 10330 7944
rect 10394 7880 10412 7944
rect 10476 7880 10494 7944
rect 10558 7880 10576 7944
rect 10640 7880 10657 7944
rect 10721 7880 10738 7944
rect 10802 7880 10819 7944
rect 10883 7880 10900 7944
rect 10964 7880 10981 7944
rect 11045 7880 11062 7944
rect 11126 7880 11143 7944
rect 11207 7880 11224 7944
rect 11288 7880 11305 7944
rect 11369 7880 11386 7944
rect 11450 7880 11467 7944
rect 11531 7880 11548 7944
rect 11612 7880 11629 7944
rect 11693 7880 11710 7944
rect 11774 7880 11791 7944
rect 11855 7880 11872 7944
rect 11936 7880 11953 7944
rect 12017 7880 12034 7944
rect 12098 7880 12115 7944
rect 12179 7880 12196 7944
rect 12260 7880 12277 7944
rect 12341 7880 12358 7944
rect 12422 7880 12439 7944
rect 12503 7880 12520 7944
rect 12584 7880 12601 7944
rect 12665 7880 12682 7944
rect 12746 7880 12763 7944
rect 12827 7880 12844 7944
rect 12908 7880 12925 7944
rect 12989 7880 13006 7944
rect 13070 7880 13087 7944
rect 13151 7880 13168 7944
rect 13232 7880 13249 7944
rect 13313 7880 13330 7944
rect 13394 7880 13411 7944
rect 13475 7880 13492 7944
rect 13556 7880 13573 7944
rect 13637 7880 13654 7944
rect 13718 7880 13735 7944
rect 13799 7880 13816 7944
rect 13880 7880 13897 7944
rect 13961 7880 13978 7944
rect 14042 7880 14059 7944
rect 14123 7880 14140 7944
rect 14204 7880 14221 7944
rect 14285 7880 14302 7944
rect 14366 7880 14383 7944
rect 14447 7880 14464 7944
rect 14528 7880 14545 7944
rect 14609 7880 14626 7944
rect 14690 7880 14707 7944
rect 14771 7880 14788 7944
rect 14852 7880 15000 7944
rect 10083 7856 15000 7880
rect 10083 7792 10084 7856
rect 10148 7792 10166 7856
rect 10230 7792 10248 7856
rect 10312 7792 10330 7856
rect 10394 7792 10412 7856
rect 10476 7792 10494 7856
rect 10558 7792 10576 7856
rect 10640 7792 10657 7856
rect 10721 7792 10738 7856
rect 10802 7792 10819 7856
rect 10883 7792 10900 7856
rect 10964 7792 10981 7856
rect 11045 7792 11062 7856
rect 11126 7792 11143 7856
rect 11207 7792 11224 7856
rect 11288 7792 11305 7856
rect 11369 7792 11386 7856
rect 11450 7792 11467 7856
rect 11531 7792 11548 7856
rect 11612 7792 11629 7856
rect 11693 7792 11710 7856
rect 11774 7792 11791 7856
rect 11855 7792 11872 7856
rect 11936 7792 11953 7856
rect 12017 7792 12034 7856
rect 12098 7792 12115 7856
rect 12179 7792 12196 7856
rect 12260 7792 12277 7856
rect 12341 7792 12358 7856
rect 12422 7792 12439 7856
rect 12503 7792 12520 7856
rect 12584 7792 12601 7856
rect 12665 7792 12682 7856
rect 12746 7792 12763 7856
rect 12827 7792 12844 7856
rect 12908 7792 12925 7856
rect 12989 7792 13006 7856
rect 13070 7792 13087 7856
rect 13151 7792 13168 7856
rect 13232 7792 13249 7856
rect 13313 7792 13330 7856
rect 13394 7792 13411 7856
rect 13475 7792 13492 7856
rect 13556 7792 13573 7856
rect 13637 7792 13654 7856
rect 13718 7792 13735 7856
rect 13799 7792 13816 7856
rect 13880 7792 13897 7856
rect 13961 7792 13978 7856
rect 14042 7792 14059 7856
rect 14123 7792 14140 7856
rect 14204 7792 14221 7856
rect 14285 7792 14302 7856
rect 14366 7792 14383 7856
rect 14447 7792 14464 7856
rect 14528 7792 14545 7856
rect 14609 7792 14626 7856
rect 14690 7792 14707 7856
rect 14771 7792 14788 7856
rect 14852 7792 15000 7856
rect 10083 7768 15000 7792
rect 10083 7704 10084 7768
rect 10148 7704 10166 7768
rect 10230 7704 10248 7768
rect 10312 7704 10330 7768
rect 10394 7704 10412 7768
rect 10476 7704 10494 7768
rect 10558 7704 10576 7768
rect 10640 7704 10657 7768
rect 10721 7704 10738 7768
rect 10802 7704 10819 7768
rect 10883 7704 10900 7768
rect 10964 7704 10981 7768
rect 11045 7704 11062 7768
rect 11126 7704 11143 7768
rect 11207 7704 11224 7768
rect 11288 7704 11305 7768
rect 11369 7704 11386 7768
rect 11450 7704 11467 7768
rect 11531 7704 11548 7768
rect 11612 7704 11629 7768
rect 11693 7704 11710 7768
rect 11774 7704 11791 7768
rect 11855 7704 11872 7768
rect 11936 7704 11953 7768
rect 12017 7704 12034 7768
rect 12098 7704 12115 7768
rect 12179 7704 12196 7768
rect 12260 7704 12277 7768
rect 12341 7704 12358 7768
rect 12422 7704 12439 7768
rect 12503 7704 12520 7768
rect 12584 7704 12601 7768
rect 12665 7704 12682 7768
rect 12746 7704 12763 7768
rect 12827 7704 12844 7768
rect 12908 7704 12925 7768
rect 12989 7704 13006 7768
rect 13070 7704 13087 7768
rect 13151 7704 13168 7768
rect 13232 7704 13249 7768
rect 13313 7704 13330 7768
rect 13394 7704 13411 7768
rect 13475 7704 13492 7768
rect 13556 7704 13573 7768
rect 13637 7704 13654 7768
rect 13718 7704 13735 7768
rect 13799 7704 13816 7768
rect 13880 7704 13897 7768
rect 13961 7704 13978 7768
rect 14042 7704 14059 7768
rect 14123 7704 14140 7768
rect 14204 7704 14221 7768
rect 14285 7704 14302 7768
rect 14366 7704 14383 7768
rect 14447 7704 14464 7768
rect 14528 7704 14545 7768
rect 14609 7704 14626 7768
rect 14690 7704 14707 7768
rect 14771 7704 14788 7768
rect 14852 7704 15000 7768
rect 10083 7680 15000 7704
rect 10083 7616 10084 7680
rect 10148 7616 10166 7680
rect 10230 7616 10248 7680
rect 10312 7616 10330 7680
rect 10394 7616 10412 7680
rect 10476 7616 10494 7680
rect 10558 7616 10576 7680
rect 10640 7616 10657 7680
rect 10721 7616 10738 7680
rect 10802 7616 10819 7680
rect 10883 7616 10900 7680
rect 10964 7616 10981 7680
rect 11045 7616 11062 7680
rect 11126 7616 11143 7680
rect 11207 7616 11224 7680
rect 11288 7616 11305 7680
rect 11369 7616 11386 7680
rect 11450 7616 11467 7680
rect 11531 7616 11548 7680
rect 11612 7616 11629 7680
rect 11693 7616 11710 7680
rect 11774 7616 11791 7680
rect 11855 7616 11872 7680
rect 11936 7616 11953 7680
rect 12017 7616 12034 7680
rect 12098 7616 12115 7680
rect 12179 7616 12196 7680
rect 12260 7616 12277 7680
rect 12341 7616 12358 7680
rect 12422 7616 12439 7680
rect 12503 7616 12520 7680
rect 12584 7616 12601 7680
rect 12665 7616 12682 7680
rect 12746 7616 12763 7680
rect 12827 7616 12844 7680
rect 12908 7616 12925 7680
rect 12989 7616 13006 7680
rect 13070 7616 13087 7680
rect 13151 7616 13168 7680
rect 13232 7616 13249 7680
rect 13313 7616 13330 7680
rect 13394 7616 13411 7680
rect 13475 7616 13492 7680
rect 13556 7616 13573 7680
rect 13637 7616 13654 7680
rect 13718 7616 13735 7680
rect 13799 7616 13816 7680
rect 13880 7616 13897 7680
rect 13961 7616 13978 7680
rect 14042 7616 14059 7680
rect 14123 7616 14140 7680
rect 14204 7616 14221 7680
rect 14285 7616 14302 7680
rect 14366 7616 14383 7680
rect 14447 7616 14464 7680
rect 14528 7616 14545 7680
rect 14609 7616 14626 7680
rect 14690 7616 14707 7680
rect 14771 7616 14788 7680
rect 14852 7616 15000 7680
rect 10083 7592 15000 7616
rect 10083 7528 10084 7592
rect 10148 7528 10166 7592
rect 10230 7528 10248 7592
rect 10312 7528 10330 7592
rect 10394 7528 10412 7592
rect 10476 7528 10494 7592
rect 10558 7528 10576 7592
rect 10640 7528 10657 7592
rect 10721 7528 10738 7592
rect 10802 7528 10819 7592
rect 10883 7528 10900 7592
rect 10964 7528 10981 7592
rect 11045 7528 11062 7592
rect 11126 7528 11143 7592
rect 11207 7528 11224 7592
rect 11288 7528 11305 7592
rect 11369 7528 11386 7592
rect 11450 7528 11467 7592
rect 11531 7528 11548 7592
rect 11612 7528 11629 7592
rect 11693 7528 11710 7592
rect 11774 7528 11791 7592
rect 11855 7528 11872 7592
rect 11936 7528 11953 7592
rect 12017 7528 12034 7592
rect 12098 7528 12115 7592
rect 12179 7528 12196 7592
rect 12260 7528 12277 7592
rect 12341 7528 12358 7592
rect 12422 7528 12439 7592
rect 12503 7528 12520 7592
rect 12584 7528 12601 7592
rect 12665 7528 12682 7592
rect 12746 7528 12763 7592
rect 12827 7528 12844 7592
rect 12908 7528 12925 7592
rect 12989 7528 13006 7592
rect 13070 7528 13087 7592
rect 13151 7528 13168 7592
rect 13232 7528 13249 7592
rect 13313 7528 13330 7592
rect 13394 7528 13411 7592
rect 13475 7528 13492 7592
rect 13556 7528 13573 7592
rect 13637 7528 13654 7592
rect 13718 7528 13735 7592
rect 13799 7528 13816 7592
rect 13880 7528 13897 7592
rect 13961 7528 13978 7592
rect 14042 7528 14059 7592
rect 14123 7528 14140 7592
rect 14204 7528 14221 7592
rect 14285 7528 14302 7592
rect 14366 7528 14383 7592
rect 14447 7528 14464 7592
rect 14528 7528 14545 7592
rect 14609 7528 14626 7592
rect 14690 7528 14707 7592
rect 14771 7528 14788 7592
rect 14852 7528 15000 7592
rect 10083 7504 15000 7528
rect 10083 7440 10084 7504
rect 10148 7440 10166 7504
rect 10230 7440 10248 7504
rect 10312 7440 10330 7504
rect 10394 7440 10412 7504
rect 10476 7440 10494 7504
rect 10558 7440 10576 7504
rect 10640 7440 10657 7504
rect 10721 7440 10738 7504
rect 10802 7440 10819 7504
rect 10883 7440 10900 7504
rect 10964 7440 10981 7504
rect 11045 7440 11062 7504
rect 11126 7440 11143 7504
rect 11207 7440 11224 7504
rect 11288 7440 11305 7504
rect 11369 7440 11386 7504
rect 11450 7440 11467 7504
rect 11531 7440 11548 7504
rect 11612 7440 11629 7504
rect 11693 7440 11710 7504
rect 11774 7440 11791 7504
rect 11855 7440 11872 7504
rect 11936 7440 11953 7504
rect 12017 7440 12034 7504
rect 12098 7440 12115 7504
rect 12179 7440 12196 7504
rect 12260 7440 12277 7504
rect 12341 7440 12358 7504
rect 12422 7440 12439 7504
rect 12503 7440 12520 7504
rect 12584 7440 12601 7504
rect 12665 7440 12682 7504
rect 12746 7440 12763 7504
rect 12827 7440 12844 7504
rect 12908 7440 12925 7504
rect 12989 7440 13006 7504
rect 13070 7440 13087 7504
rect 13151 7440 13168 7504
rect 13232 7440 13249 7504
rect 13313 7440 13330 7504
rect 13394 7440 13411 7504
rect 13475 7440 13492 7504
rect 13556 7440 13573 7504
rect 13637 7440 13654 7504
rect 13718 7440 13735 7504
rect 13799 7440 13816 7504
rect 13880 7440 13897 7504
rect 13961 7440 13978 7504
rect 14042 7440 14059 7504
rect 14123 7440 14140 7504
rect 14204 7440 14221 7504
rect 14285 7440 14302 7504
rect 14366 7440 14383 7504
rect 14447 7440 14464 7504
rect 14528 7440 14545 7504
rect 14609 7440 14626 7504
rect 14690 7440 14707 7504
rect 14771 7440 14788 7504
rect 14852 7440 15000 7504
rect 10083 7416 15000 7440
rect 10083 7352 10084 7416
rect 10148 7352 10166 7416
rect 10230 7352 10248 7416
rect 10312 7352 10330 7416
rect 10394 7352 10412 7416
rect 10476 7352 10494 7416
rect 10558 7352 10576 7416
rect 10640 7352 10657 7416
rect 10721 7352 10738 7416
rect 10802 7352 10819 7416
rect 10883 7352 10900 7416
rect 10964 7352 10981 7416
rect 11045 7352 11062 7416
rect 11126 7352 11143 7416
rect 11207 7352 11224 7416
rect 11288 7352 11305 7416
rect 11369 7352 11386 7416
rect 11450 7352 11467 7416
rect 11531 7352 11548 7416
rect 11612 7352 11629 7416
rect 11693 7352 11710 7416
rect 11774 7352 11791 7416
rect 11855 7352 11872 7416
rect 11936 7352 11953 7416
rect 12017 7352 12034 7416
rect 12098 7352 12115 7416
rect 12179 7352 12196 7416
rect 12260 7352 12277 7416
rect 12341 7352 12358 7416
rect 12422 7352 12439 7416
rect 12503 7352 12520 7416
rect 12584 7352 12601 7416
rect 12665 7352 12682 7416
rect 12746 7352 12763 7416
rect 12827 7352 12844 7416
rect 12908 7352 12925 7416
rect 12989 7352 13006 7416
rect 13070 7352 13087 7416
rect 13151 7352 13168 7416
rect 13232 7352 13249 7416
rect 13313 7352 13330 7416
rect 13394 7352 13411 7416
rect 13475 7352 13492 7416
rect 13556 7352 13573 7416
rect 13637 7352 13654 7416
rect 13718 7352 13735 7416
rect 13799 7352 13816 7416
rect 13880 7352 13897 7416
rect 13961 7352 13978 7416
rect 14042 7352 14059 7416
rect 14123 7352 14140 7416
rect 14204 7352 14221 7416
rect 14285 7352 14302 7416
rect 14366 7352 14383 7416
rect 14447 7352 14464 7416
rect 14528 7352 14545 7416
rect 14609 7352 14626 7416
rect 14690 7352 14707 7416
rect 14771 7352 14788 7416
rect 14852 7352 15000 7416
rect 10083 7347 15000 7352
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 5167 254 6097
rect 14746 5167 15000 6097
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 2987 193 3677
rect 14807 2987 15000 3677
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 18997
rect 14746 14007 15000 18997
rect 0 12837 254 13687
rect 14746 12837 15000 13687
rect 0 11667 254 12517
rect 14746 11667 15000 12517
rect 0 9547 254 11347
rect 14746 9547 15000 11347
rect 0 8337 254 9227
rect 14746 8337 15000 9227
rect 0 7368 254 8017
rect 14746 7368 15000 8017
rect 0 6397 254 7047
rect 14746 6397 15000 7047
rect 0 5187 254 6077
rect 14746 5187 15000 6077
rect 0 3977 254 4867
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 14746 1797 15000 2687
rect 0 427 254 1477
rect 14746 427 15000 1477
use sky130_fd_io__com_bus_hookup  sky130_fd_io__com_bus_hookup_0
timestamp 1619729480
transform 1 0 0 0 1 549
box 0 -142 15000 39451
<< labels >>
flabel metal5 s 0 3007 193 3657 3 FreeSans 520 0 0 0 VDDA
port 12 nsew power bidirectional
flabel metal5 s 14746 14007 15000 18997 3 FreeSans 520 180 0 0 VDDIO
port 16 nsew power bidirectional
flabel metal5 s 14746 3977 15000 4867 3 FreeSans 520 180 0 0 VDDIO
port 17 nsew power bidirectional
flabel metal5 s 0 427 254 1477 3 FreeSans 520 0 0 0 VCCHIB
port 8 nsew power bidirectional
flabel metal5 s 0 14007 254 18997 3 FreeSans 520 0 0 0 VDDIO
port 18 nsew power bidirectional
flabel metal5 s 0 3977 254 4867 3 FreeSans 520 0 0 0 VDDIO
port 19 nsew power bidirectional
flabel metal5 s 14746 12837 15000 13687 3 FreeSans 520 180 0 0 VDDIO_Q
port 24 nsew power bidirectional
flabel metal5 s 0 12837 254 13687 3 FreeSans 520 0 0 0 VDDIO_Q
port 25 nsew power bidirectional
flabel metal5 s 14746 35157 15000 40000 3 FreeSans 520 180 0 0 VSSIO
port 44 nsew ground bidirectional
flabel metal5 s 14746 5187 15000 6077 3 FreeSans 520 180 0 0 VSSIO
port 45 nsew ground bidirectional
flabel metal5 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 46 nsew ground bidirectional
flabel metal5 s 0 5187 254 6077 3 FreeSans 520 0 0 0 VSSIO
port 47 nsew ground bidirectional
flabel metal5 s 14746 11667 15000 12517 3 FreeSans 520 180 0 0 VSSIO_Q
port 52 nsew ground bidirectional
flabel metal5 s 0 11667 254 12517 3 FreeSans 520 0 0 0 VSSIO_Q
port 53 nsew ground bidirectional
flabel metal5 s 14746 6397 15000 7047 3 FreeSans 520 180 0 0 VSWITCH
port 56 nsew power bidirectional
flabel metal5 s 14746 1797 15000 2687 3 FreeSans 520 180 0 0 VCCD
port 4 nsew power bidirectional
flabel metal5 s 0 1797 254 2687 3 FreeSans 520 0 0 0 VCCD
port 5 nsew power bidirectional
flabel metal5 s 14746 427 15000 1477 3 FreeSans 520 180 0 0 VCCHIB
port 9 nsew power bidirectional
flabel metal5 s 14807 3007 15000 3657 3 FreeSans 520 180 0 0 VDDA
port 13 nsew power bidirectional
flabel metal5 s 14746 9547 15000 11347 3 FreeSans 520 180 0 0 VSSA
port 28 nsew ground bidirectional
flabel metal5 s 14746 7368 15000 8017 3 FreeSans 520 180 0 0 VSSA
port 29 nsew ground bidirectional
flabel metal5 s 0 9547 254 11347 3 FreeSans 520 0 0 0 VSSA
port 30 nsew ground bidirectional
flabel metal5 s 0 7368 254 8017 3 FreeSans 520 0 0 0 VSSA
port 31 nsew ground bidirectional
flabel metal5 s 14746 8337 15000 9227 3 FreeSans 520 180 0 0 VSSD
port 40 nsew ground bidirectional
flabel metal5 s 0 8337 254 9227 3 FreeSans 520 0 0 0 VSSD
port 41 nsew ground bidirectional
flabel metal5 s 0 6397 254 7047 3 FreeSans 520 0 0 0 VSWITCH
port 57 nsew power bidirectional
flabel metal4 s 14746 10625 15000 11221 3 FreeSans 520 180 0 0 AMUXBUS_A
port 0 nsew signal bidirectional
flabel metal4 s 0 1777 254 2707 3 FreeSans 520 0 0 0 VCCD
port 6 nsew power bidirectional
flabel metal4 s 14746 3957 15000 4887 3 FreeSans 520 180 0 0 VDDIO
port 20 nsew power bidirectional
flabel metal4 s 14746 14007 15000 19000 3 FreeSans 520 180 0 0 VDDIO
port 21 nsew power bidirectional
flabel metal4 s 0 3957 254 4887 3 FreeSans 520 0 0 0 VDDIO
port 22 nsew power bidirectional
flabel metal4 s 0 14007 254 19000 3 FreeSans 520 0 0 0 VDDIO
port 23 nsew power bidirectional
flabel metal4 s 14807 2987 15000 3677 3 FreeSans 520 180 0 0 VDDA
port 14 nsew power bidirectional
flabel metal4 s 14746 12817 15000 13707 3 FreeSans 520 180 0 0 VDDIO_Q
port 26 nsew power bidirectional
flabel metal4 s 0 12817 254 13707 3 FreeSans 520 0 0 0 VDDIO_Q
port 27 nsew power bidirectional
flabel metal4 s 14746 7347 15000 8037 3 FreeSans 520 180 0 0 VSSA
port 32 nsew ground bidirectional
flabel metal4 s 14746 35157 15000 40000 3 FreeSans 520 180 0 0 VSSIO
port 48 nsew ground bidirectional
flabel metal4 s 14746 5167 15000 6097 3 FreeSans 520 180 0 0 VSSIO
port 49 nsew ground bidirectional
flabel metal4 s 0 35157 254 40000 3 FreeSans 520 0 0 0 VSSIO
port 50 nsew ground bidirectional
flabel metal4 s 0 5167 254 6097 3 FreeSans 520 0 0 0 VSSIO
port 51 nsew ground bidirectional
flabel metal4 s 14746 11647 15000 12537 3 FreeSans 520 180 0 0 VSSIO_Q
port 54 nsew ground bidirectional
flabel metal4 s 0 11647 254 12537 3 FreeSans 520 0 0 0 VSSIO_Q
port 55 nsew ground bidirectional
flabel metal4 s 14746 6377 15000 7067 3 FreeSans 520 180 0 0 VSWITCH
port 58 nsew power bidirectional
flabel metal4 s 0 6377 254 7067 3 FreeSans 520 0 0 0 VSWITCH
port 59 nsew power bidirectional
flabel metal4 s 0 10625 254 11221 3 FreeSans 520 0 0 0 AMUXBUS_A
port 1 nsew signal bidirectional
flabel metal4 s 14746 9673 15000 10269 3 FreeSans 520 180 0 0 AMUXBUS_B
port 2 nsew signal bidirectional
flabel metal4 s 0 9673 254 10269 3 FreeSans 520 0 0 0 AMUXBUS_B
port 3 nsew signal bidirectional
flabel metal4 s 14746 1777 15000 2707 3 FreeSans 520 180 0 0 VCCD
port 7 nsew power bidirectional
flabel metal4 s 14746 407 15000 1497 3 FreeSans 520 180 0 0 VCCHIB
port 10 nsew power bidirectional
flabel metal4 s 0 407 254 1497 3 FreeSans 520 0 0 0 VCCHIB
port 11 nsew power bidirectional
flabel metal4 s 0 9547 254 9613 3 FreeSans 520 0 0 0 VSSA
port 33 nsew ground bidirectional
flabel metal4 s 0 10329 254 10565 3 FreeSans 520 0 0 0 VSSA
port 34 nsew ground bidirectional
flabel metal4 s 0 11281 254 11347 3 FreeSans 520 0 0 0 VSSA
port 35 nsew ground bidirectional
flabel metal4 s 0 7347 254 8037 3 FreeSans 520 0 0 0 VSSA
port 36 nsew ground bidirectional
flabel metal4 s 14746 8317 15000 9247 3 FreeSans 520 180 0 0 VSSD
port 42 nsew ground bidirectional
flabel metal4 s 0 8317 254 9247 3 FreeSans 520 0 0 0 VSSD
port 43 nsew ground bidirectional
flabel metal4 s 14746 9547 15000 9613 3 FreeSans 520 180 0 0 VSSA
port 37 nsew ground bidirectional
flabel metal4 s 14746 11281 15000 11347 3 FreeSans 520 180 0 0 VSSA
port 38 nsew ground bidirectional
flabel metal4 s 14746 10329 15000 10565 3 FreeSans 520 180 0 0 VSSA
port 39 nsew ground bidirectional
flabel metal4 s 0 2987 193 3677 3 FreeSans 520 0 0 0 VDDA
port 15 nsew power bidirectional
rlabel metal4 s 105 10415 169 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 105 10415 169 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 105 10499 169 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 105 10499 169 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 112 9548 176 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 112 9548 176 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 112 11282 176 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 112 11282 176 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 187 10331 251 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 187 10331 251 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 187 10415 251 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 187 10415 251 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 187 10499 251 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 187 10499 251 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 193 9548 257 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 193 9548 257 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 193 11282 257 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 193 11282 257 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 200 7352 264 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 200 7352 264 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 200 7440 264 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 200 7440 264 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 200 7528 264 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 200 7528 264 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 200 7616 264 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 200 7616 264 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 200 7704 264 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 200 7704 264 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 200 7792 264 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 200 7792 264 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 200 7880 264 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 200 7880 264 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 200 7968 264 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 200 7968 264 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 269 10331 333 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 269 10331 333 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 269 10415 333 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 269 10415 333 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 269 10499 333 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 269 10499 333 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 274 9548 338 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 274 9548 338 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 274 11282 338 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 274 11282 338 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 281 7352 345 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 281 7352 345 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 281 7440 345 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 281 7440 345 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 281 7528 345 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 281 7528 345 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 281 7616 345 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 281 7616 345 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 281 7704 345 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 281 7704 345 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 281 7792 345 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 281 7792 345 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 281 7880 345 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 281 7880 345 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 281 7968 345 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 281 7968 345 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 351 10331 415 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 351 10331 415 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 351 10415 415 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 351 10415 415 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 351 10499 415 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 351 10499 415 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 355 9548 419 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 355 9548 419 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 355 11282 419 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 355 11282 419 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 362 7352 426 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 362 7352 426 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 362 7440 426 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 362 7440 426 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 362 7528 426 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 362 7528 426 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 362 7616 426 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 362 7616 426 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 362 7704 426 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 362 7704 426 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 362 7792 426 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 362 7792 426 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 362 7880 426 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 362 7880 426 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 362 7968 426 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 362 7968 426 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2055 10331 2119 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2055 10331 2119 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2055 10415 2119 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2055 10415 2119 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2055 10499 2119 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2055 10499 2119 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2056 9548 2120 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2056 9548 2120 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2056 11282 2120 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2056 11282 2120 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2063 7352 2127 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2063 7352 2127 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2063 7440 2127 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2063 7440 2127 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2063 7528 2127 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2063 7528 2127 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2063 7616 2127 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2063 7616 2127 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2063 7704 2127 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2063 7704 2127 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2063 7792 2127 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2063 7792 2127 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2063 7880 2127 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2063 7880 2127 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2063 7968 2127 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2063 7968 2127 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2136 10331 2200 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2136 10331 2200 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2136 10415 2200 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2136 10415 2200 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2136 10499 2200 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2136 10499 2200 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2137 9548 2201 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2137 9548 2201 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2137 11282 2201 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2137 11282 2201 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2144 7352 2208 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2144 7352 2208 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2144 7440 2208 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2144 7440 2208 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2144 7528 2208 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2144 7528 2208 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2144 7616 2208 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2144 7616 2208 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2144 7704 2208 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2144 7704 2208 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2144 7792 2208 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2144 7792 2208 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2144 7880 2208 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2144 7880 2208 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2144 7968 2208 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2144 7968 2208 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2217 10331 2281 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2217 10331 2281 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2217 10415 2281 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2217 10415 2281 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2217 10499 2281 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2217 10499 2281 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2218 9548 2282 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2218 9548 2282 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2218 11282 2282 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2218 11282 2282 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2225 7352 2289 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2225 7352 2289 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2225 7440 2289 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2225 7440 2289 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2225 7528 2289 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2225 7528 2289 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2225 7616 2289 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2225 7616 2289 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2225 7704 2289 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2225 7704 2289 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2225 7792 2289 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2225 7792 2289 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2225 7880 2289 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2225 7880 2289 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2225 7968 2289 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2225 7968 2289 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2298 10331 2362 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2298 10331 2362 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2298 10415 2362 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2298 10415 2362 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2298 10499 2362 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2298 10499 2362 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2299 9548 2363 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2299 9548 2363 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2299 11282 2363 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2299 11282 2363 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2306 7352 2370 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2306 7352 2370 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2306 7440 2370 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2306 7440 2370 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2306 7528 2370 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2306 7528 2370 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2306 7616 2370 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2306 7616 2370 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2306 7704 2370 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2306 7704 2370 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2306 7792 2370 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2306 7792 2370 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2306 7880 2370 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2306 7880 2370 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2306 7968 2370 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2306 7968 2370 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2379 10331 2443 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2379 10331 2443 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2379 10415 2443 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2379 10415 2443 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2379 10499 2443 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2379 10499 2443 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2380 9548 2444 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2380 9548 2444 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2380 11282 2444 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2380 11282 2444 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2387 7352 2451 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2387 7352 2451 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2387 7440 2451 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2387 7440 2451 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2387 7528 2451 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2387 7528 2451 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2387 7616 2451 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2387 7616 2451 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2387 7704 2451 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2387 7704 2451 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2387 7792 2451 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2387 7792 2451 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2387 7880 2451 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2387 7880 2451 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2387 7968 2451 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2387 7968 2451 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2460 10331 2524 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2460 10331 2524 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2460 10415 2524 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2460 10415 2524 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2460 10499 2524 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2460 10499 2524 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2461 9548 2525 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2461 9548 2525 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2461 11282 2525 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2461 11282 2525 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2468 7352 2532 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2468 7352 2532 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2468 7440 2532 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2468 7440 2532 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2468 7528 2532 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2468 7528 2532 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2468 7616 2532 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2468 7616 2532 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2468 7704 2532 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2468 7704 2532 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2468 7792 2532 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2468 7792 2532 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2468 7880 2532 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2468 7880 2532 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2468 7968 2532 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2468 7968 2532 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2541 10331 2605 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2541 10331 2605 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2541 10415 2605 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2541 10415 2605 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2541 10499 2605 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2541 10499 2605 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2542 9548 2606 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2542 9548 2606 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2542 11282 2606 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2542 11282 2606 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2549 7352 2613 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2549 7352 2613 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2549 7440 2613 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2549 7440 2613 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2549 7528 2613 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2549 7528 2613 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2549 7616 2613 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2549 7616 2613 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2549 7704 2613 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2549 7704 2613 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2549 7792 2613 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2549 7792 2613 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2549 7880 2613 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2549 7880 2613 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2549 7968 2613 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2549 7968 2613 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2622 10331 2686 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2622 10331 2686 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2622 10415 2686 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2622 10415 2686 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2622 10499 2686 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2622 10499 2686 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2623 9548 2687 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2623 9548 2687 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2623 11282 2687 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2623 11282 2687 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2630 7352 2694 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2630 7352 2694 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2630 7440 2694 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2630 7440 2694 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2630 7528 2694 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2630 7528 2694 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2630 7616 2694 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2630 7616 2694 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2630 7704 2694 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2630 7704 2694 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2630 7792 2694 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2630 7792 2694 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2630 7880 2694 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2630 7880 2694 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2630 7968 2694 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2630 7968 2694 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2703 10331 2767 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2703 10331 2767 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2703 10415 2767 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2703 10415 2767 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2703 10499 2767 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2703 10499 2767 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2704 9548 2768 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2704 9548 2768 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2704 11282 2768 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2704 11282 2768 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2711 7352 2775 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2711 7352 2775 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2711 7440 2775 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2711 7440 2775 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2711 7528 2775 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2711 7528 2775 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2711 7616 2775 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2711 7616 2775 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2711 7704 2775 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2711 7704 2775 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2711 7792 2775 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2711 7792 2775 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2711 7880 2775 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2711 7880 2775 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2711 7968 2775 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2711 7968 2775 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2784 10331 2848 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2784 10331 2848 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2784 10415 2848 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2784 10415 2848 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2784 10499 2848 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2784 10499 2848 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2785 9548 2849 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2785 9548 2849 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2785 11282 2849 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2785 11282 2849 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2792 7352 2856 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2792 7352 2856 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2792 7440 2856 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2792 7440 2856 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2792 7528 2856 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2792 7528 2856 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2792 7616 2856 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2792 7616 2856 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2792 7704 2856 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2792 7704 2856 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2792 7792 2856 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2792 7792 2856 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2792 7880 2856 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2792 7880 2856 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2792 7968 2856 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2792 7968 2856 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2865 10331 2929 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2865 10331 2929 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2865 10415 2929 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2865 10415 2929 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2865 10499 2929 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2865 10499 2929 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2866 9548 2930 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2866 9548 2930 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2866 11282 2930 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2866 11282 2930 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2873 7352 2937 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2873 7352 2937 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2873 7440 2937 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2873 7440 2937 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2873 7528 2937 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2873 7528 2937 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2873 7616 2937 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2873 7616 2937 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2873 7704 2937 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2873 7704 2937 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2873 7792 2937 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2873 7792 2937 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2873 7880 2937 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2873 7880 2937 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2873 7968 2937 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2873 7968 2937 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2946 10331 3010 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2946 10331 3010 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2946 10415 3010 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2946 10415 3010 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2946 10499 3010 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2946 10499 3010 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2947 9548 3011 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2947 9548 3011 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2947 11282 3011 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2947 11282 3011 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2954 7352 3018 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2954 7352 3018 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2954 7440 3018 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2954 7440 3018 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2954 7528 3018 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2954 7528 3018 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2954 7616 3018 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2954 7616 3018 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2954 7704 3018 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2954 7704 3018 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2954 7792 3018 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2954 7792 3018 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2954 7880 3018 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2954 7880 3018 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 2954 7968 3018 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 2954 7968 3018 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3027 10331 3091 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3027 10331 3091 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3027 10415 3091 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3027 10415 3091 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3027 10499 3091 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3027 10499 3091 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3028 9548 3092 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3028 9548 3092 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3028 11282 3092 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3028 11282 3092 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3035 7352 3099 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3035 7352 3099 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3035 7440 3099 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3035 7440 3099 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3035 7528 3099 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3035 7528 3099 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3035 7616 3099 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3035 7616 3099 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3035 7704 3099 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3035 7704 3099 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3035 7792 3099 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3035 7792 3099 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3035 7880 3099 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3035 7880 3099 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3035 7968 3099 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3035 7968 3099 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3108 10331 3172 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3108 10331 3172 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3108 10415 3172 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3108 10415 3172 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3108 10499 3172 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3108 10499 3172 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3109 9548 3173 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3109 9548 3173 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3109 11282 3173 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3109 11282 3173 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3116 7352 3180 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3116 7352 3180 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3116 7440 3180 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3116 7440 3180 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3116 7528 3180 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3116 7528 3180 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3116 7616 3180 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3116 7616 3180 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3116 7704 3180 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3116 7704 3180 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3116 7792 3180 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3116 7792 3180 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3116 7880 3180 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3116 7880 3180 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3116 7968 3180 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3116 7968 3180 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3189 10331 3253 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3189 10331 3253 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3189 10415 3253 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3189 10415 3253 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3189 10499 3253 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3189 10499 3253 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3190 9548 3254 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3190 9548 3254 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3190 11282 3254 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3190 11282 3254 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3197 7352 3261 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3197 7352 3261 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3197 7440 3261 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3197 7440 3261 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3197 7528 3261 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3197 7528 3261 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3197 7616 3261 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3197 7616 3261 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3197 7704 3261 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3197 7704 3261 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3197 7792 3261 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3197 7792 3261 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3197 7880 3261 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3197 7880 3261 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3197 7968 3261 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3197 7968 3261 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3270 10331 3334 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3270 10331 3334 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3270 10415 3334 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3270 10415 3334 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3270 10499 3334 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3270 10499 3334 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3271 9548 3335 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3271 9548 3335 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3271 11282 3335 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3271 11282 3335 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3278 7352 3342 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3278 7352 3342 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3278 7440 3342 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3278 7440 3342 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3278 7528 3342 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3278 7528 3342 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3278 7616 3342 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3278 7616 3342 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3278 7704 3342 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3278 7704 3342 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3278 7792 3342 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3278 7792 3342 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3278 7880 3342 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3278 7880 3342 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3278 7968 3342 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3278 7968 3342 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3351 10331 3415 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3351 10331 3415 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3351 10415 3415 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3351 10415 3415 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3351 10499 3415 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3351 10499 3415 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3352 9548 3416 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3352 9548 3416 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3352 11282 3416 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3352 11282 3416 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3359 7352 3423 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3359 7352 3423 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3359 7440 3423 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3359 7440 3423 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3359 7528 3423 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3359 7528 3423 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3359 7616 3423 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3359 7616 3423 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3359 7704 3423 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3359 7704 3423 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3359 7792 3423 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3359 7792 3423 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3359 7880 3423 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3359 7880 3423 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3359 7968 3423 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3359 7968 3423 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3432 10331 3496 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3432 10331 3496 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3432 10415 3496 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3432 10415 3496 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3432 10499 3496 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3432 10499 3496 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3433 9548 3497 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3433 9548 3497 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3433 11282 3497 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3433 11282 3497 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3440 7352 3504 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3440 7352 3504 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3440 7440 3504 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3440 7440 3504 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3440 7528 3504 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3440 7528 3504 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3440 7616 3504 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3440 7616 3504 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3440 7704 3504 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3440 7704 3504 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3440 7792 3504 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3440 7792 3504 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3440 7880 3504 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3440 7880 3504 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3440 7968 3504 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3440 7968 3504 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3513 10331 3577 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3513 10331 3577 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3513 10415 3577 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3513 10415 3577 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3513 10499 3577 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3513 10499 3577 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3514 9548 3578 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3514 9548 3578 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3514 11282 3578 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3514 11282 3578 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3521 7352 3585 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3521 7352 3585 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3521 7440 3585 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3521 7440 3585 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3521 7528 3585 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3521 7528 3585 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3521 7616 3585 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3521 7616 3585 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3521 7704 3585 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3521 7704 3585 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3521 7792 3585 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3521 7792 3585 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3521 7880 3585 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3521 7880 3585 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3521 7968 3585 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3521 7968 3585 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3594 10331 3658 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3594 10331 3658 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3594 10415 3658 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3594 10415 3658 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3594 10499 3658 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3594 10499 3658 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3595 9548 3659 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3595 9548 3659 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3595 11282 3659 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3595 11282 3659 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3602 7352 3666 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3602 7352 3666 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3602 7440 3666 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3602 7440 3666 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3602 7528 3666 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3602 7528 3666 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3602 7616 3666 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3602 7616 3666 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3602 7704 3666 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3602 7704 3666 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3602 7792 3666 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3602 7792 3666 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3602 7880 3666 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3602 7880 3666 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3602 7968 3666 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3602 7968 3666 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3675 10331 3739 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3675 10331 3739 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3675 10415 3739 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3675 10415 3739 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3675 10499 3739 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3675 10499 3739 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3676 9548 3740 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3676 9548 3740 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3676 11282 3740 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3676 11282 3740 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3683 7352 3747 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3683 7352 3747 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3683 7440 3747 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3683 7440 3747 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3683 7528 3747 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3683 7528 3747 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3683 7616 3747 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3683 7616 3747 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3683 7704 3747 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3683 7704 3747 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3683 7792 3747 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3683 7792 3747 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3683 7880 3747 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3683 7880 3747 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3683 7968 3747 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3683 7968 3747 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3756 10331 3820 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3756 10331 3820 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3756 10415 3820 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3756 10415 3820 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3756 10499 3820 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3756 10499 3820 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3757 9548 3821 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3757 9548 3821 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3757 11282 3821 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3757 11282 3821 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3764 7352 3828 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3764 7352 3828 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3764 7440 3828 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3764 7440 3828 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3764 7528 3828 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3764 7528 3828 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3764 7616 3828 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3764 7616 3828 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3764 7704 3828 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3764 7704 3828 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3764 7792 3828 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3764 7792 3828 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3764 7880 3828 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3764 7880 3828 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3764 7968 3828 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3764 7968 3828 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3837 10331 3901 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3837 10331 3901 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3837 10415 3901 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3837 10415 3901 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3837 10499 3901 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3837 10499 3901 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3838 9548 3902 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3838 9548 3902 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3838 11282 3902 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3838 11282 3902 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3845 7352 3909 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3845 7352 3909 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3845 7440 3909 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3845 7440 3909 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3845 7528 3909 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3845 7528 3909 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3845 7616 3909 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3845 7616 3909 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3845 7704 3909 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3845 7704 3909 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3845 7792 3909 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3845 7792 3909 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3845 7880 3909 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3845 7880 3909 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3845 7968 3909 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3845 7968 3909 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3918 10331 3982 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3918 10331 3982 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3918 10415 3982 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3918 10415 3982 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3918 10499 3982 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3918 10499 3982 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3919 9548 3983 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3919 9548 3983 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3919 11282 3983 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3919 11282 3983 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3926 7352 3990 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3926 7352 3990 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3926 7440 3990 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3926 7440 3990 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3926 7528 3990 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3926 7528 3990 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3926 7616 3990 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3926 7616 3990 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3926 7704 3990 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3926 7704 3990 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3926 7792 3990 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3926 7792 3990 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3926 7880 3990 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3926 7880 3990 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3926 7968 3990 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3926 7968 3990 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3999 10331 4063 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3999 10331 4063 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3999 10415 4063 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3999 10415 4063 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 3999 10499 4063 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 3999 10499 4063 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 433 10331 497 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 433 10331 497 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 433 10415 497 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 433 10415 497 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 433 10499 497 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 433 10499 497 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 436 9548 500 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 436 9548 500 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 436 11282 500 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 436 11282 500 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 443 7352 507 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 443 7352 507 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 443 7440 507 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 443 7440 507 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 443 7528 507 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 443 7528 507 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 443 7616 507 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 443 7616 507 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 443 7704 507 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 443 7704 507 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 443 7792 507 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 443 7792 507 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 443 7880 507 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 443 7880 507 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 443 7968 507 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 443 7968 507 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 515 10331 579 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 515 10331 579 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 515 10415 579 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 515 10415 579 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 515 10499 579 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 515 10499 579 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 517 9548 581 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 517 9548 581 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 517 11282 581 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 517 11282 581 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 524 7352 588 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 524 7352 588 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 524 7440 588 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 524 7440 588 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 524 7528 588 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 524 7528 588 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 524 7616 588 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 524 7616 588 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 524 7704 588 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 524 7704 588 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 524 7792 588 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 524 7792 588 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 524 7880 588 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 524 7880 588 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 524 7968 588 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 524 7968 588 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 597 10331 661 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 597 10331 661 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 597 10415 661 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 597 10415 661 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 597 10499 661 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 597 10499 661 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 598 9548 662 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 598 9548 662 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 598 11282 662 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 598 11282 662 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4000 9548 4064 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4000 9548 4064 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4000 11282 4064 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4000 11282 4064 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4007 7352 4071 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4007 7352 4071 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4007 7440 4071 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4007 7440 4071 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4007 7528 4071 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4007 7528 4071 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4007 7616 4071 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4007 7616 4071 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4007 7704 4071 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4007 7704 4071 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4007 7792 4071 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4007 7792 4071 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4007 7880 4071 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4007 7880 4071 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4007 7968 4071 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4007 7968 4071 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4080 10331 4144 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4080 10331 4144 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4080 10415 4144 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4080 10415 4144 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4080 10499 4144 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4080 10499 4144 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4081 9548 4145 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4081 9548 4145 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4081 11282 4145 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4081 11282 4145 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4088 7352 4152 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4088 7352 4152 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4088 7440 4152 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4088 7440 4152 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4088 7528 4152 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4088 7528 4152 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4088 7616 4152 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4088 7616 4152 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4088 7704 4152 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4088 7704 4152 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4088 7792 4152 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4088 7792 4152 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4088 7880 4152 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4088 7880 4152 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4088 7968 4152 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4088 7968 4152 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4161 10331 4225 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4161 10331 4225 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4161 10415 4225 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4161 10415 4225 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4161 10499 4225 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4161 10499 4225 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4162 9548 4226 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4162 9548 4226 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4162 11282 4226 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4162 11282 4226 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4169 7352 4233 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4169 7352 4233 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4169 7440 4233 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4169 7440 4233 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4169 7528 4233 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4169 7528 4233 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4169 7616 4233 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4169 7616 4233 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4169 7704 4233 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4169 7704 4233 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4169 7792 4233 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4169 7792 4233 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4169 7880 4233 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4169 7880 4233 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4169 7968 4233 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4169 7968 4233 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4242 10331 4306 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4242 10331 4306 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4242 10415 4306 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4242 10415 4306 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4242 10499 4306 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4242 10499 4306 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4243 9548 4307 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4243 9548 4307 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4243 11282 4307 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4243 11282 4307 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4249 7352 4313 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4249 7352 4313 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4249 7440 4313 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4249 7440 4313 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4249 7528 4313 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4249 7528 4313 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4249 7616 4313 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4249 7616 4313 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4249 7704 4313 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4249 7704 4313 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4249 7792 4313 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4249 7792 4313 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4249 7880 4313 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4249 7880 4313 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4249 7968 4313 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4249 7968 4313 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4323 10331 4387 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4323 10331 4387 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4323 10415 4387 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4323 10415 4387 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4323 10499 4387 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4323 10499 4387 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4324 9548 4388 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4324 9548 4388 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4324 11282 4388 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4324 11282 4388 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4329 7352 4393 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4329 7352 4393 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4329 7440 4393 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4329 7440 4393 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4329 7528 4393 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4329 7528 4393 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4329 7616 4393 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4329 7616 4393 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4329 7704 4393 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4329 7704 4393 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4329 7792 4393 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4329 7792 4393 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4329 7880 4393 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4329 7880 4393 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4329 7968 4393 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4329 7968 4393 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4404 10331 4468 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4404 10331 4468 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4404 10415 4468 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4404 10415 4468 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4404 10499 4468 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4404 10499 4468 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4405 9548 4469 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4405 9548 4469 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4405 11282 4469 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4405 11282 4469 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4409 7352 4473 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4409 7352 4473 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4409 7440 4473 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4409 7440 4473 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4409 7528 4473 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4409 7528 4473 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4409 7616 4473 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4409 7616 4473 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4409 7704 4473 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4409 7704 4473 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4409 7792 4473 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4409 7792 4473 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4409 7880 4473 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4409 7880 4473 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4409 7968 4473 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4409 7968 4473 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4485 10331 4549 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4485 10331 4549 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4485 10415 4549 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4485 10415 4549 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4485 10499 4549 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4485 10499 4549 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4486 9548 4550 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4486 9548 4550 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4486 11282 4550 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4486 11282 4550 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4489 7352 4553 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4489 7352 4553 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4489 7440 4553 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4489 7440 4553 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4489 7528 4553 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4489 7528 4553 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4489 7616 4553 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4489 7616 4553 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4489 7704 4553 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4489 7704 4553 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4489 7792 4553 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4489 7792 4553 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4489 7880 4553 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4489 7880 4553 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4489 7968 4553 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4489 7968 4553 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4566 10331 4630 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4566 10331 4630 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4566 10415 4630 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4566 10415 4630 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4566 10499 4630 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4566 10499 4630 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4567 9548 4631 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4567 9548 4631 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4567 11282 4631 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4567 11282 4631 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4569 7352 4633 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4569 7352 4633 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4569 7440 4633 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4569 7440 4633 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4569 7528 4633 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4569 7528 4633 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4569 7616 4633 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4569 7616 4633 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4569 7704 4633 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4569 7704 4633 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4569 7792 4633 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4569 7792 4633 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4569 7880 4633 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4569 7880 4633 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4569 7968 4633 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4569 7968 4633 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4647 10331 4711 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4647 10331 4711 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4647 10415 4711 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4647 10415 4711 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4647 10499 4711 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4647 10499 4711 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4648 9548 4712 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4648 9548 4712 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4648 11282 4712 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4648 11282 4712 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4649 7352 4713 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4649 7352 4713 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4649 7440 4713 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4649 7440 4713 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4649 7528 4713 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4649 7528 4713 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4649 7616 4713 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4649 7616 4713 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4649 7704 4713 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4649 7704 4713 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4649 7792 4713 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4649 7792 4713 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4649 7880 4713 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4649 7880 4713 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4649 7968 4713 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4649 7968 4713 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4728 10331 4792 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4728 10331 4792 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4728 10415 4792 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4728 10415 4792 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4728 10499 4792 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4728 10499 4792 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4729 7352 4793 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4729 7352 4793 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4729 7440 4793 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4729 7440 4793 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4729 7528 4793 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4729 7528 4793 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4729 7616 4793 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4729 7616 4793 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4729 7704 4793 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4729 7704 4793 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4729 7792 4793 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4729 7792 4793 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4729 7880 4793 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4729 7880 4793 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4729 7968 4793 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4729 7968 4793 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4729 9548 4793 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4729 9548 4793 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4729 11282 4793 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4729 11282 4793 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4809 7352 4873 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4809 7352 4873 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4809 7440 4873 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4809 7440 4873 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4809 7528 4873 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4809 7528 4873 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4809 7616 4873 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4809 7616 4873 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4809 7704 4873 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4809 7704 4873 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4809 7792 4873 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4809 7792 4873 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4809 7880 4873 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4809 7880 4873 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4809 7968 4873 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4809 7968 4873 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4809 9548 4873 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4809 9548 4873 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4809 10331 4873 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4809 10331 4873 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4809 10415 4873 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4809 10415 4873 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4809 10499 4873 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4809 10499 4873 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 4809 11282 4873 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 4809 11282 4873 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 605 7352 669 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 605 7352 669 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 605 7440 669 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 605 7440 669 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 605 7528 669 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 605 7528 669 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 605 7616 669 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 605 7616 669 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 605 7704 669 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 605 7704 669 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 605 7792 669 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 605 7792 669 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 605 7880 669 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 605 7880 669 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 605 7968 669 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 605 7968 669 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 678 10331 742 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 678 10331 742 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 678 10415 742 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 678 10415 742 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 678 10499 742 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 678 10499 742 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 679 9548 743 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 679 9548 743 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 679 11282 743 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 679 11282 743 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 686 7352 750 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 686 7352 750 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 686 7440 750 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 686 7440 750 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 686 7528 750 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 686 7528 750 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 686 7616 750 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 686 7616 750 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 686 7704 750 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 686 7704 750 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 686 7792 750 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 686 7792 750 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 686 7880 750 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 686 7880 750 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 686 7968 750 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 686 7968 750 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 759 10331 823 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 759 10331 823 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 759 10415 823 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 759 10415 823 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 759 10499 823 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 759 10499 823 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 760 9548 824 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 760 9548 824 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 760 11282 824 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 760 11282 824 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 767 7352 831 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 767 7352 831 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 767 7440 831 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 767 7440 831 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 767 7528 831 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 767 7528 831 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 767 7616 831 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 767 7616 831 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 767 7704 831 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 767 7704 831 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 767 7792 831 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 767 7792 831 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 767 7880 831 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 767 7880 831 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 767 7968 831 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 767 7968 831 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 840 10331 904 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 840 10331 904 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 840 10415 904 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 840 10415 904 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 840 10499 904 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 840 10499 904 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 841 9548 905 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 841 9548 905 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 841 11282 905 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 841 11282 905 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 848 7352 912 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 848 7352 912 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 848 7440 912 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 848 7440 912 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 848 7528 912 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 848 7528 912 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 848 7616 912 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 848 7616 912 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 848 7704 912 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 848 7704 912 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 848 7792 912 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 848 7792 912 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 848 7880 912 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 848 7880 912 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 848 7968 912 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 848 7968 912 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 921 10331 985 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 921 10331 985 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 921 10415 985 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 921 10415 985 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 921 10499 985 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 921 10499 985 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 922 9548 986 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 922 9548 986 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 922 11282 986 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 922 11282 986 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 929 7352 993 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 929 7352 993 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 929 7440 993 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 929 7440 993 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 929 7528 993 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 929 7528 993 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 929 7616 993 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 929 7616 993 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 929 7704 993 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 929 7704 993 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 929 7792 993 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 929 7792 993 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 929 7880 993 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 929 7880 993 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 929 7968 993 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 929 7968 993 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1002 10331 1066 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1002 10331 1066 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1002 10415 1066 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1002 10415 1066 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1002 10499 1066 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1002 10499 1066 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1003 9548 1067 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1003 9548 1067 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1003 11282 1067 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1003 11282 1067 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1010 7352 1074 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1010 7352 1074 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1010 7440 1074 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1010 7440 1074 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1010 7528 1074 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1010 7528 1074 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1010 7616 1074 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1010 7616 1074 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1010 7704 1074 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1010 7704 1074 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1010 7792 1074 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1010 7792 1074 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1010 7880 1074 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1010 7880 1074 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1010 7968 1074 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1010 7968 1074 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1083 10331 1147 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1083 10331 1147 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1083 10415 1147 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1083 10415 1147 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1083 10499 1147 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1083 10499 1147 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1084 9548 1148 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1084 9548 1148 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1084 11282 1148 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1084 11282 1148 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1091 7352 1155 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1091 7352 1155 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1091 7440 1155 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1091 7440 1155 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1091 7528 1155 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1091 7528 1155 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1091 7616 1155 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1091 7616 1155 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1091 7704 1155 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1091 7704 1155 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1091 7792 1155 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1091 7792 1155 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1091 7880 1155 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1091 7880 1155 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1091 7968 1155 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1091 7968 1155 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1164 10331 1228 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1164 10331 1228 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1164 10415 1228 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1164 10415 1228 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1164 10499 1228 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1164 10499 1228 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1165 9548 1229 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1165 9548 1229 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1165 11282 1229 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1165 11282 1229 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1172 7352 1236 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1172 7352 1236 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1172 7440 1236 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1172 7440 1236 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1172 7528 1236 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1172 7528 1236 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1172 7616 1236 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1172 7616 1236 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1172 7704 1236 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1172 7704 1236 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1172 7792 1236 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1172 7792 1236 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1172 7880 1236 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1172 7880 1236 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1172 7968 1236 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1172 7968 1236 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10084 7352 10148 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10084 7352 10148 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10084 7440 10148 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10084 7440 10148 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10084 7528 10148 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10084 7528 10148 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10084 7616 10148 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10084 7616 10148 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10084 7704 10148 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10084 7704 10148 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10084 7792 10148 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10084 7792 10148 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10084 7880 10148 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10084 7880 10148 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10084 7968 10148 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10084 7968 10148 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10084 9548 10148 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10084 9548 10148 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10084 10331 10148 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10084 10331 10148 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10084 10415 10148 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10084 10415 10148 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10084 10499 10148 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10084 10499 10148 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10084 11282 10148 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10084 11282 10148 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10165 9548 10229 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10165 9548 10229 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10165 11282 10229 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10165 11282 10229 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10166 7352 10230 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10166 7352 10230 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10166 7440 10230 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10166 7440 10230 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10166 7528 10230 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10166 7528 10230 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10166 7616 10230 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10166 7616 10230 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10166 7704 10230 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10166 7704 10230 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10166 7792 10230 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10166 7792 10230 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10166 7880 10230 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10166 7880 10230 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10166 7968 10230 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10166 7968 10230 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10166 10331 10230 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10166 10331 10230 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10166 10415 10230 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10166 10415 10230 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10166 10499 10230 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10166 10499 10230 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10246 9548 10310 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10246 9548 10310 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10246 11282 10310 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10246 11282 10310 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10248 7352 10312 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10248 7352 10312 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10248 7440 10312 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10248 7440 10312 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10248 7528 10312 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10248 7528 10312 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10248 7616 10312 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10248 7616 10312 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10248 7704 10312 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10248 7704 10312 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10248 7792 10312 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10248 7792 10312 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10248 7880 10312 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10248 7880 10312 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10248 7968 10312 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10248 7968 10312 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10248 10331 10312 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10248 10331 10312 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10248 10415 10312 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10248 10415 10312 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10248 10499 10312 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10248 10499 10312 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10327 9548 10391 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10327 9548 10391 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10327 11282 10391 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10327 11282 10391 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10330 7352 10394 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10330 7352 10394 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10330 7440 10394 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10330 7440 10394 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10330 7528 10394 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10330 7528 10394 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10330 7616 10394 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10330 7616 10394 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10330 7704 10394 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10330 7704 10394 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10330 7792 10394 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10330 7792 10394 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10330 7880 10394 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10330 7880 10394 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10330 7968 10394 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10330 7968 10394 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10330 10331 10394 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10330 10331 10394 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10330 10415 10394 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10330 10415 10394 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10330 10499 10394 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10330 10499 10394 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10408 9548 10472 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10408 9548 10472 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10408 11282 10472 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10408 11282 10472 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10412 7352 10476 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10412 7352 10476 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10412 7440 10476 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10412 7440 10476 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10412 7528 10476 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10412 7528 10476 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10412 7616 10476 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10412 7616 10476 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10412 7704 10476 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10412 7704 10476 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10412 7792 10476 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10412 7792 10476 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10412 7880 10476 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10412 7880 10476 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10412 7968 10476 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10412 7968 10476 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10412 10331 10476 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10412 10331 10476 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10412 10415 10476 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10412 10415 10476 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10412 10499 10476 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10412 10499 10476 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10489 9548 10553 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10489 9548 10553 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10489 11282 10553 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10489 11282 10553 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10494 7352 10558 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10494 7352 10558 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10494 7440 10558 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10494 7440 10558 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10494 7528 10558 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10494 7528 10558 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10494 7616 10558 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10494 7616 10558 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10494 7704 10558 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10494 7704 10558 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10494 7792 10558 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10494 7792 10558 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10494 7880 10558 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10494 7880 10558 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10494 7968 10558 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10494 7968 10558 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10494 10331 10558 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10494 10331 10558 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10494 10415 10558 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10494 10415 10558 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10494 10499 10558 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10494 10499 10558 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10570 9548 10634 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10570 9548 10634 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10570 11282 10634 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10570 11282 10634 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10576 7352 10640 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10576 7352 10640 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10576 7440 10640 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10576 7440 10640 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10576 7528 10640 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10576 7528 10640 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10576 7616 10640 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10576 7616 10640 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10576 7704 10640 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10576 7704 10640 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10576 7792 10640 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10576 7792 10640 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10576 7880 10640 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10576 7880 10640 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10576 7968 10640 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10576 7968 10640 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10576 10331 10640 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10576 10331 10640 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10576 10415 10640 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10576 10415 10640 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10576 10499 10640 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10576 10499 10640 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10651 9548 10715 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10651 9548 10715 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10651 11282 10715 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10651 11282 10715 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10657 7352 10721 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10657 7352 10721 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10657 7440 10721 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10657 7440 10721 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10657 7528 10721 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10657 7528 10721 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10657 7616 10721 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10657 7616 10721 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10657 7704 10721 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10657 7704 10721 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10657 7792 10721 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10657 7792 10721 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10657 7880 10721 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10657 7880 10721 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10657 7968 10721 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10657 7968 10721 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10657 10331 10721 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10657 10331 10721 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10657 10415 10721 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10657 10415 10721 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10657 10499 10721 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10657 10499 10721 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10732 9548 10796 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10732 9548 10796 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10732 11282 10796 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10732 11282 10796 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10738 7352 10802 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10738 7352 10802 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10738 7440 10802 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10738 7440 10802 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10738 7528 10802 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10738 7528 10802 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10738 7616 10802 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10738 7616 10802 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10738 7704 10802 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10738 7704 10802 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10738 7792 10802 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10738 7792 10802 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10738 7880 10802 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10738 7880 10802 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10738 7968 10802 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10738 7968 10802 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10738 10331 10802 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10738 10331 10802 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10738 10415 10802 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10738 10415 10802 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10738 10499 10802 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10738 10499 10802 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10813 9548 10877 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10813 9548 10877 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10813 11282 10877 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10813 11282 10877 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10819 7352 10883 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10819 7352 10883 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10819 7440 10883 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10819 7440 10883 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10819 7528 10883 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10819 7528 10883 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10819 7616 10883 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10819 7616 10883 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10819 7704 10883 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10819 7704 10883 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10819 7792 10883 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10819 7792 10883 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10819 7880 10883 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10819 7880 10883 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10819 7968 10883 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10819 7968 10883 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10819 10331 10883 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10819 10331 10883 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10819 10415 10883 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10819 10415 10883 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10819 10499 10883 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10819 10499 10883 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10894 9548 10958 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10894 9548 10958 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10894 11282 10958 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10894 11282 10958 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10900 7352 10964 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10900 7352 10964 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10900 7440 10964 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10900 7440 10964 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10900 7528 10964 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10900 7528 10964 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10900 7616 10964 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10900 7616 10964 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10900 7704 10964 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10900 7704 10964 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10900 7792 10964 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10900 7792 10964 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10900 7880 10964 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10900 7880 10964 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10900 7968 10964 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10900 7968 10964 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10900 10331 10964 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10900 10331 10964 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10900 10415 10964 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10900 10415 10964 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10900 10499 10964 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10900 10499 10964 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10975 9548 11039 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10975 9548 11039 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10975 11282 11039 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10975 11282 11039 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10981 7352 11045 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10981 7352 11045 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10981 7440 11045 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10981 7440 11045 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10981 7528 11045 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10981 7528 11045 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10981 7616 11045 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10981 7616 11045 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10981 7704 11045 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10981 7704 11045 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10981 7792 11045 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10981 7792 11045 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10981 7880 11045 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10981 7880 11045 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10981 7968 11045 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10981 7968 11045 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10981 10331 11045 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10981 10331 11045 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10981 10415 11045 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10981 10415 11045 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 10981 10499 11045 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 10981 10499 11045 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11056 9548 11120 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11056 9548 11120 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11056 11282 11120 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11056 11282 11120 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11062 7352 11126 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11062 7352 11126 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11062 7440 11126 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11062 7440 11126 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11062 7528 11126 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11062 7528 11126 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11062 7616 11126 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11062 7616 11126 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11062 7704 11126 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11062 7704 11126 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11062 7792 11126 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11062 7792 11126 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11062 7880 11126 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11062 7880 11126 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11062 7968 11126 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11062 7968 11126 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11062 10331 11126 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11062 10331 11126 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11062 10415 11126 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11062 10415 11126 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11062 10499 11126 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11062 10499 11126 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11137 9548 11201 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11137 9548 11201 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11137 11282 11201 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11137 11282 11201 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11143 7352 11207 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11143 7352 11207 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11143 7440 11207 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11143 7440 11207 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11143 7528 11207 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11143 7528 11207 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11143 7616 11207 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11143 7616 11207 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11143 7704 11207 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11143 7704 11207 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11143 7792 11207 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11143 7792 11207 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11143 7880 11207 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11143 7880 11207 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11143 7968 11207 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11143 7968 11207 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11143 10331 11207 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11143 10331 11207 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11143 10415 11207 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11143 10415 11207 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11143 10499 11207 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11143 10499 11207 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11218 9548 11282 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11218 9548 11282 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11218 11282 11282 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11218 11282 11282 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11224 7352 11288 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11224 7352 11288 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11224 7440 11288 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11224 7440 11288 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11224 7528 11288 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11224 7528 11288 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11224 7616 11288 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11224 7616 11288 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11224 7704 11288 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11224 7704 11288 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11224 7792 11288 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11224 7792 11288 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11224 7880 11288 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11224 7880 11288 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11224 7968 11288 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11224 7968 11288 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11224 10331 11288 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11224 10331 11288 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11224 10415 11288 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11224 10415 11288 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11224 10499 11288 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11224 10499 11288 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11299 9548 11363 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11299 9548 11363 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11299 11282 11363 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11299 11282 11363 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11305 7352 11369 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11305 7352 11369 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11305 7440 11369 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11305 7440 11369 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11305 7528 11369 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11305 7528 11369 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11305 7616 11369 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11305 7616 11369 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11305 7704 11369 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11305 7704 11369 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11305 7792 11369 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11305 7792 11369 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11305 7880 11369 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11305 7880 11369 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11305 7968 11369 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11305 7968 11369 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11305 10331 11369 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11305 10331 11369 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11305 10415 11369 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11305 10415 11369 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11305 10499 11369 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11305 10499 11369 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11380 9548 11444 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11380 9548 11444 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11380 11282 11444 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11380 11282 11444 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11386 7352 11450 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11386 7352 11450 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11386 7440 11450 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11386 7440 11450 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11386 7528 11450 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11386 7528 11450 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11386 7616 11450 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11386 7616 11450 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11386 7704 11450 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11386 7704 11450 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11386 7792 11450 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11386 7792 11450 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11386 7880 11450 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11386 7880 11450 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11386 7968 11450 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11386 7968 11450 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11386 10331 11450 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11386 10331 11450 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11386 10415 11450 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11386 10415 11450 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11386 10499 11450 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11386 10499 11450 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11461 9548 11525 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11461 9548 11525 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11461 11282 11525 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11461 11282 11525 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11467 7352 11531 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11467 7352 11531 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11467 7440 11531 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11467 7440 11531 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11467 7528 11531 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11467 7528 11531 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11467 7616 11531 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11467 7616 11531 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11467 7704 11531 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11467 7704 11531 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11467 7792 11531 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11467 7792 11531 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11467 7880 11531 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11467 7880 11531 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11467 7968 11531 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11467 7968 11531 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11467 10331 11531 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11467 10331 11531 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11467 10415 11531 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11467 10415 11531 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11467 10499 11531 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11467 10499 11531 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11542 9548 11606 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11542 9548 11606 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11542 11282 11606 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11542 11282 11606 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11548 7352 11612 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11548 7352 11612 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11548 7440 11612 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11548 7440 11612 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11548 7528 11612 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11548 7528 11612 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11548 7616 11612 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11548 7616 11612 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11548 7704 11612 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11548 7704 11612 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11548 7792 11612 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11548 7792 11612 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11548 7880 11612 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11548 7880 11612 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11548 7968 11612 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11548 7968 11612 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11548 10331 11612 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11548 10331 11612 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11548 10415 11612 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11548 10415 11612 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11548 10499 11612 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11548 10499 11612 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11623 9548 11687 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11623 9548 11687 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11623 11282 11687 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11623 11282 11687 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11629 7352 11693 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11629 7352 11693 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11629 7440 11693 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11629 7440 11693 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11629 7528 11693 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11629 7528 11693 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11629 7616 11693 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11629 7616 11693 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11629 7704 11693 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11629 7704 11693 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11629 7792 11693 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11629 7792 11693 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11629 7880 11693 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11629 7880 11693 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11629 7968 11693 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11629 7968 11693 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11629 10331 11693 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11629 10331 11693 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11629 10415 11693 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11629 10415 11693 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11629 10499 11693 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11629 10499 11693 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11704 9548 11768 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11704 9548 11768 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11704 11282 11768 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11704 11282 11768 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11710 7352 11774 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11710 7352 11774 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11710 7440 11774 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11710 7440 11774 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11710 7528 11774 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11710 7528 11774 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11710 7616 11774 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11710 7616 11774 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11710 7704 11774 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11710 7704 11774 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11710 7792 11774 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11710 7792 11774 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11710 7880 11774 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11710 7880 11774 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11710 7968 11774 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11710 7968 11774 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11710 10331 11774 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11710 10331 11774 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11710 10415 11774 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11710 10415 11774 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11710 10499 11774 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11710 10499 11774 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11785 9548 11849 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11785 9548 11849 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11785 11282 11849 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11785 11282 11849 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11791 7352 11855 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11791 7352 11855 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11791 7440 11855 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11791 7440 11855 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11791 7528 11855 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11791 7528 11855 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11791 7616 11855 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11791 7616 11855 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11791 7704 11855 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11791 7704 11855 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11791 7792 11855 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11791 7792 11855 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11791 7880 11855 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11791 7880 11855 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11791 7968 11855 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11791 7968 11855 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11791 10331 11855 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11791 10331 11855 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11791 10415 11855 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11791 10415 11855 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11791 10499 11855 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11791 10499 11855 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11866 9548 11930 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11866 9548 11930 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11866 11282 11930 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11866 11282 11930 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11872 7352 11936 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11872 7352 11936 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11872 7440 11936 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11872 7440 11936 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11872 7528 11936 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11872 7528 11936 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11872 7616 11936 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11872 7616 11936 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11872 7704 11936 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11872 7704 11936 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11872 7792 11936 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11872 7792 11936 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11872 7880 11936 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11872 7880 11936 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11872 7968 11936 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11872 7968 11936 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11872 10331 11936 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11872 10331 11936 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11872 10415 11936 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11872 10415 11936 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11872 10499 11936 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11872 10499 11936 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11947 9548 12011 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11947 9548 12011 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11947 11282 12011 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11947 11282 12011 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11953 7352 12017 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11953 7352 12017 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11953 7440 12017 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11953 7440 12017 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11953 7528 12017 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11953 7528 12017 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11953 7616 12017 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11953 7616 12017 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11953 7704 12017 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11953 7704 12017 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11953 7792 12017 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11953 7792 12017 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11953 7880 12017 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11953 7880 12017 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11953 7968 12017 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11953 7968 12017 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11953 10331 12017 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11953 10331 12017 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11953 10415 12017 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11953 10415 12017 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 11953 10499 12017 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 11953 10499 12017 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1245 10331 1309 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1245 10331 1309 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1245 10415 1309 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1245 10415 1309 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1245 10499 1309 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1245 10499 1309 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1246 9548 1310 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1246 9548 1310 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1246 11282 1310 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1246 11282 1310 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1253 7352 1317 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1253 7352 1317 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1253 7440 1317 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1253 7440 1317 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1253 7528 1317 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1253 7528 1317 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1253 7616 1317 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1253 7616 1317 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1253 7704 1317 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1253 7704 1317 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1253 7792 1317 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1253 7792 1317 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1253 7880 1317 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1253 7880 1317 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1253 7968 1317 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1253 7968 1317 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1326 10331 1390 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1326 10331 1390 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1326 10415 1390 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1326 10415 1390 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1326 10499 1390 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1326 10499 1390 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1327 9548 1391 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1327 9548 1391 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1327 11282 1391 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1327 11282 1391 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1334 7352 1398 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1334 7352 1398 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1334 7440 1398 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1334 7440 1398 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1334 7528 1398 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1334 7528 1398 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1334 7616 1398 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1334 7616 1398 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1334 7704 1398 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1334 7704 1398 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1334 7792 1398 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1334 7792 1398 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1334 7880 1398 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1334 7880 1398 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1334 7968 1398 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1334 7968 1398 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12028 9548 12092 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12028 9548 12092 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12028 11282 12092 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12028 11282 12092 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12034 7352 12098 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12034 7352 12098 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12034 7440 12098 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12034 7440 12098 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12034 7528 12098 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12034 7528 12098 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12034 7616 12098 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12034 7616 12098 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12034 7704 12098 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12034 7704 12098 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12034 7792 12098 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12034 7792 12098 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12034 7880 12098 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12034 7880 12098 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12034 7968 12098 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12034 7968 12098 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12034 10331 12098 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12034 10331 12098 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12034 10415 12098 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12034 10415 12098 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12034 10499 12098 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12034 10499 12098 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12109 9548 12173 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12109 9548 12173 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12109 11282 12173 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12109 11282 12173 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12115 7352 12179 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12115 7352 12179 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12115 7440 12179 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12115 7440 12179 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12115 7528 12179 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12115 7528 12179 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12115 7616 12179 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12115 7616 12179 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12115 7704 12179 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12115 7704 12179 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12115 7792 12179 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12115 7792 12179 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12115 7880 12179 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12115 7880 12179 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12115 7968 12179 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12115 7968 12179 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12115 10331 12179 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12115 10331 12179 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12115 10415 12179 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12115 10415 12179 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12115 10499 12179 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12115 10499 12179 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12190 9548 12254 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12190 9548 12254 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12190 11282 12254 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12190 11282 12254 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12196 7352 12260 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12196 7352 12260 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12196 7440 12260 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12196 7440 12260 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12196 7528 12260 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12196 7528 12260 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12196 7616 12260 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12196 7616 12260 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12196 7704 12260 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12196 7704 12260 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12196 7792 12260 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12196 7792 12260 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12196 7880 12260 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12196 7880 12260 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12196 7968 12260 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12196 7968 12260 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12196 10331 12260 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12196 10331 12260 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12196 10415 12260 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12196 10415 12260 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12196 10499 12260 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12196 10499 12260 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12271 9548 12335 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12271 9548 12335 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12271 11282 12335 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12271 11282 12335 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12277 7352 12341 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12277 7352 12341 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12277 7440 12341 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12277 7440 12341 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12277 7528 12341 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12277 7528 12341 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12277 7616 12341 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12277 7616 12341 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12277 7704 12341 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12277 7704 12341 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12277 7792 12341 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12277 7792 12341 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12277 7880 12341 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12277 7880 12341 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12277 7968 12341 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12277 7968 12341 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12277 10331 12341 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12277 10331 12341 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12277 10415 12341 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12277 10415 12341 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12277 10499 12341 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12277 10499 12341 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12352 9548 12416 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12352 9548 12416 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12352 11282 12416 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12352 11282 12416 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12358 7352 12422 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12358 7352 12422 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12358 7440 12422 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12358 7440 12422 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12358 7528 12422 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12358 7528 12422 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12358 7616 12422 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12358 7616 12422 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12358 7704 12422 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12358 7704 12422 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12358 7792 12422 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12358 7792 12422 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12358 7880 12422 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12358 7880 12422 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12358 7968 12422 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12358 7968 12422 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12358 10331 12422 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12358 10331 12422 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12358 10415 12422 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12358 10415 12422 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12358 10499 12422 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12358 10499 12422 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12433 9548 12497 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12433 9548 12497 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12433 11282 12497 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12433 11282 12497 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12439 7352 12503 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12439 7352 12503 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12439 7440 12503 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12439 7440 12503 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12439 7528 12503 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12439 7528 12503 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12439 7616 12503 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12439 7616 12503 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12439 7704 12503 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12439 7704 12503 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12439 7792 12503 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12439 7792 12503 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12439 7880 12503 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12439 7880 12503 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12439 7968 12503 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12439 7968 12503 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12439 10331 12503 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12439 10331 12503 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12439 10415 12503 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12439 10415 12503 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12439 10499 12503 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12439 10499 12503 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12514 9548 12578 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12514 9548 12578 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12514 11282 12578 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12514 11282 12578 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12520 7352 12584 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12520 7352 12584 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12520 7440 12584 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12520 7440 12584 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12520 7528 12584 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12520 7528 12584 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12520 7616 12584 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12520 7616 12584 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12520 7704 12584 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12520 7704 12584 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12520 7792 12584 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12520 7792 12584 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12520 7880 12584 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12520 7880 12584 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12520 7968 12584 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12520 7968 12584 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12520 10331 12584 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12520 10331 12584 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12520 10415 12584 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12520 10415 12584 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12520 10499 12584 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12520 10499 12584 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12595 9548 12659 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12595 9548 12659 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12595 11282 12659 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12595 11282 12659 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12601 7352 12665 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12601 7352 12665 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12601 7440 12665 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12601 7440 12665 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12601 7528 12665 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12601 7528 12665 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12601 7616 12665 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12601 7616 12665 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12601 7704 12665 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12601 7704 12665 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12601 7792 12665 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12601 7792 12665 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12601 7880 12665 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12601 7880 12665 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12601 7968 12665 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12601 7968 12665 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12601 10331 12665 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12601 10331 12665 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12601 10415 12665 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12601 10415 12665 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12601 10499 12665 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12601 10499 12665 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12676 9548 12740 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12676 9548 12740 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12676 11282 12740 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12676 11282 12740 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12682 7352 12746 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12682 7352 12746 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12682 7440 12746 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12682 7440 12746 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12682 7528 12746 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12682 7528 12746 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12682 7616 12746 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12682 7616 12746 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12682 7704 12746 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12682 7704 12746 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12682 7792 12746 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12682 7792 12746 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12682 7880 12746 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12682 7880 12746 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12682 7968 12746 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12682 7968 12746 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12682 10331 12746 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12682 10331 12746 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12682 10415 12746 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12682 10415 12746 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12682 10499 12746 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12682 10499 12746 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12757 9548 12821 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12757 9548 12821 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12757 11282 12821 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12757 11282 12821 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12763 7352 12827 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12763 7352 12827 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12763 7440 12827 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12763 7440 12827 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12763 7528 12827 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12763 7528 12827 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12763 7616 12827 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12763 7616 12827 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12763 7704 12827 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12763 7704 12827 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12763 7792 12827 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12763 7792 12827 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12763 7880 12827 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12763 7880 12827 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12763 7968 12827 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12763 7968 12827 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12763 10331 12827 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12763 10331 12827 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12763 10415 12827 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12763 10415 12827 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12763 10499 12827 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12763 10499 12827 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12838 9548 12902 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12838 9548 12902 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12838 11282 12902 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12838 11282 12902 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12844 7352 12908 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12844 7352 12908 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12844 7440 12908 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12844 7440 12908 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12844 7528 12908 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12844 7528 12908 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12844 7616 12908 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12844 7616 12908 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12844 7704 12908 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12844 7704 12908 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12844 7792 12908 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12844 7792 12908 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12844 7880 12908 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12844 7880 12908 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12844 7968 12908 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12844 7968 12908 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12844 10331 12908 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12844 10331 12908 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12844 10415 12908 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12844 10415 12908 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12844 10499 12908 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12844 10499 12908 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12919 9548 12983 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12919 9548 12983 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12919 11282 12983 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12919 11282 12983 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12925 7352 12989 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12925 7352 12989 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12925 7440 12989 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12925 7440 12989 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12925 7528 12989 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12925 7528 12989 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12925 7616 12989 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12925 7616 12989 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12925 7704 12989 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12925 7704 12989 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12925 7792 12989 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12925 7792 12989 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12925 7880 12989 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12925 7880 12989 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12925 7968 12989 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12925 7968 12989 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12925 10331 12989 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12925 10331 12989 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12925 10415 12989 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12925 10415 12989 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 12925 10499 12989 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 12925 10499 12989 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13000 9548 13064 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13000 9548 13064 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13000 11282 13064 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13000 11282 13064 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13006 7352 13070 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13006 7352 13070 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13006 7440 13070 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13006 7440 13070 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13006 7528 13070 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13006 7528 13070 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13006 7616 13070 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13006 7616 13070 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13006 7704 13070 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13006 7704 13070 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13006 7792 13070 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13006 7792 13070 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13006 7880 13070 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13006 7880 13070 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13006 7968 13070 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13006 7968 13070 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13006 10331 13070 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13006 10331 13070 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13006 10415 13070 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13006 10415 13070 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13006 10499 13070 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13006 10499 13070 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13081 9548 13145 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13081 9548 13145 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13081 11282 13145 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13081 11282 13145 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13087 7352 13151 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13087 7352 13151 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13087 7440 13151 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13087 7440 13151 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13087 7528 13151 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13087 7528 13151 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13087 7616 13151 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13087 7616 13151 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13087 7704 13151 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13087 7704 13151 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13087 7792 13151 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13087 7792 13151 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13087 7880 13151 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13087 7880 13151 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13087 7968 13151 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13087 7968 13151 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13087 10331 13151 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13087 10331 13151 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13087 10415 13151 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13087 10415 13151 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13087 10499 13151 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13087 10499 13151 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13162 9548 13226 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13162 9548 13226 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13162 11282 13226 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13162 11282 13226 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13168 7352 13232 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13168 7352 13232 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13168 7440 13232 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13168 7440 13232 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13168 7528 13232 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13168 7528 13232 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13168 7616 13232 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13168 7616 13232 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13168 7704 13232 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13168 7704 13232 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13168 7792 13232 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13168 7792 13232 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13168 7880 13232 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13168 7880 13232 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13168 7968 13232 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13168 7968 13232 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13168 10331 13232 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13168 10331 13232 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13168 10415 13232 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13168 10415 13232 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13168 10499 13232 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13168 10499 13232 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13243 9548 13307 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13243 9548 13307 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13243 11282 13307 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13243 11282 13307 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13249 7352 13313 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13249 7352 13313 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13249 7440 13313 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13249 7440 13313 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13249 7528 13313 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13249 7528 13313 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13249 7616 13313 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13249 7616 13313 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13249 7704 13313 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13249 7704 13313 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13249 7792 13313 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13249 7792 13313 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13249 7880 13313 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13249 7880 13313 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13249 7968 13313 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13249 7968 13313 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13249 10331 13313 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13249 10331 13313 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13249 10415 13313 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13249 10415 13313 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13249 10499 13313 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13249 10499 13313 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13324 9548 13388 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13324 9548 13388 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13324 11282 13388 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13324 11282 13388 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13330 7352 13394 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13330 7352 13394 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13330 7440 13394 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13330 7440 13394 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13330 7528 13394 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13330 7528 13394 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13330 7616 13394 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13330 7616 13394 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13330 7704 13394 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13330 7704 13394 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13330 7792 13394 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13330 7792 13394 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13330 7880 13394 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13330 7880 13394 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13330 7968 13394 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13330 7968 13394 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13330 10331 13394 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13330 10331 13394 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13330 10415 13394 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13330 10415 13394 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13330 10499 13394 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13330 10499 13394 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13405 9548 13469 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13405 9548 13469 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13405 11282 13469 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13405 11282 13469 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13411 7352 13475 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13411 7352 13475 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13411 7440 13475 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13411 7440 13475 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13411 7528 13475 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13411 7528 13475 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13411 7616 13475 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13411 7616 13475 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13411 7704 13475 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13411 7704 13475 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13411 7792 13475 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13411 7792 13475 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13411 7880 13475 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13411 7880 13475 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13411 7968 13475 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13411 7968 13475 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13411 10331 13475 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13411 10331 13475 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13411 10415 13475 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13411 10415 13475 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13411 10499 13475 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13411 10499 13475 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13486 9548 13550 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13486 9548 13550 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13486 11282 13550 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13486 11282 13550 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13492 7352 13556 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13492 7352 13556 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13492 7440 13556 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13492 7440 13556 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13492 7528 13556 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13492 7528 13556 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13492 7616 13556 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13492 7616 13556 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13492 7704 13556 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13492 7704 13556 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13492 7792 13556 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13492 7792 13556 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13492 7880 13556 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13492 7880 13556 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13492 7968 13556 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13492 7968 13556 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13492 10331 13556 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13492 10331 13556 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13492 10415 13556 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13492 10415 13556 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13492 10499 13556 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13492 10499 13556 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13567 9548 13631 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13567 9548 13631 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13567 11282 13631 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13567 11282 13631 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13573 7352 13637 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13573 7352 13637 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13573 7440 13637 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13573 7440 13637 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13573 7528 13637 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13573 7528 13637 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13573 7616 13637 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13573 7616 13637 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13573 7704 13637 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13573 7704 13637 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13573 7792 13637 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13573 7792 13637 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13573 7880 13637 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13573 7880 13637 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13573 7968 13637 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13573 7968 13637 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13573 10331 13637 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13573 10331 13637 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13573 10415 13637 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13573 10415 13637 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13573 10499 13637 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13573 10499 13637 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13648 9548 13712 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13648 9548 13712 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13648 11282 13712 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13648 11282 13712 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13654 7352 13718 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13654 7352 13718 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13654 7440 13718 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13654 7440 13718 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13654 7528 13718 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13654 7528 13718 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13654 7616 13718 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13654 7616 13718 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13654 7704 13718 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13654 7704 13718 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13654 7792 13718 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13654 7792 13718 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13654 7880 13718 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13654 7880 13718 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13654 7968 13718 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13654 7968 13718 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13654 10331 13718 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13654 10331 13718 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13654 10415 13718 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13654 10415 13718 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13654 10499 13718 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13654 10499 13718 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13729 9548 13793 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13729 9548 13793 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13729 11282 13793 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13729 11282 13793 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13735 7352 13799 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13735 7352 13799 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13735 7440 13799 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13735 7440 13799 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13735 7528 13799 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13735 7528 13799 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13735 7616 13799 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13735 7616 13799 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13735 7704 13799 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13735 7704 13799 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13735 7792 13799 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13735 7792 13799 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13735 7880 13799 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13735 7880 13799 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13735 7968 13799 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13735 7968 13799 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13735 10331 13799 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13735 10331 13799 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13735 10415 13799 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13735 10415 13799 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13735 10499 13799 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13735 10499 13799 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13810 9548 13874 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13810 9548 13874 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13810 11282 13874 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13810 11282 13874 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13816 7352 13880 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13816 7352 13880 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13816 7440 13880 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13816 7440 13880 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13816 7528 13880 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13816 7528 13880 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13816 7616 13880 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13816 7616 13880 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13816 7704 13880 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13816 7704 13880 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13816 7792 13880 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13816 7792 13880 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13816 7880 13880 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13816 7880 13880 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13816 7968 13880 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13816 7968 13880 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13816 10331 13880 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13816 10331 13880 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13816 10415 13880 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13816 10415 13880 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13816 10499 13880 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13816 10499 13880 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13891 9548 13955 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13891 9548 13955 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13891 11282 13955 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13891 11282 13955 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13897 7352 13961 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13897 7352 13961 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13897 7440 13961 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13897 7440 13961 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13897 7528 13961 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13897 7528 13961 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13897 7616 13961 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13897 7616 13961 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13897 7704 13961 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13897 7704 13961 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13897 7792 13961 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13897 7792 13961 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13897 7880 13961 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13897 7880 13961 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13897 7968 13961 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13897 7968 13961 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13897 10331 13961 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13897 10331 13961 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13897 10415 13961 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13897 10415 13961 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13897 10499 13961 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13897 10499 13961 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13972 9548 14036 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13972 9548 14036 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13972 11282 14036 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13972 11282 14036 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13978 7352 14042 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13978 7352 14042 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13978 7440 14042 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13978 7440 14042 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13978 7528 14042 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13978 7528 14042 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13978 7616 14042 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13978 7616 14042 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13978 7704 14042 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13978 7704 14042 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13978 7792 14042 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13978 7792 14042 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13978 7880 14042 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13978 7880 14042 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13978 7968 14042 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13978 7968 14042 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13978 10331 14042 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13978 10331 14042 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13978 10415 14042 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13978 10415 14042 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 13978 10499 14042 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 13978 10499 14042 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1407 10331 1471 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1407 10331 1471 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1407 10415 1471 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1407 10415 1471 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1407 10499 1471 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1407 10499 1471 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1408 9548 1472 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1408 9548 1472 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1408 11282 1472 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1408 11282 1472 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1415 7352 1479 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1415 7352 1479 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1415 7440 1479 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1415 7440 1479 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1415 7528 1479 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1415 7528 1479 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1415 7616 1479 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1415 7616 1479 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1415 7704 1479 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1415 7704 1479 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1415 7792 1479 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1415 7792 1479 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1415 7880 1479 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1415 7880 1479 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1415 7968 1479 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1415 7968 1479 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1488 10331 1552 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1488 10331 1552 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1488 10415 1552 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1488 10415 1552 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1488 10499 1552 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1488 10499 1552 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1489 9548 1553 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1489 9548 1553 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1489 11282 1553 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1489 11282 1553 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1496 7352 1560 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1496 7352 1560 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1496 7440 1560 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1496 7440 1560 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1496 7528 1560 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1496 7528 1560 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1496 7616 1560 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1496 7616 1560 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1496 7704 1560 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1496 7704 1560 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1496 7792 1560 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1496 7792 1560 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1496 7880 1560 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1496 7880 1560 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1496 7968 1560 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1496 7968 1560 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1569 10331 1633 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1569 10331 1633 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1569 10415 1633 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1569 10415 1633 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1569 10499 1633 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1569 10499 1633 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1570 9548 1634 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1570 9548 1634 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1570 11282 1634 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1570 11282 1634 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1577 7352 1641 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1577 7352 1641 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1577 7440 1641 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1577 7440 1641 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1577 7528 1641 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1577 7528 1641 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1577 7616 1641 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1577 7616 1641 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1577 7704 1641 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1577 7704 1641 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1577 7792 1641 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1577 7792 1641 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1577 7880 1641 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1577 7880 1641 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1577 7968 1641 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1577 7968 1641 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14053 9548 14117 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14053 9548 14117 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14053 11282 14117 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14053 11282 14117 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14059 7352 14123 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14059 7352 14123 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14059 7440 14123 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14059 7440 14123 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14059 7528 14123 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14059 7528 14123 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14059 7616 14123 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14059 7616 14123 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14059 7704 14123 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14059 7704 14123 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14059 7792 14123 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14059 7792 14123 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14059 7880 14123 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14059 7880 14123 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14059 7968 14123 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14059 7968 14123 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14059 10331 14123 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14059 10331 14123 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14059 10415 14123 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14059 10415 14123 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14059 10499 14123 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14059 10499 14123 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14134 9548 14198 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14134 9548 14198 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14134 11282 14198 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14134 11282 14198 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14140 7352 14204 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14140 7352 14204 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14140 7440 14204 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14140 7440 14204 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14140 7528 14204 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14140 7528 14204 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14140 7616 14204 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14140 7616 14204 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14140 7704 14204 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14140 7704 14204 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14140 7792 14204 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14140 7792 14204 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14140 7880 14204 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14140 7880 14204 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14140 7968 14204 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14140 7968 14204 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14140 10331 14204 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14140 10331 14204 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14140 10415 14204 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14140 10415 14204 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14140 10499 14204 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14140 10499 14204 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14215 9548 14279 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14215 9548 14279 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14215 11282 14279 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14215 11282 14279 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14221 7352 14285 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14221 7352 14285 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14221 7440 14285 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14221 7440 14285 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14221 7528 14285 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14221 7528 14285 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14221 7616 14285 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14221 7616 14285 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14221 7704 14285 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14221 7704 14285 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14221 7792 14285 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14221 7792 14285 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14221 7880 14285 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14221 7880 14285 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14221 7968 14285 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14221 7968 14285 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14221 10331 14285 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14221 10331 14285 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14221 10415 14285 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14221 10415 14285 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14221 10499 14285 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14221 10499 14285 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14296 9548 14360 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14296 9548 14360 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14296 11282 14360 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14296 11282 14360 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14302 7352 14366 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14302 7352 14366 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14302 7440 14366 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14302 7440 14366 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14302 7528 14366 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14302 7528 14366 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14302 7616 14366 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14302 7616 14366 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14302 7704 14366 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14302 7704 14366 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14302 7792 14366 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14302 7792 14366 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14302 7880 14366 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14302 7880 14366 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14302 7968 14366 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14302 7968 14366 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14302 10331 14366 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14302 10331 14366 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14302 10415 14366 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14302 10415 14366 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14302 10499 14366 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14302 10499 14366 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14378 9548 14442 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14378 9548 14442 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14378 11282 14442 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14378 11282 14442 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14383 7352 14447 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14383 7352 14447 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14383 7440 14447 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14383 7440 14447 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14383 7528 14447 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14383 7528 14447 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14383 7616 14447 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14383 7616 14447 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14383 7704 14447 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14383 7704 14447 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14383 7792 14447 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14383 7792 14447 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14383 7880 14447 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14383 7880 14447 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14383 7968 14447 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14383 7968 14447 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14383 10331 14447 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14383 10331 14447 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14383 10415 14447 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14383 10415 14447 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14383 10499 14447 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14383 10499 14447 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14460 9548 14524 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14460 9548 14524 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14460 11282 14524 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14460 11282 14524 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14464 7352 14528 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14464 7352 14528 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14464 7440 14528 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14464 7440 14528 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14464 7528 14528 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14464 7528 14528 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14464 7616 14528 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14464 7616 14528 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14464 7704 14528 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14464 7704 14528 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14464 7792 14528 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14464 7792 14528 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14464 7880 14528 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14464 7880 14528 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14464 7968 14528 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14464 7968 14528 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14464 10331 14528 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14464 10331 14528 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14464 10415 14528 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14464 10415 14528 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14464 10499 14528 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14464 10499 14528 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14542 9548 14606 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14542 9548 14606 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14542 11282 14606 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14542 11282 14606 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14545 7352 14609 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14545 7352 14609 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14545 7440 14609 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14545 7440 14609 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14545 7528 14609 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14545 7528 14609 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14545 7616 14609 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14545 7616 14609 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14545 7704 14609 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14545 7704 14609 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14545 7792 14609 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14545 7792 14609 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14545 7880 14609 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14545 7880 14609 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14545 7968 14609 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14545 7968 14609 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14545 10331 14609 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14545 10331 14609 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14545 10415 14609 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14545 10415 14609 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14545 10499 14609 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14545 10499 14609 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14624 9548 14688 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14624 9548 14688 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14624 11282 14688 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14624 11282 14688 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14626 7352 14690 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14626 7352 14690 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14626 7440 14690 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14626 7440 14690 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14626 7528 14690 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14626 7528 14690 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14626 7616 14690 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14626 7616 14690 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14626 7704 14690 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14626 7704 14690 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14626 7792 14690 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14626 7792 14690 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14626 7880 14690 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14626 7880 14690 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14626 7968 14690 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14626 7968 14690 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14626 10331 14690 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14626 10331 14690 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14626 10415 14690 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14626 10415 14690 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14626 10499 14690 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14626 10499 14690 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14706 9548 14770 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14706 9548 14770 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14706 11282 14770 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14706 11282 14770 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14707 7352 14771 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14707 7352 14771 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14707 7440 14771 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14707 7440 14771 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14707 7528 14771 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14707 7528 14771 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14707 7616 14771 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14707 7616 14771 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14707 7704 14771 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14707 7704 14771 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14707 7792 14771 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14707 7792 14771 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14707 7880 14771 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14707 7880 14771 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14707 7968 14771 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14707 7968 14771 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14707 10331 14771 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14707 10331 14771 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14707 10415 14771 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14707 10415 14771 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14707 10499 14771 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14707 10499 14771 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14788 7352 14852 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14788 7352 14852 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14788 7440 14852 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14788 7440 14852 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14788 7528 14852 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14788 7528 14852 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14788 7616 14852 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14788 7616 14852 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14788 7704 14852 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14788 7704 14852 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14788 7792 14852 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14788 7792 14852 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14788 7880 14852 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14788 7880 14852 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14788 7968 14852 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14788 7968 14852 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14788 9548 14852 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14788 9548 14852 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14788 10331 14852 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14788 10331 14852 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14788 10415 14852 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14788 10415 14852 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14788 10499 14852 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14788 10499 14852 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 14788 11282 14852 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 14788 11282 14852 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1650 10331 1714 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1650 10331 1714 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1650 10415 1714 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1650 10415 1714 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1650 10499 1714 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1650 10499 1714 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1651 9548 1715 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1651 9548 1715 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1651 11282 1715 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1651 11282 1715 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1658 7352 1722 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1658 7352 1722 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1658 7440 1722 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1658 7440 1722 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1658 7528 1722 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1658 7528 1722 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1658 7616 1722 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1658 7616 1722 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1658 7704 1722 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1658 7704 1722 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1658 7792 1722 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1658 7792 1722 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1658 7880 1722 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1658 7880 1722 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1658 7968 1722 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1658 7968 1722 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1731 10331 1795 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1731 10331 1795 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1731 10415 1795 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1731 10415 1795 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1731 10499 1795 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1731 10499 1795 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1732 9548 1796 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1732 9548 1796 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1732 11282 1796 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1732 11282 1796 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1739 7352 1803 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1739 7352 1803 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1739 7440 1803 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1739 7440 1803 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1739 7528 1803 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1739 7528 1803 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1739 7616 1803 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1739 7616 1803 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1739 7704 1803 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1739 7704 1803 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1739 7792 1803 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1739 7792 1803 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1739 7880 1803 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1739 7880 1803 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1739 7968 1803 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1739 7968 1803 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1812 10331 1876 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1812 10331 1876 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1812 10415 1876 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1812 10415 1876 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1812 10499 1876 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1812 10499 1876 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1813 9548 1877 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1813 9548 1877 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1813 11282 1877 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1813 11282 1877 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1820 7352 1884 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1820 7352 1884 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1820 7440 1884 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1820 7440 1884 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1820 7528 1884 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1820 7528 1884 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1820 7616 1884 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1820 7616 1884 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1820 7704 1884 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1820 7704 1884 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1820 7792 1884 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1820 7792 1884 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1820 7880 1884 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1820 7880 1884 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1820 7968 1884 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1820 7968 1884 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1893 10331 1957 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1893 10331 1957 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1893 10415 1957 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1893 10415 1957 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1893 10499 1957 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1893 10499 1957 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1894 9548 1958 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1894 9548 1958 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1894 11282 1958 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1894 11282 1958 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1901 7352 1965 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1901 7352 1965 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1901 7440 1965 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1901 7440 1965 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1901 7528 1965 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1901 7528 1965 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1901 7616 1965 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1901 7616 1965 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1901 7704 1965 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1901 7704 1965 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1901 7792 1965 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1901 7792 1965 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1901 7880 1965 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1901 7880 1965 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1901 7968 1965 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1901 7968 1965 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1974 10331 2038 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1974 10331 2038 10395 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1974 10415 2038 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1974 10415 2038 10479 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1974 10499 2038 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1974 10499 2038 10563 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1975 9548 2039 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1975 9548 2039 9612 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1975 11282 2039 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1975 11282 2039 11346 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1982 7352 2046 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1982 7352 2046 7416 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1982 7440 2046 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1982 7440 2046 7504 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1982 7528 2046 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1982 7528 2046 7592 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1982 7616 2046 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1982 7616 2046 7680 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1982 7704 2046 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1982 7704 2046 7768 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1982 7792 2046 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1982 7792 2046 7856 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1982 7880 2046 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1982 7880 2046 7944 1 VSSA
port 39 nsew ground bidirectional
rlabel metal4 s 1982 7968 2046 8032 1 VSSA
port 39 nsew ground bidirectional
rlabel metal3 s 1982 7968 2046 8032 1 VSSA
port 39 nsew ground bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 15000 40000
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string LEFsymmetry X Y R90
string GDS_END 31743216
string GDS_START 31636320
<< end >>
