magic
tech sky130A
magscale 1 2
timestamp 1640697980
<< nwell >>
rect -38 261 1786 582
<< pwell >>
rect 63 21 1745 203
rect 29 -17 63 17
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 39 291 83 527
rect 217 291 266 527
rect 409 367 459 527
rect 577 367 627 527
rect 745 367 795 527
rect 913 367 963 527
rect 1081 323 1131 425
rect 1249 323 1299 425
rect 1417 323 1467 425
rect 1585 323 1635 425
rect 1081 289 1731 323
rect 17 213 115 257
rect 1054 215 1602 255
rect 17 51 53 213
rect 87 17 131 179
rect 1636 181 1731 289
rect 265 17 367 181
rect 401 145 1731 181
rect 401 51 467 145
rect 501 17 535 111
rect 569 51 635 145
rect 669 17 703 111
rect 737 51 803 145
rect 837 17 871 111
rect 905 51 971 145
rect 1005 17 1039 111
rect 1073 51 1139 145
rect 1173 17 1207 111
rect 1241 51 1307 145
rect 1341 17 1375 111
rect 1409 51 1475 145
rect 1509 17 1543 111
rect 1577 51 1643 145
rect 1677 17 1731 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< obsli1 >>
rect 117 291 183 493
rect 311 333 375 493
rect 493 333 543 493
rect 661 333 711 493
rect 829 333 879 493
rect 997 459 1719 493
rect 997 333 1047 459
rect 311 291 1047 333
rect 1165 357 1215 459
rect 1333 357 1383 459
rect 1501 357 1551 459
rect 1669 357 1719 459
rect 149 257 183 291
rect 149 215 1000 257
rect 149 213 231 215
rect 165 51 231 213
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
rlabel locali s 17 51 53 213 6 A
port 1 nsew signal input
rlabel locali s 17 213 115 257 6 A
port 1 nsew signal input
rlabel locali s 1054 215 1602 255 6 SLEEP
port 2 nsew signal input
rlabel metal1 s 0 -48 1748 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1685 -17 1719 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1593 -17 1627 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1501 -17 1535 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1409 -17 1443 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1317 -17 1351 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1225 -17 1259 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1133 -17 1167 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 1041 -17 1075 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 949 -17 983 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 857 -17 891 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 765 -17 799 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 673 -17 707 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 581 -17 615 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 489 -17 523 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 397 -17 431 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 305 -17 339 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 213 -17 247 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 121 -17 155 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel viali s 29 -17 63 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 0 -17 1748 17 8 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1677 17 1731 111 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1509 17 1543 111 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1341 17 1375 111 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1173 17 1207 111 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 1005 17 1039 111 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 837 17 871 111 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 669 17 703 111 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 501 17 535 111 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 265 17 367 181 6 VGND
port 3 nsew ground bidirectional abutment
rlabel locali s 87 17 131 179 6 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1786 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1748 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 1685 527 1719 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 1593 527 1627 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 1501 527 1535 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 1409 527 1443 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 1317 527 1351 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 1225 527 1259 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 1133 527 1167 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 1041 527 1075 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 949 527 983 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 857 527 891 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 765 527 799 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 673 527 707 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 581 527 615 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 489 527 523 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 397 527 431 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 305 527 339 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 213 527 247 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 121 527 155 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel viali s 29 527 63 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 913 367 963 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 745 367 795 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 577 367 627 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 409 367 459 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 217 291 266 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 39 291 83 527 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 0 527 1748 561 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1577 51 1643 145 6 X
port 7 nsew signal output
rlabel locali s 1409 51 1475 145 6 X
port 7 nsew signal output
rlabel locali s 1241 51 1307 145 6 X
port 7 nsew signal output
rlabel locali s 1073 51 1139 145 6 X
port 7 nsew signal output
rlabel locali s 905 51 971 145 6 X
port 7 nsew signal output
rlabel locali s 737 51 803 145 6 X
port 7 nsew signal output
rlabel locali s 569 51 635 145 6 X
port 7 nsew signal output
rlabel locali s 401 51 467 145 6 X
port 7 nsew signal output
rlabel locali s 401 145 1731 181 6 X
port 7 nsew signal output
rlabel locali s 1636 181 1731 289 6 X
port 7 nsew signal output
rlabel locali s 1081 289 1731 323 6 X
port 7 nsew signal output
rlabel locali s 1585 323 1635 425 6 X
port 7 nsew signal output
rlabel locali s 1417 323 1467 425 6 X
port 7 nsew signal output
rlabel locali s 1249 323 1299 425 6 X
port 7 nsew signal output
rlabel locali s 1081 323 1131 425 6 X
port 7 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1748 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2398866
string GDS_START 2385564
<< end >>
